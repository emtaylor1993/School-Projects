# 
# LEF OUT API 
# User Name : edbab 
# Date : Fri Aug 28 17:39:05 2009
# 
VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
 TIME NANOSECONDS 1 ;
 CAPACITANCE PICOFARADS 1 ;
 RESISTANCE OHMS 1 ;
 DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;
LAYER NWELL
 TYPE MASTERSLICE ;
END NWELL

LAYER DIFF
 TYPE MASTERSLICE ;
END DIFF

LAYER PIMP
 TYPE MASTERSLICE ;
END PIMP

LAYER NIMP
 TYPE MASTERSLICE ;
END NIMP

LAYER DIFF_25
 TYPE MASTERSLICE ;
END DIFF_25

LAYER SBLK
 TYPE MASTERSLICE ;
END SBLK

LAYER M1PIN
 TYPE MASTERSLICE ;
END M1PIN

LAYER M2PIN
 TYPE MASTERSLICE ;
END M2PIN

LAYER M3PIN
 TYPE MASTERSLICE ;
END M3PIN

LAYER M4PIN
 TYPE MASTERSLICE ;
END M4PIN

LAYER M5PIN
 TYPE MASTERSLICE ;
END M5PIN

LAYER M6PIN
 TYPE MASTERSLICE ;
END M6PIN

LAYER M7PIN
 TYPE MASTERSLICE ;
END M7PIN

LAYER M8PIN
 TYPE MASTERSLICE ;
END M8PIN

LAYER M9PIN
 TYPE MASTERSLICE ;
END M9PIN

LAYER IP
 TYPE MASTERSLICE ;
END IP

LAYER PO
 TYPE MASTERSLICE ;
END PO

LAYER CO
 TYPE CUT ;
 SPACING 0.13 ;
END CO

LAYER M1
 TYPE ROUTING ;
 PITCH 0.32 ;
 OFFSET 0.16 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.14 ;
 SPACING 0.14 ;
 ANTENNASIDEAREARATIO 1000 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.06 1000 ) ( 0.060001 43027.4 ) ( 1.06 43483.4 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
END M1

LAYER VIA1
 TYPE CUT ;
 SPACING 0.16 ;
END VIA1

LAYER M2
 TYPE ROUTING ;
 PITCH 0.32 ;
 OFFSET 0.16 ;
 DIRECTION VERTICAL ;
 WIDTH 0.16 ;
 SPACING 0.16 ;
 ANTENNASIDEAREARATIO 1000 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.06 1000 ) ( 0.060001 43027.4 ) ( 1.06 43483.4 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
END M2

LAYER VIA2
 TYPE CUT ;
 SPACING 0.16 ;
END VIA2

LAYER M3
 TYPE ROUTING ;
 PITCH 0.32 ;
 OFFSET 0.16 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.16 ;
 SPACING 0.16 ;
 ANTENNASIDEAREARATIO 1000 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.06 1000 ) ( 0.060001 43027.4 ) ( 1.06 43483.4 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
END M3

LAYER VIA3
 TYPE CUT ;
 SPACING 0.16 ;
END VIA3

LAYER M4
 TYPE ROUTING ;
 PITCH 0.32 ;
 OFFSET 0.16 ;
 DIRECTION VERTICAL ;
 WIDTH 0.16 ;
 SPACING 0.16 ;
 ANTENNASIDEAREARATIO 1000 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.06 1000 ) ( 0.060001 43027.4 ) ( 1.06 43483.4 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
END M4

LAYER VIA4
 TYPE CUT ;
 SPACING 0.16 ;
END VIA4

LAYER M5
 TYPE ROUTING ;
 PITCH 0.32 ;
 OFFSET 0.16 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.16 ;
 SPACING 0.16 ;
 ANTENNASIDEAREARATIO 1000 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.06 1000 ) ( 0.060001 43027.4 ) ( 1.06 43483.4 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
END M5

LAYER VIA5
 TYPE CUT ;
 SPACING 0.16 ;
END VIA5

LAYER M6
 TYPE ROUTING ;
 PITCH 0.32 ;
 OFFSET 0.16 ;
 DIRECTION VERTICAL ;
 WIDTH 0.16 ;
 SPACING 0.16 ;
 ANTENNASIDEAREARATIO 1000 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.06 1000 ) ( 0.060001 43027.4 ) ( 1.06 43483.4 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
END M6

LAYER VIA6
 TYPE CUT ;
 SPACING 0.16 ;
END VIA6

LAYER M7
 TYPE ROUTING ;
 PITCH 0.32 ;
 OFFSET 0.16 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.16 ;
 SPACING 0.16 ;
 ANTENNASIDEAREARATIO 1000 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.06 1000 ) ( 0.060001 43027.4 ) ( 1.06 43483.4 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
END M7

LAYER VIA7
 TYPE CUT ;
 SPACING 0.16 ;
END VIA7

LAYER M8
 TYPE ROUTING ;
 PITCH 0.32 ;
 OFFSET 0.16 ;
 DIRECTION VERTICAL ;
 WIDTH 0.16 ;
 SPACING 0.16 ;
 ANTENNASIDEAREARATIO 1000 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.06 1000 ) ( 0.060001 43027.4 ) ( 1.06 43483.4 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
END M8

LAYER VIA8
 TYPE CUT ;
 SPACING 0.34 ;
END VIA8

LAYER M9
 TYPE ROUTING ;
 PITCH 0.32 ;
 OFFSET 0.16 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.45 ;
 SPACING 0.45 ;
 ANTENNASIDEAREARATIO 1000 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.06 1000 ) ( 0.060001 50480 ) ( 1.06 58480 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
END M9

LAYER OverlapCheck
 TYPE OVERLAP ;
END OverlapCheck

VIA VIA12A DEFAULT
 RESISTANCE 1.6 ;
 LAYER VIA1 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 LAYER M1 ;
 RECT -0.12 -0.075 0.12 0.075 ;
 LAYER M2 ;
 RECT -0.12 -0.075 0.12 0.075 ;
END VIA12A

VIARULE VIA12A GENERATE
 LAYER M1 ;
 DIRECTION HORIZONTAL ;
 OVERHANG 0.05 ;
 LAYER M2 ;
 DIRECTION VERTICAL ;
 OVERHANG 0.005 ;
 LAYER VIA1 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 SPACING 0.3 BY 0.3 ;
 RESISTANCE 1.6 ;
END VIA12A

VIA VIA23 DEFAULT
 RESISTANCE 1.6 ;
 LAYER VIA2 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 LAYER M2 ;
 RECT -0.12 -0.075 0.12 0.075 ;
 LAYER M3 ;
 RECT -0.12 -0.075 0.12 0.075 ;
END VIA23

VIARULE VIA23 GENERATE
 LAYER M2 ;
 DIRECTION HORIZONTAL ;
 OVERHANG 0.05 ;
 LAYER M3 ;
 DIRECTION VERTICAL ;
 OVERHANG 0.005 ;
 LAYER VIA2 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 SPACING 0.3 BY 0.3 ;
 RESISTANCE 1.6 ;
END VIA23

VIA VIA34 DEFAULT
 RESISTANCE 1.6 ;
 LAYER VIA3 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 LAYER M3 ;
 RECT -0.12 -0.075 0.12 0.075 ;
 LAYER M4 ;
 RECT -0.12 -0.075 0.12 0.075 ;
END VIA34

VIARULE VIA34 GENERATE
 LAYER M3 ;
 DIRECTION HORIZONTAL ;
 OVERHANG 0.05 ;
 LAYER M4 ;
 DIRECTION VERTICAL ;
 OVERHANG 0.005 ;
 LAYER VIA3 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 SPACING 0.3 BY 0.3 ;
 RESISTANCE 1.6 ;
END VIA34

VIA VIA45 DEFAULT
 RESISTANCE 1.6 ;
 LAYER VIA4 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 LAYER M4 ;
 RECT -0.12 -0.075 0.12 0.075 ;
 LAYER M5 ;
 RECT -0.12 -0.075 0.12 0.075 ;
END VIA45

VIARULE VIA45 GENERATE
 LAYER M4 ;
 DIRECTION HORIZONTAL ;
 OVERHANG 0.05 ;
 LAYER M5 ;
 DIRECTION VERTICAL ;
 OVERHANG 0.005 ;
 LAYER VIA4 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 SPACING 0.3 BY 0.3 ;
 RESISTANCE 1.6 ;
END VIA45

VIA VIA56 DEFAULT
 RESISTANCE 1.6 ;
 LAYER VIA5 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 LAYER M5 ;
 RECT -0.12 -0.075 0.12 0.075 ;
 LAYER M6 ;
 RECT -0.12 -0.075 0.12 0.075 ;
END VIA56

VIARULE VIA56 GENERATE
 LAYER M5 ;
 DIRECTION HORIZONTAL ;
 OVERHANG 0.05 ;
 LAYER M6 ;
 DIRECTION VERTICAL ;
 OVERHANG 0.005 ;
 LAYER VIA5 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 SPACING 0.3 BY 0.3 ;
 RESISTANCE 1.6 ;
END VIA56

VIA VIA67 DEFAULT
 RESISTANCE 1.6 ;
 LAYER VIA6 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 LAYER M6 ;
 RECT -0.12 -0.075 0.12 0.075 ;
 LAYER M7 ;
 RECT -0.12 -0.075 0.12 0.075 ;
END VIA67

VIARULE VIA67 GENERATE
 LAYER M6 ;
 DIRECTION HORIZONTAL ;
 OVERHANG 0.05 ;
 LAYER M7 ;
 DIRECTION VERTICAL ;
 OVERHANG 0.005 ;
 LAYER VIA6 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 SPACING 0.3 BY 0.3 ;
 RESISTANCE 1.6 ;
END VIA67

VIA VIA78 DEFAULT
 RESISTANCE 1.6 ;
 LAYER VIA7 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 LAYER M7 ;
 RECT -0.12 -0.075 0.12 0.075 ;
 LAYER M8 ;
 RECT -0.12 -0.075 0.12 0.075 ;
END VIA78

VIARULE VIA78 GENERATE
 LAYER M7 ;
 DIRECTION HORIZONTAL ;
 OVERHANG 0.05 ;
 LAYER M8 ;
 DIRECTION VERTICAL ;
 OVERHANG 0.005 ;
 LAYER VIA7 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 SPACING 0.3 BY 0.3 ;
 RESISTANCE 1.6 ;
END VIA78

VIA VIA89 DEFAULT
 RESISTANCE 1.6 ;
 LAYER VIA8 ;
 RECT -0.18 -0.18 0.18 0.18 ;
 LAYER M8 ;
 RECT -0.26 -0.21 0.26 0.21 ;
 LAYER M9 ;
 RECT -0.26 -0.21 0.26 0.21 ;
END VIA89

VIARULE VIA89 GENERATE
 LAYER M8 ;
 DIRECTION HORIZONTAL ;
 OVERHANG 0.08 ;
 LAYER M9 ;
 DIRECTION VERTICAL ;
 OVERHANG 0.03 ;
 LAYER VIA8 ;
 RECT -0.18 -0.18 0.18 0.18 ;
 SPACING 0.7 BY 0.7 ;
 RESISTANCE 1.6 ;
END VIA89

VIA POLYCON 
 LAYER CO ;
 RECT -0.065 -0.065 0.065 0.065 ;
 LAYER PO ;
 RECT -0.115 -0.105 0.115 0.105 ;
 LAYER M1 ;
 RECT -0.115 -0.105 0.115 0.105 ;
END POLYCON

VIARULE POLYCON GENERATE
 LAYER PO ;
 DIRECTION HORIZONTAL ;
 OVERHANG 0.05 ;
 LAYER M1 ;
 DIRECTION VERTICAL ;
 OVERHANG 0.04 ;
 LAYER CO ;
 RECT -0.065 -0.065 0.065 0.065 ;
 SPACING 0.26 BY 0.26 ;
END POLYCON

VIA VIA12B DEFAULT
 RESISTANCE 1.6 ;
 LAYER VIA1 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 LAYER M1 ;
 RECT -0.075 -0.12 0.075 0.12 ;
 LAYER M2 ;
 RECT -0.12 -0.075 0.12 0.075 ;
END VIA12B

VIARULE VIA12B GENERATE
 LAYER M1 ;
 DIRECTION HORIZONTAL ;
 OVERHANG 0.005 ;
 LAYER M2 ;
 DIRECTION VERTICAL ;
 OVERHANG 0.005 ;
 LAYER VIA1 ;
 RECT -0.07 -0.07 0.07 0.07 ;
 SPACING 0.3 BY 0.3 ;
 RESISTANCE 1.6 ;
END VIA12B

SPACING
 SAMENET PO CO 0.12 ;
 SAMENET CO M1 0 ;
 SAMENET CO VIA1 0 STACK ;
 SAMENET M1 VIA1 0 ;
 SAMENET VIA1 M2 0 ;
 SAMENET VIA1 VIA2 0 STACK ;
 SAMENET M2 VIA2 0 ;
 SAMENET VIA2 M3 0 ;
 SAMENET M3 VIA3 0 ;
 SAMENET VIA2 VIA3 0 STACK ;
 SAMENET VIA3 M4 0 ;
 SAMENET VIA3 VIA4 0 STACK ;
 SAMENET M4 VIA4 0 ;
 SAMENET VIA4 M5 0 ;
 SAMENET M5 VIA5 0 ;
 SAMENET VIA4 VIA5 0 STACK ;
 SAMENET VIA5 M6 0 ;
 SAMENET M6 VIA6 0 ;
 SAMENET VIA5 VIA6 0 STACK ;
 SAMENET VIA6 M7 0 ;
 SAMENET M7 VIA7 0 ;
 SAMENET VIA6 VIA7 0 STACK ;
 SAMENET VIA7 M8 0 ;
 SAMENET M8 VIA8 0 ;
 SAMENET VIA7 VIA8 0 STACK ;
 SAMENET VIA8 M9 0 ;
END SPACING

END LIBRARY
