`timescale 1ns / 1ps

module mux2g(
    input a,
    input b,
    input s,
    output z
    );

endmodule
