# 
# LEF OUT API 
# User Name : stud732 
# Date : Tue Aug 31 09:49:08 2010
# 
VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
SITE unit
 CLASS CORE ;
 SIZE 0.32 BY 2.88 ;
END unit

MACRO CGLPPSX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.96 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.96 2.96 ;
 RECT 4.57 1.525 4.8 1.665 ;
 RECT 1.55 2.625 1.78 2.8 ;
 RECT 0.755 1.575 0.895 2.8 ;
 RECT 3.305 2.345 3.445 2.8 ;
 RECT 5.555 2.135 5.695 2.8 ;
 RECT 7 1.715 7.14 2.8 ;
 RECT 7.94 1.45 8.08 2.8 ;
 RECT 6.495 1.46 6.635 2.8 ;
 RECT 4.615 1.665 4.755 2.8 ;
 RECT 8.435 1.5 8.575 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 2.09 0.615 2.36 ;
 END
 ANTENNAGATEAREA 0.063 ;
 END CLK

 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 1.16 1.925 1.4 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.96 0.08 ;
 RECT 4.57 0.515 4.8 0.655 ;
 RECT 1.545 0.585 1.8 0.725 ;
 RECT 7 0.08 7.14 0.68 ;
 RECT 7.94 0.08 8.08 0.98 ;
 RECT 3.305 0.08 3.445 0.74 ;
 RECT 0.755 0.08 0.895 0.985 ;
 RECT 5.86 0.08 6 0.7 ;
 RECT 1.66 0.08 1.8 0.585 ;
 RECT 8.4 0.08 8.54 0.85 ;
 RECT 4.615 0.655 4.755 0.665 ;
 RECT 4.615 0.08 4.755 0.515 ;
 END
 END VSS

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.47 2.36 7.61 2.53 ;
 RECT 7.47 2.12 7.8 2.36 ;
 RECT 7.47 0.39 7.61 2.12 ;
 END
 ANTENNADIFFAREA 0.622 ;
 END GCLK

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.425 0.84 4.99 1.105 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END SE

 OBS
 LAYER PO ;
 RECT 4.4 0.93 4.69 1.14 ;
 RECT 4.4 0.28 4.5 0.93 ;
 RECT 4.4 1.14 4.5 1.88 ;
 RECT 4.87 0.29 4.97 2.09 ;
 RECT 3.56 1.1 3.66 2.09 ;
 RECT 3.555 2.09 4.97 2.19 ;
 RECT 3.56 0.35 3.66 0.89 ;
 RECT 3.405 0.89 3.66 1.1 ;
 RECT 1.85 1.4 1.95 2.14 ;
 RECT 1.85 0.37 1.95 1.19 ;
 RECT 1.685 1.19 1.95 1.4 ;
 RECT 2.79 0.315 2.89 0.89 ;
 RECT 2.32 1.26 2.42 2.03 ;
 RECT 2.71 0.89 2.89 0.99 ;
 RECT 2.71 0.99 2.81 1.16 ;
 RECT 2.32 1.16 2.81 1.26 ;
 RECT 2.245 2.03 2.475 2.24 ;
 RECT 2.79 1.56 2.89 2.35 ;
 RECT 2.73 2.35 2.94 2.58 ;
 RECT 3.09 0.315 3.19 1.17 ;
 RECT 3.09 1.38 3.19 2.14 ;
 RECT 2.99 1.17 3.22 1.38 ;
 RECT 5.17 1.2 5.405 1.23 ;
 RECT 5.17 0.295 5.27 1.2 ;
 RECT 5.175 1.33 5.44 1.41 ;
 RECT 5.34 1.41 5.44 1.88 ;
 RECT 5.17 1.23 5.44 1.33 ;
 RECT 5.81 0.85 5.91 2.52 ;
 RECT 6.115 0.28 6.215 0.75 ;
 RECT 4.245 2.41 4.475 2.52 ;
 RECT 4.245 2.52 5.91 2.62 ;
 RECT 5.81 0.75 6.215 0.85 ;
 RECT 6.945 1.02 7.355 1.23 ;
 RECT 7.255 0.195 7.355 1.02 ;
 RECT 7.725 0.195 7.825 1.23 ;
 RECT 7.725 1.33 7.825 2.76 ;
 RECT 7.255 1.33 7.355 2.76 ;
 RECT 7.255 1.23 7.825 1.33 ;
 RECT 6.415 0.28 6.515 1.28 ;
 RECT 6.28 1.38 6.38 1.82 ;
 RECT 6.28 1.28 6.515 1.38 ;
 RECT 6.12 1.82 6.38 2.03 ;
 RECT 0.82 1.15 1.11 1.36 ;
 RECT 1.01 0.19 1.11 1.15 ;
 RECT 1.01 1.36 1.11 2.31 ;
 RECT 2.32 0.19 2.42 0.885 ;
 RECT 0.13 0.09 2.42 0.19 ;
 RECT 1.01 2.31 1.285 2.52 ;
 RECT 0.13 0.19 0.36 0.4 ;
 RECT 0.54 0.57 0.64 2.12 ;
 RECT 0.385 2.12 0.64 2.33 ;
 LAYER CO ;
 RECT 3.455 0.93 3.585 1.06 ;
 RECT 7.475 0.5 7.605 0.63 ;
 RECT 0.29 1.585 0.42 1.715 ;
 RECT 0.29 0.79 0.42 0.92 ;
 RECT 7.005 0.5 7.135 0.63 ;
 RECT 1.105 2.35 1.235 2.48 ;
 RECT 3.04 1.21 3.17 1.34 ;
 RECT 7.005 2.03 7.135 2.16 ;
 RECT 6.635 0.5 6.765 0.63 ;
 RECT 3.31 2.395 3.44 2.525 ;
 RECT 7.945 0.505 8.075 0.635 ;
 RECT 0.76 0.79 0.89 0.92 ;
 RECT 2.295 2.07 2.425 2.2 ;
 RECT 7.945 1.5 8.075 1.63 ;
 RECT 4.51 0.97 4.64 1.1 ;
 RECT 8.44 2.07 8.57 2.2 ;
 RECT 7.945 0.765 8.075 0.895 ;
 RECT 6.5 1.51 6.63 1.64 ;
 RECT 1.23 0.79 1.36 0.92 ;
 RECT 1.23 2.04 1.36 2.17 ;
 RECT 7.475 2.03 7.605 2.16 ;
 RECT 1.6 2.63 1.73 2.76 ;
 RECT 2.77 2.4 2.9 2.53 ;
 RECT 3.78 0.6 3.91 0.73 ;
 RECT 7.475 2.29 7.605 2.42 ;
 RECT 7.475 1.5 7.605 1.63 ;
 RECT 2.07 1.78 2.2 1.91 ;
 RECT 5.225 1.24 5.355 1.37 ;
 RECT 4.295 2.45 4.425 2.58 ;
 RECT 6.17 1.86 6.3 1.99 ;
 RECT 5.56 2.185 5.69 2.315 ;
 RECT 4.62 1.53 4.75 1.66 ;
 RECT 6.03 1.51 6.16 1.64 ;
 RECT 0.87 1.19 1 1.32 ;
 RECT 0.435 2.16 0.565 2.29 ;
 RECT 5.865 0.5 5.995 0.63 ;
 RECT 4.15 1.53 4.28 1.66 ;
 RECT 4.15 0.52 4.28 0.65 ;
 RECT 0.76 1.625 0.89 1.755 ;
 RECT 7.945 2.29 8.075 2.42 ;
 RECT 7.475 0.765 7.605 0.895 ;
 RECT 2.54 0.535 2.67 0.665 ;
 RECT 4.62 0.52 4.75 0.65 ;
 RECT 1.74 1.23 1.87 1.36 ;
 RECT 7.475 1.765 7.605 1.895 ;
 RECT 6.995 1.06 7.125 1.19 ;
 RECT 5.39 0.52 5.52 0.65 ;
 RECT 8.405 0.41 8.535 0.54 ;
 RECT 5.09 1.53 5.22 1.66 ;
 RECT 7.005 2.29 7.135 2.42 ;
 RECT 8.44 1.55 8.57 1.68 ;
 RECT 2.07 0.59 2.2 0.72 ;
 RECT 8.44 1.81 8.57 1.94 ;
 RECT 7.945 2.03 8.075 2.16 ;
 RECT 7.945 1.765 8.075 1.895 ;
 RECT 0.18 0.23 0.31 0.36 ;
 RECT 3.31 0.535 3.44 0.665 ;
 RECT 3.78 1.78 3.91 1.91 ;
 RECT 2.54 1.78 2.67 1.91 ;
 RECT 1.6 0.59 1.73 0.72 ;
 RECT 8.405 0.67 8.535 0.8 ;
 RECT 7.005 1.765 7.135 1.895 ;
 LAYER M1 ;
 RECT 4.145 0.45 4.285 1.245 ;
 RECT 4.145 1.385 4.285 1.71 ;
 RECT 4.145 1.245 5.405 1.375 ;
 RECT 5.175 1.235 5.405 1.245 ;
 RECT 4.145 1.375 5.355 1.385 ;
 RECT 2.535 1.065 2.675 1.775 ;
 RECT 2.535 0.455 2.675 0.925 ;
 RECT 2.49 1.775 2.72 1.915 ;
 RECT 2.535 0.925 3.635 1.065 ;
 RECT 3.775 1.345 3.915 1.775 ;
 RECT 2.99 1.205 3.915 1.345 ;
 RECT 3.775 0.365 3.915 1.205 ;
 RECT 3.73 1.775 3.96 1.915 ;
 RECT 2.065 0.53 2.205 1.775 ;
 RECT 2.02 1.775 2.25 1.915 ;
 RECT 5.55 0.655 5.69 1.525 ;
 RECT 5.34 0.515 5.69 0.655 ;
 RECT 5.55 1.665 5.69 1.855 ;
 RECT 5.04 1.525 5.69 1.665 ;
 RECT 5.55 1.855 6.35 1.995 ;
 RECT 6.025 1.19 6.165 1.71 ;
 RECT 6.025 1.05 6.77 1.055 ;
 RECT 6.63 0.45 6.77 1.05 ;
 RECT 6.025 1.055 7.185 1.19 ;
 RECT 6.645 1.19 7.185 1.195 ;
 RECT 1.05 2.35 2.905 2.485 ;
 RECT 1.05 2.345 2.9 2.35 ;
 RECT 2.765 2.485 2.905 2.58 ;
 RECT 1.19 0.985 1.33 1.97 ;
 RECT 1.13 1.97 1.41 2.065 ;
 RECT 1.19 0.715 1.365 0.985 ;
 RECT 4.25 2.205 4.39 2.445 ;
 RECT 4.25 2.585 4.39 2.59 ;
 RECT 1.13 2.065 4.39 2.205 ;
 RECT 4.245 2.445 4.475 2.585 ;
 RECT 0.285 0.365 0.425 1.185 ;
 RECT 0.285 1.325 0.425 1.79 ;
 RECT 0.13 0.225 0.425 0.365 ;
 RECT 0.285 1.185 1.05 1.325 ;
 RECT 0.82 1.15 1.05 1.185 ;
 RECT 0.82 1.325 1.05 1.36 ;
 END
END CGLPPSX2

MACRO CGLPPSX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.92 BY 2.88 ;
 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.475 1.435 8.795 1.735 ;
 RECT 8.56 1.735 8.7 2.45 ;
 RECT 7.62 1.12 8.7 1.26 ;
 RECT 8.56 1.26 8.7 1.435 ;
 RECT 8.56 0.475 8.7 1.12 ;
 RECT 7.62 1.26 7.76 2.45 ;
 RECT 7.62 0.475 7.76 1.12 ;
 END
 ANTENNADIFFAREA 1.244 ;
 END GCLK

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.92 2.96 ;
 RECT 4.72 1.525 4.95 1.665 ;
 RECT 1.7 2.625 1.93 2.8 ;
 RECT 0.86 2.625 1.09 2.8 ;
 RECT 8.09 1.43 8.23 2.8 ;
 RECT 7.15 1.43 7.29 2.8 ;
 RECT 3.455 1.73 3.595 2.8 ;
 RECT 5.745 2.045 5.885 2.8 ;
 RECT 9.03 1.43 9.17 2.8 ;
 RECT 6.78 1.44 6.92 2.8 ;
 RECT 4.765 1.665 4.905 2.8 ;
 RECT 9.47 1.5 9.61 2.8 ;
 END
 END VDD

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.61 0.84 4.92 1.105 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END SE

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.475 2.07 0.835 2.39 ;
 END
 ANTENNAGATEAREA 0.063 ;
 END CLK

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.92 0.08 ;
 RECT 4.72 0.555 4.95 0.695 ;
 RECT 1.695 0.585 1.95 0.725 ;
 RECT 0.905 0.08 1.045 0.985 ;
 RECT 9.03 0.08 9.17 0.975 ;
 RECT 7.15 0.08 7.29 0.94 ;
 RECT 3.455 0.08 3.595 0.74 ;
 RECT 6.01 0.08 6.15 0.98 ;
 RECT 1.81 0.08 1.95 0.585 ;
 RECT 8.09 0.08 8.23 0.975 ;
 RECT 9.47 0.08 9.61 0.85 ;
 RECT 4.765 0.695 4.905 0.7 ;
 RECT 4.765 0.08 4.905 0.555 ;
 END
 END VSS

 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.755 1.12 2.07 1.445 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 OBS
 LAYER PO ;
 RECT 5.32 0.31 5.42 1.2 ;
 RECT 5.49 1.41 5.59 1.88 ;
 RECT 5.32 1.2 5.59 1.41 ;
 RECT 6.565 0.53 6.665 2.215 ;
 RECT 6.435 2.215 6.665 2.445 ;
 RECT 6.095 1.19 6.195 2.535 ;
 RECT 6.265 0.53 6.365 1.09 ;
 RECT 3.085 2.43 3.295 2.535 ;
 RECT 3.085 2.635 3.295 2.66 ;
 RECT 3.085 2.535 6.195 2.635 ;
 RECT 6.095 1.09 6.365 1.19 ;
 RECT 4.55 0.93 4.84 1.14 ;
 RECT 4.55 0.305 4.65 0.93 ;
 RECT 4.55 1.14 4.65 1.88 ;
 RECT 5.02 1.83 5.125 1.88 ;
 RECT 5.025 1.88 5.125 2.09 ;
 RECT 5.02 0.265 5.12 1.83 ;
 RECT 3.71 1.1 3.81 2.09 ;
 RECT 3.71 0.255 3.81 0.89 ;
 RECT 3.555 0.89 3.81 1.1 ;
 RECT 3.7 2.09 5.125 2.19 ;
 RECT 7.24 1.08 7.505 1.15 ;
 RECT 7.24 1.25 7.505 1.29 ;
 RECT 7.405 1.29 7.505 2.74 ;
 RECT 7.405 0.215 7.505 1.08 ;
 RECT 8.815 1.25 8.915 2.74 ;
 RECT 8.815 0.215 8.915 1.15 ;
 RECT 8.345 0.215 8.445 1.15 ;
 RECT 8.345 1.25 8.445 2.74 ;
 RECT 7.875 0.215 7.975 1.15 ;
 RECT 7.875 1.25 7.975 2.74 ;
 RECT 7.24 1.15 8.915 1.25 ;
 RECT 2 1.4 2.1 2.14 ;
 RECT 2 0.37 2.1 1.19 ;
 RECT 1.84 1.19 2.1 1.4 ;
 RECT 3.24 0.315 3.34 1.17 ;
 RECT 3.24 1.38 3.34 2.14 ;
 RECT 3.14 1.17 3.37 1.38 ;
 RECT 2.94 1.56 3.04 2.14 ;
 RECT 2.805 2.24 2.905 2.43 ;
 RECT 2.54 2.53 2.75 2.66 ;
 RECT 2.54 2.43 2.905 2.53 ;
 RECT 2.805 2.14 3.04 2.24 ;
 RECT 2.94 0.315 3.04 0.89 ;
 RECT 2.47 1.26 2.57 2.03 ;
 RECT 2.86 0.89 3.04 0.99 ;
 RECT 2.86 0.99 2.96 1.16 ;
 RECT 2.47 1.16 2.96 1.26 ;
 RECT 2.395 2.03 2.625 2.24 ;
 RECT 0.99 1.125 1.26 1.335 ;
 RECT 1.16 1.335 1.26 2.31 ;
 RECT 2.47 0.19 2.57 0.885 ;
 RECT 1.16 0.19 1.26 1.125 ;
 RECT 1.16 2.31 1.39 2.52 ;
 RECT 1.16 0.09 2.57 0.19 ;
 RECT 0.69 0.57 0.79 2.12 ;
 RECT 0.56 2.12 0.79 2.33 ;
 LAYER CO ;
 RECT 2.69 1.78 2.82 1.91 ;
 RECT 8.095 0.785 8.225 0.915 ;
 RECT 0.91 0.79 1.04 0.92 ;
 RECT 2.22 0.59 2.35 0.72 ;
 RECT 9.475 0.41 9.605 0.54 ;
 RECT 3.605 0.93 3.735 1.06 ;
 RECT 2.445 2.07 2.575 2.2 ;
 RECT 8.095 2.27 8.225 2.4 ;
 RECT 7.155 1.74 7.285 1.87 ;
 RECT 3.93 0.6 4.06 0.73 ;
 RECT 7.625 0.785 7.755 0.915 ;
 RECT 5.375 1.24 5.505 1.37 ;
 RECT 8.565 1.48 8.695 1.61 ;
 RECT 9.035 1.48 9.165 1.61 ;
 RECT 8.565 2.27 8.695 2.4 ;
 RECT 8.565 1.745 8.695 1.875 ;
 RECT 9.035 1.745 9.165 1.875 ;
 RECT 9.475 1.81 9.605 1.94 ;
 RECT 3.46 0.535 3.59 0.665 ;
 RECT 7.155 0.76 7.285 0.89 ;
 RECT 1.75 2.63 1.88 2.76 ;
 RECT 6.315 1.49 6.445 1.62 ;
 RECT 7.625 2.01 7.755 2.14 ;
 RECT 7.625 0.525 7.755 0.655 ;
 RECT 1.38 0.79 1.51 0.92 ;
 RECT 6.485 2.26 6.615 2.39 ;
 RECT 9.035 0.785 9.165 0.915 ;
 RECT 6.785 1.49 6.915 1.62 ;
 RECT 9.035 2.27 9.165 2.4 ;
 RECT 3.46 1.78 3.59 1.91 ;
 RECT 7.625 1.745 7.755 1.875 ;
 RECT 3.19 1.21 3.32 1.34 ;
 RECT 7.29 1.12 7.42 1.25 ;
 RECT 1.04 1.165 1.17 1.295 ;
 RECT 0.61 2.16 0.74 2.29 ;
 RECT 5.75 2.095 5.88 2.225 ;
 RECT 1.89 1.23 2.02 1.36 ;
 RECT 7.155 2.27 7.285 2.4 ;
 RECT 3.93 1.78 4.06 1.91 ;
 RECT 5.24 1.53 5.37 1.66 ;
 RECT 3.125 2.48 3.255 2.61 ;
 RECT 6.785 0.785 6.915 0.915 ;
 RECT 6.015 0.79 6.145 0.92 ;
 RECT 8.095 0.525 8.225 0.655 ;
 RECT 8.095 1.745 8.225 1.875 ;
 RECT 2.58 2.48 2.71 2.61 ;
 RECT 7.155 0.495 7.285 0.625 ;
 RECT 8.095 2.01 8.225 2.14 ;
 RECT 8.565 0.785 8.695 0.915 ;
 RECT 8.565 0.525 8.695 0.655 ;
 RECT 7.155 2.01 7.285 2.14 ;
 RECT 0.44 0.79 0.57 0.92 ;
 RECT 7.625 2.27 7.755 2.4 ;
 RECT 4.77 1.53 4.9 1.66 ;
 RECT 8.095 1.48 8.225 1.61 ;
 RECT 9.475 0.67 9.605 0.8 ;
 RECT 4.3 1.53 4.43 1.66 ;
 RECT 7.625 1.48 7.755 1.61 ;
 RECT 9.475 2.07 9.605 2.2 ;
 RECT 2.22 1.78 2.35 1.91 ;
 RECT 0.44 1.585 0.57 1.715 ;
 RECT 7.155 1.48 7.285 1.61 ;
 RECT 4.3 0.56 4.43 0.69 ;
 RECT 1.38 1.5 1.51 1.63 ;
 RECT 8.565 2.01 8.695 2.14 ;
 RECT 4.77 0.56 4.9 0.69 ;
 RECT 2.69 0.535 2.82 0.665 ;
 RECT 9.035 0.525 9.165 0.655 ;
 RECT 5.54 0.56 5.67 0.69 ;
 RECT 1.21 2.35 1.34 2.48 ;
 RECT 9.475 1.55 9.605 1.68 ;
 RECT 0.91 2.63 1.04 2.76 ;
 RECT 1.75 0.59 1.88 0.72 ;
 RECT 9.035 2.01 9.165 2.14 ;
 RECT 4.66 0.97 4.79 1.1 ;
 LAYER M1 ;
 RECT 2.215 0.53 2.355 1.775 ;
 RECT 2.17 1.775 2.4 1.915 ;
 RECT 6.78 0.72 6.92 1.11 ;
 RECT 6.77 1.11 6.92 1.115 ;
 RECT 6.31 1.255 6.45 1.485 ;
 RECT 6.265 1.485 6.495 1.625 ;
 RECT 6.31 1.115 7.47 1.255 ;
 RECT 5.7 1.665 5.84 1.765 ;
 RECT 5.7 0.695 5.84 1.525 ;
 RECT 5.19 1.525 5.84 1.665 ;
 RECT 5.49 0.555 5.84 0.695 ;
 RECT 6.48 1.905 6.62 2.445 ;
 RECT 5.7 1.765 6.62 1.905 ;
 RECT 1.16 2.345 2.715 2.485 ;
 RECT 2.575 2.485 2.715 2.66 ;
 RECT 2.685 1.065 2.825 1.775 ;
 RECT 2.685 0.455 2.825 0.925 ;
 RECT 2.64 1.775 2.87 1.915 ;
 RECT 2.685 0.925 3.785 1.065 ;
 RECT 4.295 0.425 4.435 1.245 ;
 RECT 4.295 1.385 4.435 1.71 ;
 RECT 5.325 1.235 5.555 1.245 ;
 RECT 4.295 1.245 5.555 1.385 ;
 RECT 3.925 1.345 4.065 1.775 ;
 RECT 3.14 1.205 4.065 1.345 ;
 RECT 3.925 0.365 4.065 1.205 ;
 RECT 3.88 1.775 4.11 1.915 ;
 RECT 1.375 0.715 1.515 2.065 ;
 RECT 3.12 2.205 3.26 2.66 ;
 RECT 1.375 2.065 3.26 2.205 ;
 RECT 0.435 0.635 0.575 1.16 ;
 RECT 0.435 1.3 0.575 1.785 ;
 RECT 0.99 1.125 1.22 1.16 ;
 RECT 0.99 1.3 1.22 1.335 ;
 RECT 0.435 1.16 1.22 1.3 ;
 END
END CGLPPSX4

MACRO ISOLANDX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.515 1.445 0.905 1.725 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END ISO

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.455 1.115 1.735 1.325 ;
 RECT 1.455 1.325 1.84 1.405 ;
 RECT 1.555 1.405 1.84 1.72 ;
 END
 ANTENNAGATEAREA 0.058 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.235 1.195 2.965 1.425 ;
 RECT 2.675 1.16 2.965 1.195 ;
 RECT 2.235 1.425 2.375 2.505 ;
 RECT 2.32 0.365 2.46 1.195 ;
 END
 ANTENNADIFFAREA 0.83 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 1.645 1.885 1.785 2.8 ;
 RECT 0.63 2.14 0.845 2.28 ;
 RECT 0.91 2.48 1.395 2.8 ;
 RECT 0.63 2.28 0.77 2.8 ;
 RECT 2.8 1.61 2.94 2.8 ;
 RECT 0.705 1.87 0.845 2.14 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 0.64 0.75 0.905 0.89 ;
 RECT 1.025 0.08 1.515 0.42 ;
 RECT 1.85 0.08 1.99 0.57 ;
 RECT 2.8 0.08 2.94 0.57 ;
 RECT 0.705 0.08 0.845 0.75 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.96 0.51 1.06 1.06 ;
 RECT 0.96 1.29 1.06 2.4 ;
 RECT 0.83 1.06 1.06 1.29 ;
 RECT 0.49 0.515 0.59 1.47 ;
 RECT 0.49 1.7 0.59 2.41 ;
 RECT 0.485 1.47 0.715 1.7 ;
 RECT 1.26 1.125 1.675 1.265 ;
 RECT 1.26 0.51 1.36 1.125 ;
 RECT 1.43 1.265 1.675 1.355 ;
 RECT 1.43 1.355 1.53 2.405 ;
 RECT 1.9 0.99 2.675 1.09 ;
 RECT 2.575 0.1 2.675 0.99 ;
 RECT 1.9 0.86 2.205 0.99 ;
 RECT 2.575 1.09 2.675 2.775 ;
 RECT 1.9 1.09 2 2.775 ;
 RECT 2.105 0.1 2.205 0.86 ;
 LAYER CO ;
 RECT 2.805 0.39 2.935 0.52 ;
 RECT 2.805 1.66 2.935 1.79 ;
 RECT 2.805 2.305 2.935 2.435 ;
 RECT 2.805 1.965 2.935 2.095 ;
 RECT 1.335 0.255 1.465 0.385 ;
 RECT 1.075 0.255 1.205 0.385 ;
 RECT 1.22 2.53 1.35 2.66 ;
 RECT 0.96 2.53 1.09 2.66 ;
 RECT 1.95 0.91 2.08 1.04 ;
 RECT 1.495 1.175 1.625 1.305 ;
 RECT 0.88 1.11 1.01 1.24 ;
 RECT 2.325 0.42 2.455 0.55 ;
 RECT 2.24 1.6 2.37 1.73 ;
 RECT 2.24 1.93 2.37 2.06 ;
 RECT 2.24 2.305 2.37 2.435 ;
 RECT 1.855 0.39 1.985 0.52 ;
 RECT 1.65 2.305 1.78 2.435 ;
 RECT 0.535 1.52 0.665 1.65 ;
 RECT 1.48 0.755 1.61 0.885 ;
 RECT 1.65 1.965 1.78 2.095 ;
 RECT 1.18 1.93 1.31 2.06 ;
 RECT 0.71 0.755 0.84 0.885 ;
 RECT 0.71 1.93 0.84 2.06 ;
 RECT 0.24 0.755 0.37 0.885 ;
 RECT 0.24 1.93 0.37 2.06 ;
 LAYER M1 ;
 RECT 0.235 0.645 0.375 1.105 ;
 RECT 0.235 1.245 0.375 2.11 ;
 RECT 0.875 1.04 1.015 1.105 ;
 RECT 0.875 1.245 1.015 1.3 ;
 RECT 0.235 1.105 1.015 1.245 ;
 RECT 1.175 0.89 1.315 2.11 ;
 RECT 1.88 0.89 2.13 1.045 ;
 RECT 1.175 0.75 2.13 0.89 ;
 END
END ISOLANDX2

MACRO ISOLANDX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.395 1.445 0.76 1.725 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END ISO

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.335 1.275 1.715 1.615 ;
 RECT 1.335 1.115 1.615 1.275 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.115 1.215 3.29 1.355 ;
 RECT 2.505 1.355 2.935 1.425 ;
 RECT 2.505 1.16 2.935 1.215 ;
 RECT 2.115 1.355 2.255 2.505 ;
 RECT 2.2 0.365 2.34 1.215 ;
 RECT 3.15 1.355 3.29 2.505 ;
 RECT 3.15 0.295 3.29 1.215 ;
 END
 ANTENNADIFFAREA 1.446 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 0.51 2.14 0.725 2.28 ;
 RECT 0.79 2.48 1.275 2.8 ;
 RECT 0.51 2.28 0.65 2.8 ;
 RECT 1.525 1.805 1.665 2.8 ;
 RECT 2.68 1.61 2.82 2.8 ;
 RECT 3.65 1.61 3.79 2.8 ;
 RECT 0.585 1.87 0.725 2.14 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 0.52 0.76 0.785 0.9 ;
 RECT 0.905 0.08 1.395 0.42 ;
 RECT 1.73 0.08 1.87 0.57 ;
 RECT 2.68 0.08 2.82 0.57 ;
 RECT 3.64 0.08 3.78 0.57 ;
 RECT 0.585 0.08 0.725 0.76 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.84 0.51 0.94 1.06 ;
 RECT 0.84 1.29 0.94 2.315 ;
 RECT 0.71 1.06 0.94 1.29 ;
 RECT 0.37 0.515 0.47 1.47 ;
 RECT 0.37 1.7 0.47 2.405 ;
 RECT 0.37 1.47 0.595 1.7 ;
 RECT 1.14 1.125 1.555 1.265 ;
 RECT 1.14 0.51 1.24 1.125 ;
 RECT 1.31 1.265 1.555 1.355 ;
 RECT 1.31 1.355 1.41 2.37 ;
 RECT 1.78 0.99 3.515 1.09 ;
 RECT 3.415 0.1 3.515 0.99 ;
 RECT 2.935 0.1 3.035 0.99 ;
 RECT 2.455 0.1 2.555 0.99 ;
 RECT 1.78 0.89 2.085 0.99 ;
 RECT 3.415 1.09 3.515 2.775 ;
 RECT 2.935 1.09 3.035 2.775 ;
 RECT 2.455 1.09 2.555 2.775 ;
 RECT 1.78 1.12 1.88 2.775 ;
 RECT 1.985 0.1 2.085 0.89 ;
 RECT 1.78 1.09 2.01 1.12 ;
 LAYER CO ;
 RECT 3.645 0.39 3.775 0.52 ;
 RECT 3.155 0.39 3.285 0.52 ;
 RECT 3.655 1.66 3.785 1.79 ;
 RECT 3.655 2.305 3.785 2.435 ;
 RECT 3.655 1.965 3.785 2.095 ;
 RECT 3.155 1.6 3.285 1.73 ;
 RECT 3.155 1.93 3.285 2.06 ;
 RECT 3.155 2.305 3.285 2.435 ;
 RECT 2.685 0.39 2.815 0.52 ;
 RECT 2.685 1.66 2.815 1.79 ;
 RECT 2.685 2.305 2.815 2.435 ;
 RECT 2.685 1.965 2.815 2.095 ;
 RECT 1.215 0.255 1.345 0.385 ;
 RECT 0.955 0.255 1.085 0.385 ;
 RECT 1.1 2.53 1.23 2.66 ;
 RECT 0.84 2.53 0.97 2.66 ;
 RECT 1.83 0.94 1.96 1.07 ;
 RECT 1.375 1.175 1.505 1.305 ;
 RECT 0.76 1.11 0.89 1.24 ;
 RECT 2.205 0.42 2.335 0.55 ;
 RECT 2.12 1.6 2.25 1.73 ;
 RECT 2.12 1.93 2.25 2.06 ;
 RECT 2.12 2.305 2.25 2.435 ;
 RECT 1.735 0.39 1.865 0.52 ;
 RECT 1.53 2.305 1.66 2.435 ;
 RECT 0.415 1.52 0.545 1.65 ;
 RECT 1.36 0.765 1.49 0.895 ;
 RECT 1.53 1.965 1.66 2.095 ;
 RECT 1.06 1.93 1.19 2.06 ;
 RECT 0.59 0.765 0.72 0.895 ;
 RECT 0.59 1.93 0.72 2.06 ;
 RECT 0.12 0.765 0.25 0.895 ;
 RECT 0.12 1.93 0.25 2.06 ;
 LAYER M1 ;
 RECT 0.115 0.645 0.255 1.105 ;
 RECT 0.115 1.245 0.255 2.11 ;
 RECT 0.755 1.04 0.895 1.105 ;
 RECT 0.755 1.245 0.895 1.3 ;
 RECT 0.115 1.105 0.895 1.245 ;
 RECT 1.055 0.9 1.195 2.11 ;
 RECT 1.76 0.75 2.01 0.76 ;
 RECT 1.76 0.9 2.01 1.075 ;
 RECT 1.055 0.76 2.01 0.9 ;
 RECT 1.825 1.075 1.965 1.09 ;
 END
END ISOLANDX4

MACRO ISOLANDX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.4 BY 2.88 ;
 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.715 1.445 1.125 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END ISO

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.655 1.275 2.095 1.63 ;
 RECT 1.655 1.115 1.935 1.275 ;
 END
 ANTENNAGATEAREA 0.11 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.78 1.355 4.21 1.425 ;
 RECT 3.78 1.145 4.21 1.215 ;
 RECT 2.435 1.355 2.575 2.505 ;
 RECT 2.52 0.365 2.66 1.215 ;
 RECT 3.47 1.355 3.61 2.505 ;
 RECT 3.47 0.295 3.61 1.215 ;
 RECT 5.49 1.355 5.63 2.505 ;
 RECT 2.435 1.215 5.63 1.355 ;
 RECT 5.49 0.295 5.63 1.215 ;
 RECT 4.455 1.355 4.595 2.505 ;
 RECT 4.455 0.305 4.595 1.215 ;
 END
 ANTENNADIFFAREA 2.822 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.4 2.96 ;
 RECT 3 1.61 3.14 2.8 ;
 RECT 0.83 2.14 1.045 2.28 ;
 RECT 1.11 2.48 1.595 2.8 ;
 RECT 0.83 2.28 0.97 2.8 ;
 RECT 1.845 1.855 1.985 2.8 ;
 RECT 3.97 1.61 4.11 2.8 ;
 RECT 5.99 1.61 6.13 2.8 ;
 RECT 5.02 1.61 5.16 2.8 ;
 RECT 0.905 1.87 1.045 2.14 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.4 0.08 ;
 RECT 3 0.08 3.14 0.57 ;
 RECT 0.84 0.75 1.105 0.89 ;
 RECT 0.275 0.08 0.765 0.42 ;
 RECT 2.05 0.08 2.19 0.57 ;
 RECT 3.96 0.08 4.1 0.57 ;
 RECT 5.02 0.08 5.16 0.57 ;
 RECT 5.98 0.08 6.12 0.57 ;
 RECT 0.905 0.08 1.045 0.75 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.69 0.515 0.79 1.47 ;
 RECT 0.69 1.7 0.79 2.405 ;
 RECT 0.68 1.47 0.91 1.7 ;
 RECT 2.1 0.99 5.855 1.09 ;
 RECT 4.225 1.09 4.325 2.775 ;
 RECT 4.795 1.09 4.895 2.775 ;
 RECT 5.755 0.1 5.855 0.99 ;
 RECT 5.275 0.1 5.375 0.99 ;
 RECT 3.735 0.1 3.835 0.99 ;
 RECT 3.255 0.1 3.355 0.99 ;
 RECT 2.775 0.1 2.875 0.99 ;
 RECT 2.1 0.89 2.405 0.99 ;
 RECT 2.1 1.12 2.2 2.775 ;
 RECT 4.225 0.1 4.325 0.99 ;
 RECT 4.795 0.1 4.895 0.99 ;
 RECT 5.755 1.09 5.855 2.775 ;
 RECT 5.275 1.09 5.375 2.775 ;
 RECT 3.735 1.09 3.835 2.775 ;
 RECT 3.255 1.09 3.355 2.775 ;
 RECT 2.775 1.09 2.875 2.775 ;
 RECT 2.1 1.09 2.33 1.12 ;
 RECT 2.305 0.1 2.405 0.89 ;
 RECT 1.46 1.125 1.875 1.265 ;
 RECT 1.46 0.36 1.56 1.125 ;
 RECT 1.63 1.265 1.875 1.355 ;
 RECT 1.63 1.355 1.73 2.355 ;
 RECT 1.16 0.37 1.26 1.06 ;
 RECT 1.16 1.29 1.26 2.35 ;
 RECT 1.03 1.06 1.26 1.29 ;
 LAYER CO ;
 RECT 1.85 2.305 1.98 2.435 ;
 RECT 0.73 1.52 0.86 1.65 ;
 RECT 1.68 0.755 1.81 0.885 ;
 RECT 1.85 1.965 1.98 2.095 ;
 RECT 1.38 1.93 1.51 2.06 ;
 RECT 0.91 0.755 1.04 0.885 ;
 RECT 0.91 1.93 1.04 2.06 ;
 RECT 0.44 0.755 0.57 0.885 ;
 RECT 0.44 1.93 0.57 2.06 ;
 RECT 4.46 0.39 4.59 0.52 ;
 RECT 5.985 0.39 6.115 0.52 ;
 RECT 5.025 0.39 5.155 0.52 ;
 RECT 5.495 0.39 5.625 0.52 ;
 RECT 5.025 1.66 5.155 1.79 ;
 RECT 5.995 1.66 6.125 1.79 ;
 RECT 5.025 2.305 5.155 2.435 ;
 RECT 5.995 2.305 6.125 2.435 ;
 RECT 5.025 1.965 5.155 2.095 ;
 RECT 5.995 1.965 6.125 2.095 ;
 RECT 5.495 1.6 5.625 1.73 ;
 RECT 5.495 1.93 5.625 2.06 ;
 RECT 4.46 1.6 4.59 1.73 ;
 RECT 5.495 2.305 5.625 2.435 ;
 RECT 4.46 1.93 4.59 2.06 ;
 RECT 4.46 2.305 4.59 2.435 ;
 RECT 3.965 0.39 4.095 0.52 ;
 RECT 3.475 0.39 3.605 0.52 ;
 RECT 3.975 1.66 4.105 1.79 ;
 RECT 3.975 2.305 4.105 2.435 ;
 RECT 3.975 1.965 4.105 2.095 ;
 RECT 3.475 1.6 3.605 1.73 ;
 RECT 3.475 1.93 3.605 2.06 ;
 RECT 3.475 2.305 3.605 2.435 ;
 RECT 3.005 0.39 3.135 0.52 ;
 RECT 3.005 1.66 3.135 1.79 ;
 RECT 3.005 2.305 3.135 2.435 ;
 RECT 3.005 1.965 3.135 2.095 ;
 RECT 0.585 0.255 0.715 0.385 ;
 RECT 0.325 0.255 0.455 0.385 ;
 RECT 1.42 2.53 1.55 2.66 ;
 RECT 1.16 2.53 1.29 2.66 ;
 RECT 2.15 0.94 2.28 1.07 ;
 RECT 1.695 1.175 1.825 1.305 ;
 RECT 1.08 1.11 1.21 1.24 ;
 RECT 2.525 0.42 2.655 0.55 ;
 RECT 2.44 1.6 2.57 1.73 ;
 RECT 2.44 1.93 2.57 2.06 ;
 RECT 2.44 2.305 2.57 2.435 ;
 RECT 2.055 0.39 2.185 0.52 ;
 LAYER M1 ;
 RECT 0.435 0.645 0.575 1.105 ;
 RECT 0.435 1.245 0.575 2.11 ;
 RECT 1.075 1.04 1.215 1.105 ;
 RECT 1.075 1.245 1.215 1.3 ;
 RECT 0.435 1.105 1.215 1.245 ;
 RECT 1.375 0.89 1.515 2.11 ;
 RECT 2.08 0.89 2.33 1.075 ;
 RECT 1.375 0.75 2.33 0.89 ;
 RECT 2.145 1.075 2.285 1.09 ;
 END
END ISOLANDX8

MACRO ISOLORX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 RECT 1.72 1.9 1.86 2.8 ;
 RECT 0.35 1.945 0.49 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 RECT 0.725 0.565 0.975 0.705 ;
 RECT 1.66 0.565 1.925 0.705 ;
 RECT 0.35 0.08 0.49 0.765 ;
 RECT 0.77 0.08 0.91 0.565 ;
 RECT 1.725 0.08 1.865 0.565 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 1.15 1.24 1.485 ;
 END
 ANTENNAGATEAREA 0.111 ;
 END D

 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.435 1.15 1.85 1.425 ;
 END
 ANTENNAGATEAREA 0.111 ;
 END ISO

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.27 1.76 2.41 2.46 ;
 RECT 1.99 1.445 2.41 1.76 ;
 RECT 2.27 0.505 2.41 1.445 ;
 END
 ANTENNADIFFAREA 0.48 ;
 END Q

 OBS
 LAYER PO ;
 RECT 2.055 0.1 2.155 0.955 ;
 RECT 2.055 1.185 2.155 2.75 ;
 RECT 1.945 0.955 2.175 1.185 ;
 RECT 1.505 0.33 1.605 1.125 ;
 RECT 1.415 1.355 1.515 2.7 ;
 RECT 1.415 1.125 1.69 1.355 ;
 RECT 1.025 0.325 1.125 1.22 ;
 RECT 1.025 1.45 1.125 2.7 ;
 RECT 1.005 1.22 1.235 1.45 ;
 LAYER CO ;
 RECT 0.355 0.305 0.485 0.435 ;
 RECT 0.355 0.565 0.485 0.695 ;
 RECT 0.355 2.015 0.485 2.145 ;
 RECT 0.355 2.275 0.485 2.405 ;
 RECT 2.275 2.26 2.405 2.39 ;
 RECT 2.275 1.92 2.405 2.05 ;
 RECT 1.995 1.005 2.125 1.135 ;
 RECT 2.275 0.57 2.405 0.7 ;
 RECT 1.51 1.175 1.64 1.305 ;
 RECT 1.055 1.27 1.185 1.4 ;
 RECT 1.73 0.57 1.86 0.7 ;
 RECT 1.25 0.57 1.38 0.7 ;
 RECT 0.775 0.57 0.905 0.7 ;
 RECT 1.725 2.27 1.855 2.4 ;
 RECT 1.725 1.97 1.855 2.1 ;
 RECT 0.765 1.935 0.895 2.065 ;
 RECT 0.765 2.27 0.895 2.4 ;
 LAYER M1 ;
 RECT 0.67 0.87 0.81 1.64 ;
 RECT 0.67 1.64 0.9 1.86 ;
 RECT 0.755 1.86 0.9 2.005 ;
 RECT 0.76 2.005 0.9 2.47 ;
 RECT 1.245 0.565 1.385 0.995 ;
 RECT 0.76 0.87 1.385 1.01 ;
 RECT 1.18 0.565 1.45 0.705 ;
 RECT 1.99 0.87 2.13 1.205 ;
 RECT 1.355 0.87 2.125 1.01 ;
 END
END ISOLORX1

MACRO ISOLORX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 1.72 1.9 1.86 2.8 ;
 RECT 0.35 1.945 0.49 2.8 ;
 RECT 2.755 1.9 2.895 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 0.725 0.565 0.975 0.705 ;
 RECT 1.66 0.565 1.925 0.705 ;
 RECT 0.35 0.08 0.49 0.765 ;
 RECT 2.75 0.08 2.89 0.765 ;
 RECT 0.77 0.08 0.91 0.565 ;
 RECT 1.725 0.08 1.865 0.565 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.975 1.15 1.275 1.485 ;
 END
 ANTENNAGATEAREA 0.116 ;
 END D

 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.435 1.15 1.85 1.425 ;
 END
 ANTENNAGATEAREA 0.116 ;
 END ISO

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.27 1.72 2.41 2.46 ;
 RECT 1.99 1.48 2.41 1.72 ;
 RECT 2.27 0.505 2.41 1.48 ;
 END
 ANTENNADIFFAREA 0.6 ;
 END Q

 OBS
 LAYER PO ;
 RECT 1.945 0.955 2.63 1.035 ;
 RECT 2.53 1.035 2.63 2.75 ;
 RECT 2.055 0.1 2.155 0.935 ;
 RECT 2.055 0.935 2.63 0.955 ;
 RECT 2.53 0.1 2.63 0.935 ;
 RECT 1.945 1.035 2.175 1.185 ;
 RECT 2.055 1.185 2.155 2.75 ;
 RECT 1.505 0.33 1.605 1.125 ;
 RECT 1.415 1.355 1.515 2.7 ;
 RECT 1.415 1.125 1.69 1.355 ;
 RECT 1.025 0.325 1.125 1.22 ;
 RECT 1.025 1.45 1.125 2.7 ;
 RECT 1.005 1.22 1.235 1.45 ;
 LAYER CO ;
 RECT 2.755 0.57 2.885 0.7 ;
 RECT 2.76 2.27 2.89 2.4 ;
 RECT 2.76 1.97 2.89 2.1 ;
 RECT 0.355 0.305 0.485 0.435 ;
 RECT 0.355 0.565 0.485 0.695 ;
 RECT 0.355 2.015 0.485 2.145 ;
 RECT 0.355 2.275 0.485 2.405 ;
 RECT 2.275 2.26 2.405 2.39 ;
 RECT 2.275 1.92 2.405 2.05 ;
 RECT 1.995 1.005 2.125 1.135 ;
 RECT 2.275 0.57 2.405 0.7 ;
 RECT 1.51 1.175 1.64 1.305 ;
 RECT 1.055 1.27 1.185 1.4 ;
 RECT 1.73 0.57 1.86 0.7 ;
 RECT 1.25 0.57 1.38 0.7 ;
 RECT 0.775 0.57 0.905 0.7 ;
 RECT 1.725 2.27 1.855 2.4 ;
 RECT 1.725 1.97 1.855 2.1 ;
 RECT 0.765 1.935 0.895 2.065 ;
 RECT 0.765 2.27 0.895 2.4 ;
 LAYER M1 ;
 RECT 0.67 0.87 0.81 1.885 ;
 RECT 0.76 1.855 0.9 2.47 ;
 RECT 0.67 1.79 0.9 2.09 ;
 RECT 1.245 0.565 1.385 0.995 ;
 RECT 0.76 0.87 1.385 1.01 ;
 RECT 1.18 0.565 1.45 0.705 ;
 RECT 1.99 0.87 2.13 1.205 ;
 RECT 1.355 0.87 2.125 1.01 ;
 END
END ISOLORX2

MACRO ISOLORX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 1.72 1.9 1.86 2.8 ;
 RECT 0.35 1.945 0.49 2.8 ;
 RECT 2.755 1.9 2.895 2.8 ;
 RECT 3.715 1.9 3.855 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 0.725 0.565 0.975 0.705 ;
 RECT 1.66 0.565 1.925 0.705 ;
 RECT 0.35 0.08 0.49 0.765 ;
 RECT 2.75 0.08 2.89 0.765 ;
 RECT 3.71 0.08 3.85 0.765 ;
 RECT 0.77 0.08 0.91 0.565 ;
 RECT 1.725 0.08 1.865 0.565 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.97 1.15 1.275 1.485 ;
 END
 ANTENNAGATEAREA 0.111 ;
 END D

 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.435 1.15 1.85 1.63 ;
 END
 ANTENNAGATEAREA 0.111 ;
 END ISO

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.565 1.35 2.87 1.445 ;
 RECT 2.565 1.11 2.87 1.21 ;
 RECT 2.27 1.35 2.41 2.46 ;
 RECT 2.27 0.505 2.41 1.21 ;
 RECT 2.27 1.21 3.37 1.35 ;
 RECT 3.23 1.35 3.37 2.46 ;
 RECT 3.23 0.505 3.37 1.21 ;
 END
 ANTENNADIFFAREA 1.216 ;
 END Q

 OBS
 LAYER PO ;
 RECT 2.055 0.935 3.59 0.955 ;
 RECT 1.945 0.955 3.59 1.035 ;
 RECT 2.055 0.1 2.155 0.935 ;
 RECT 3.015 0.1 3.115 0.935 ;
 RECT 3.015 1.035 3.115 2.75 ;
 RECT 3.49 0.1 3.59 0.935 ;
 RECT 3.49 1.035 3.59 2.75 ;
 RECT 2.53 0.1 2.63 0.935 ;
 RECT 2.53 1.035 2.63 2.75 ;
 RECT 1.945 1.035 2.175 1.185 ;
 RECT 2.055 1.185 2.155 2.75 ;
 RECT 1.505 0.33 1.605 1.125 ;
 RECT 1.415 1.355 1.515 2.705 ;
 RECT 1.415 1.125 1.69 1.355 ;
 RECT 1.025 0.325 1.125 1.22 ;
 RECT 1.025 1.45 1.125 2.705 ;
 RECT 1.005 1.22 1.235 1.45 ;
 LAYER CO ;
 RECT 3.235 0.57 3.365 0.7 ;
 RECT 3.715 0.57 3.845 0.7 ;
 RECT 3.72 2.27 3.85 2.4 ;
 RECT 3.72 1.97 3.85 2.1 ;
 RECT 3.235 2.26 3.365 2.39 ;
 RECT 3.235 1.92 3.365 2.05 ;
 RECT 2.755 0.57 2.885 0.7 ;
 RECT 2.76 2.27 2.89 2.4 ;
 RECT 2.76 1.97 2.89 2.1 ;
 RECT 0.355 0.305 0.485 0.435 ;
 RECT 0.355 0.565 0.485 0.695 ;
 RECT 0.355 2.015 0.485 2.145 ;
 RECT 0.355 2.275 0.485 2.405 ;
 RECT 2.275 2.26 2.405 2.39 ;
 RECT 2.275 1.92 2.405 2.05 ;
 RECT 1.995 1.005 2.125 1.135 ;
 RECT 2.275 0.57 2.405 0.7 ;
 RECT 1.51 1.175 1.64 1.305 ;
 RECT 1.055 1.27 1.185 1.4 ;
 RECT 1.73 0.57 1.86 0.7 ;
 RECT 1.25 0.57 1.38 0.7 ;
 RECT 0.775 0.57 0.905 0.7 ;
 RECT 1.725 2.27 1.855 2.4 ;
 RECT 1.725 1.97 1.855 2.1 ;
 RECT 0.765 1.935 0.895 2.065 ;
 RECT 0.765 2.27 0.895 2.4 ;
 LAYER M1 ;
 RECT 0.64 0.87 0.78 1.94 ;
 RECT 0.76 1.855 0.9 2.47 ;
 RECT 0.64 1.74 0.9 2.02 ;
 RECT 1.245 0.565 1.385 0.995 ;
 RECT 0.76 0.87 1.385 1.01 ;
 RECT 1.18 0.565 1.45 0.705 ;
 RECT 1.99 0.87 2.13 1.205 ;
 RECT 1.355 0.87 2.125 1.01 ;
 END
END ISOLORX4

MACRO ISOLORX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.08 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.08 2.96 ;
 RECT 1.72 1.9 1.86 2.8 ;
 RECT 0.35 1.945 0.49 2.8 ;
 RECT 2.755 1.9 2.895 2.8 ;
 RECT 3.715 1.9 3.855 2.8 ;
 RECT 4.68 1.9 4.82 2.8 ;
 RECT 5.64 1.9 5.78 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.08 0.08 ;
 RECT 0.725 0.565 0.975 0.705 ;
 RECT 1.66 0.565 1.925 0.705 ;
 RECT 0.35 0.08 0.49 0.765 ;
 RECT 2.75 0.08 2.89 0.765 ;
 RECT 3.71 0.08 3.85 0.765 ;
 RECT 4.675 0.08 4.815 0.765 ;
 RECT 5.635 0.08 5.775 0.765 ;
 RECT 0.77 0.08 0.91 0.565 ;
 RECT 1.725 0.08 1.865 0.565 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.955 1.15 1.275 1.43 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END D

 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.435 1.15 1.85 1.425 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END ISO

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.52 1.35 3.825 1.425 ;
 RECT 3.52 1.11 3.825 1.21 ;
 RECT 3.23 1.35 3.37 2.46 ;
 RECT 3.23 0.505 3.37 1.21 ;
 RECT 4.195 1.35 4.335 2.46 ;
 RECT 4.195 0.505 4.335 1.21 ;
 RECT 5.155 1.35 5.295 2.46 ;
 RECT 5.155 0.505 5.295 1.21 ;
 RECT 2.27 1.35 2.41 2.46 ;
 RECT 2.27 0.505 2.41 1.21 ;
 RECT 2.27 1.21 5.295 1.35 ;
 END
 ANTENNADIFFAREA 2.432 ;
 END Q

 OBS
 LAYER PO ;
 RECT 1.025 0.345 1.125 1.14 ;
 RECT 1.025 1.37 1.125 2.755 ;
 RECT 1.005 1.14 1.235 1.37 ;
 RECT 2.055 0.935 5.515 0.955 ;
 RECT 1.945 0.955 5.515 1.035 ;
 RECT 2.055 0.15 2.155 0.935 ;
 RECT 4.94 0.15 5.04 0.935 ;
 RECT 4.94 1.035 5.04 2.75 ;
 RECT 5.415 0.15 5.515 0.935 ;
 RECT 5.415 1.035 5.515 2.75 ;
 RECT 4.455 0.15 4.555 0.935 ;
 RECT 4.455 1.035 4.555 2.75 ;
 RECT 3.98 0.15 4.08 0.935 ;
 RECT 3.98 1.035 4.08 2.75 ;
 RECT 3.015 0.15 3.115 0.935 ;
 RECT 3.015 1.035 3.115 2.75 ;
 RECT 3.49 0.15 3.59 0.935 ;
 RECT 3.49 1.035 3.59 2.75 ;
 RECT 2.53 0.15 2.63 0.935 ;
 RECT 2.53 1.035 2.63 2.75 ;
 RECT 1.945 1.035 2.175 1.185 ;
 RECT 2.055 1.185 2.155 2.75 ;
 RECT 1.505 0.345 1.605 1.125 ;
 RECT 1.415 1.355 1.515 2.755 ;
 RECT 1.415 1.125 1.69 1.355 ;
 LAYER CO ;
 RECT 1.055 1.19 1.185 1.32 ;
 RECT 5.645 1.97 5.775 2.1 ;
 RECT 5.16 2.26 5.29 2.39 ;
 RECT 4.2 0.57 4.33 0.7 ;
 RECT 5.16 1.92 5.29 2.05 ;
 RECT 4.68 0.57 4.81 0.7 ;
 RECT 4.685 2.27 4.815 2.4 ;
 RECT 4.685 1.97 4.815 2.1 ;
 RECT 5.16 0.57 5.29 0.7 ;
 RECT 4.2 2.26 4.33 2.39 ;
 RECT 5.64 0.57 5.77 0.7 ;
 RECT 4.2 1.92 4.33 2.05 ;
 RECT 5.645 2.27 5.775 2.4 ;
 RECT 3.235 0.57 3.365 0.7 ;
 RECT 3.715 0.57 3.845 0.7 ;
 RECT 3.72 2.27 3.85 2.4 ;
 RECT 3.72 1.97 3.85 2.1 ;
 RECT 3.235 2.26 3.365 2.39 ;
 RECT 3.235 1.92 3.365 2.05 ;
 RECT 2.755 0.57 2.885 0.7 ;
 RECT 2.76 2.27 2.89 2.4 ;
 RECT 2.76 1.97 2.89 2.1 ;
 RECT 0.355 0.305 0.485 0.435 ;
 RECT 0.355 0.565 0.485 0.695 ;
 RECT 0.355 2.015 0.485 2.145 ;
 RECT 0.355 2.275 0.485 2.405 ;
 RECT 2.275 2.26 2.405 2.39 ;
 RECT 2.275 1.92 2.405 2.05 ;
 RECT 1.995 1.005 2.125 1.135 ;
 RECT 2.275 0.57 2.405 0.7 ;
 RECT 1.51 1.175 1.64 1.305 ;
 RECT 1.73 0.57 1.86 0.7 ;
 RECT 1.25 0.57 1.38 0.7 ;
 RECT 0.775 0.57 0.905 0.7 ;
 RECT 1.725 2.27 1.855 2.4 ;
 RECT 1.725 1.97 1.855 2.1 ;
 RECT 0.765 1.935 0.895 2.065 ;
 RECT 0.765 2.27 0.895 2.4 ;
 LAYER M1 ;
 RECT 0.64 0.87 0.78 1.875 ;
 RECT 0.76 1.855 0.9 2.47 ;
 RECT 0.635 1.715 0.9 1.99 ;
 RECT 1.245 0.565 1.385 0.995 ;
 RECT 0.76 0.87 1.385 1.01 ;
 RECT 1.18 0.565 1.45 0.705 ;
 RECT 1.99 0.87 2.13 1.205 ;
 RECT 1.355 0.87 2.125 1.01 ;
 END
END ISOLORX8

MACRO RDFFNSRASX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 30.08 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 23.045 0.59 23.415 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 28.275 1.435 28.615 1.8 ;
 RECT 26.595 1.99 28.46 2.13 ;
 RECT 24.365 2.22 26.735 2.36 ;
 RECT 26.595 1.435 26.735 1.99 ;
 RECT 28.32 1.8 28.46 1.99 ;
 RECT 24.365 1.39 24.505 2.22 ;
 RECT 25.75 1.37 25.89 2.22 ;
 RECT 26.595 2.13 26.735 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.84 2.12 1.165 2.59 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.825 0.08 2.105 0.295 ;
 RECT 26.715 0.08 26.955 0.26 ;
 RECT 5.755 0.31 6.045 0.45 ;
 RECT 9.44 0.615 9.71 0.755 ;
 RECT 13.365 0.275 14.39 0.415 ;
 RECT 19.03 0.29 19.27 0.45 ;
 RECT 18.045 0.335 18.31 0.495 ;
 RECT 14.25 0.75 15.195 0.89 ;
 RECT 0 -0.08 30.08 0.08 ;
 RECT 1.305 0.08 1.445 0.97 ;
 RECT 0.335 0.08 0.475 0.775 ;
 RECT 4.65 0.08 4.885 0.46 ;
 RECT 20.565 0.08 20.705 0.325 ;
 RECT 21.63 0.08 21.77 0.82 ;
 RECT 24.365 0.08 24.505 0.36 ;
 RECT 25.58 0.08 25.72 0.35 ;
 RECT 5.835 0.08 5.975 0.31 ;
 RECT 9.505 0.08 9.645 0.615 ;
 RECT 13.365 0.415 13.505 0.945 ;
 RECT 13.365 0.08 13.505 0.275 ;
 RECT 19.085 0.08 19.225 0.29 ;
 RECT 18.1 0.08 18.24 0.335 ;
 RECT 15.055 0.89 15.195 1.11 ;
 RECT 14.25 0.415 14.39 0.75 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 9.25 2.215 9.525 2.355 ;
 RECT 0 2.8 30.08 2.96 ;
 RECT 1.98 2.34 2.23 2.8 ;
 RECT 0.335 1.74 0.475 2.8 ;
 RECT 1.305 1.98 1.445 2.8 ;
 RECT 6.865 2 7.005 2.8 ;
 RECT 5.835 1.98 5.975 2.8 ;
 RECT 12.275 2.335 12.545 2.8 ;
 RECT 20.48 2.57 20.62 2.8 ;
 RECT 19.02 2.57 19.16 2.8 ;
 RECT 18.015 2.57 18.155 2.8 ;
 RECT 21.545 2.57 21.685 2.8 ;
 RECT 5.355 2.65 5.495 2.8 ;
 RECT 5.355 2.44 5.69 2.65 ;
 RECT 5.355 2.07 5.495 2.44 ;
 RECT 9.315 2.355 9.455 2.8 ;
 RECT 9.315 2.195 9.455 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 1.475 1.605 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.73 2.255 10.04 2.465 ;
 RECT 9.8 2.465 10.04 2.47 ;
 RECT 9.8 2.12 10.04 2.255 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.24 1.795 7.48 2.04 ;
 RECT 6.655 1.795 6.885 1.83 ;
 RECT 6.655 1.655 7.48 1.795 ;
 RECT 6.655 1.62 6.885 1.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.48 1.16 17.75 1.445 ;
 RECT 17.61 0.915 17.75 1.16 ;
 RECT 18.615 1.84 18.755 1.885 ;
 RECT 18.615 0.915 18.755 1.7 ;
 RECT 19.555 1.84 19.695 1.885 ;
 RECT 19.555 0.915 19.695 1.7 ;
 RECT 17.61 1.7 19.695 1.84 ;
 RECT 17.61 1.84 17.75 1.885 ;
 RECT 17.61 1.445 17.75 1.7 ;
 END
 ANTENNADIFFAREA 1.165 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 21.065 1.905 21.205 1.91 ;
 RECT 21.065 0.56 21.205 1.765 ;
 RECT 22.13 1.905 22.27 1.91 ;
 RECT 22.13 0.56 22.27 1.765 ;
 RECT 20.005 0.51 20.145 1.48 ;
 RECT 20.005 1.48 20.285 1.765 ;
 RECT 20.005 1.765 22.27 1.905 ;
 END
 ANTENNADIFFAREA 0.909 ;
 END Q

 OBS
 LAYER PO ;
 RECT 12.09 1.39 12.285 1.405 ;
 RECT 3.225 1.565 3.325 2.675 ;
 RECT 2.34 1.62 2.44 2.675 ;
 RECT 1.905 1.44 2.15 1.52 ;
 RECT 1.905 1.62 2.15 1.69 ;
 RECT 4.46 0.285 4.56 1.24 ;
 RECT 11.195 1.29 12.285 1.39 ;
 RECT 2.34 2.675 3.325 2.775 ;
 RECT 12.09 1.405 12.32 1.615 ;
 RECT 24.625 1.245 24.725 2.02 ;
 RECT 24.495 1.035 24.725 1.245 ;
 RECT 12.585 0.105 15.41 0.205 ;
 RECT 12.585 0.205 12.685 1.91 ;
 RECT 15.31 0.205 15.41 1.265 ;
 RECT 11.765 1.71 11.865 1.91 ;
 RECT 10.68 1.61 11.865 1.71 ;
 RECT 10.68 0.475 10.78 1.61 ;
 RECT 11.23 1.71 11.33 2.425 ;
 RECT 7.345 0.475 7.445 0.895 ;
 RECT 11.765 1.91 12.685 2.01 ;
 RECT 7.345 0.375 10.78 0.475 ;
 RECT 7.22 0.895 7.45 1.105 ;
 RECT 12.895 0.455 14.825 0.535 ;
 RECT 14.595 0.535 14.825 0.6 ;
 RECT 14.595 0.39 14.825 0.435 ;
 RECT 12.975 0.435 14.825 0.455 ;
 RECT 12.895 0.535 13.125 0.665 ;
 RECT 13.75 0.535 13.98 0.835 ;
 RECT 13.75 0.835 13.85 2.39 ;
 RECT 24.93 0.215 25.03 0.995 ;
 RECT 24.93 0.995 25.17 1.205 ;
 RECT 24.93 1.205 25.03 2 ;
 RECT 27.325 0.375 27.425 0.99 ;
 RECT 27.325 0.99 27.575 1.2 ;
 RECT 27.325 1.2 27.425 2.27 ;
 RECT 27.325 2.27 27.61 2.48 ;
 RECT 10.16 0.655 10.26 2.305 ;
 RECT 10.465 2.3 10.695 2.305 ;
 RECT 10.465 2.405 10.695 2.51 ;
 RECT 10.16 2.305 10.695 2.405 ;
 RECT 24.15 0.21 24.25 0.755 ;
 RECT 24.15 0.855 24.25 2.2 ;
 RECT 27.015 1.125 27.115 2.2 ;
 RECT 23.185 0.755 24.72 0.84 ;
 RECT 23.185 0.84 24.715 0.855 ;
 RECT 24.62 0.215 24.72 0.755 ;
 RECT 23.185 0.595 23.415 0.755 ;
 RECT 24.15 2.2 27.115 2.3 ;
 RECT 25.84 1.06 25.94 1.14 ;
 RECT 25.84 0.38 25.94 0.96 ;
 RECT 25.84 1.14 26.11 1.24 ;
 RECT 26.01 1.24 26.11 1.84 ;
 RECT 25.42 0.935 25.65 0.96 ;
 RECT 25.42 0.96 25.94 1.06 ;
 RECT 25.42 1.06 25.65 1.145 ;
 RECT 26.205 0.22 26.435 0.28 ;
 RECT 26.205 0.38 26.435 0.43 ;
 RECT 25.84 0.28 26.435 0.38 ;
 RECT 7.945 1.575 8.045 2.485 ;
 RECT 8.455 1.575 8.685 1.685 ;
 RECT 7.945 1.475 8.685 1.575 ;
 RECT 28.025 0.195 28.125 2.665 ;
 RECT 27.015 0.095 28.125 0.195 ;
 RECT 23.39 1.245 23.49 2.665 ;
 RECT 23.39 1.2 23.675 1.245 ;
 RECT 27.015 0.195 27.115 0.945 ;
 RECT 23.445 1.035 23.675 1.1 ;
 RECT 23.39 2.665 28.125 2.765 ;
 RECT 23.39 1.1 23.72 1.2 ;
 RECT 12.17 0.795 12.335 0.925 ;
 RECT 11.49 0.885 11.72 0.925 ;
 RECT 11.49 1.025 11.72 1.095 ;
 RECT 11.49 0.925 12.335 1.025 ;
 RECT 12.17 0.585 12.4 0.795 ;
 RECT 9.765 0.655 9.865 1.24 ;
 RECT 9.155 1.34 9.385 1.475 ;
 RECT 9.155 1.24 9.865 1.34 ;
 RECT 1.565 0.49 1.665 1.495 ;
 RECT 1.37 1.495 1.665 1.745 ;
 RECT 1.565 1.745 1.665 2.37 ;
 RECT 3.72 1.33 3.86 1.475 ;
 RECT 3.72 1.71 3.82 2.475 ;
 RECT 3.76 0.65 3.86 1.33 ;
 RECT 3.72 1.475 3.95 1.71 ;
 RECT 4.16 0.715 4.26 1.61 ;
 RECT 4.195 1.71 4.295 2.48 ;
 RECT 4.16 1.61 4.295 1.71 ;
 RECT 4.04 0.485 4.28 0.715 ;
 RECT 3.27 0.705 3.37 1.165 ;
 RECT 2.83 1.27 2.93 1.445 ;
 RECT 3.27 0.47 3.555 0.705 ;
 RECT 2.83 1.17 3.37 1.265 ;
 RECT 3.06 1.165 3.37 1.17 ;
 RECT 2.83 1.265 3.205 1.27 ;
 RECT 2.685 1.445 2.93 1.69 ;
 RECT 0.93 2.37 1.19 2.58 ;
 RECT 1.09 0.27 1.19 2.37 ;
 RECT 8.87 0.655 8.97 1.18 ;
 RECT 8.87 1.28 8.97 1.655 ;
 RECT 7.955 0.66 8.055 1.18 ;
 RECT 8.87 1.655 9.83 1.755 ;
 RECT 9.73 1.755 9.83 2.255 ;
 RECT 8.87 1.755 8.97 2.51 ;
 RECT 7.955 1.18 8.97 1.28 ;
 RECT 9.73 2.255 9.96 2.465 ;
 RECT 5.615 0.745 5.715 2.44 ;
 RECT 5.46 2.44 5.715 2.65 ;
 RECT 5.325 0.535 5.555 0.645 ;
 RECT 5.325 0.645 5.715 0.745 ;
 RECT 16.19 0.77 16.29 2.155 ;
 RECT 16.19 0.55 16.29 0.56 ;
 RECT 16.19 0.56 16.445 0.77 ;
 RECT 17.875 0.39 17.975 1.4 ;
 RECT 17.875 1.5 17.975 2.37 ;
 RECT 16.825 0.43 16.925 1.245 ;
 RECT 16.76 0.29 17.975 0.39 ;
 RECT 19.34 0.51 19.44 1.4 ;
 RECT 19.34 1.5 19.44 2.37 ;
 RECT 18.87 0.515 18.97 1.4 ;
 RECT 18.87 1.5 18.97 2.37 ;
 RECT 17.875 1.4 19.44 1.5 ;
 RECT 18.365 0.51 18.465 1.4 ;
 RECT 18.365 1.5 18.465 2.37 ;
 RECT 16.76 0.22 16.99 0.29 ;
 RECT 16.76 0.39 16.99 0.43 ;
 RECT 16.775 1.245 17.005 1.455 ;
 RECT 4.98 2.445 5.24 2.655 ;
 RECT 5.14 1.79 5.24 2.445 ;
 RECT 15.25 1.445 15.35 2.035 ;
 RECT 15.235 2.035 15.465 2.245 ;
 RECT 15.72 0.55 15.82 2.69 ;
 RECT 6.65 1.83 6.75 2.69 ;
 RECT 6.65 1.58 6.75 1.62 ;
 RECT 6.39 1.01 6.49 1.48 ;
 RECT 6.65 1.62 6.885 1.83 ;
 RECT 6.65 2.69 15.82 2.79 ;
 RECT 6.39 1.48 6.75 1.58 ;
 RECT 6.09 0.98 6.19 1.615 ;
 RECT 5.95 1.615 6.19 1.825 ;
 RECT 6.09 1.825 6.19 2.51 ;
 RECT 20.725 1.195 20.945 1.33 ;
 RECT 20.845 0.385 20.945 1.195 ;
 RECT 20.265 1.33 22.01 1.43 ;
 RECT 20.845 1.43 20.945 2.575 ;
 RECT 21.91 0.195 22.01 1.33 ;
 RECT 20.265 0.385 20.365 1.33 ;
 RECT 20.265 1.43 20.365 2.575 ;
 RECT 21.33 0.385 21.43 1.33 ;
 RECT 21.33 1.43 21.43 2.575 ;
 RECT 21.91 1.43 22.01 2.575 ;
 RECT 21.91 0.095 22.505 0.195 ;
 RECT 22.405 0.195 22.505 0.22 ;
 RECT 22.405 0.22 22.635 0.43 ;
 RECT 14.22 0.73 14.32 1.39 ;
 RECT 14.085 1.39 14.32 1.6 ;
 RECT 14.22 1.6 14.32 2.39 ;
 RECT 2.405 0.285 2.505 1.52 ;
 RECT 1.905 1.52 2.505 1.62 ;
 RECT 2.405 0.185 11.295 0.195 ;
 RECT 4.46 0.095 11.295 0.185 ;
 RECT 2.405 0.195 4.56 0.285 ;
 RECT 11.195 0.195 11.295 1.29 ;
 LAYER CO ;
 RECT 11.45 1.87 11.58 2 ;
 RECT 0.34 0.59 0.47 0.72 ;
 RECT 9.205 1.28 9.335 1.41 ;
 RECT 3.375 0.525 3.505 0.655 ;
 RECT 8.62 1.995 8.75 2.125 ;
 RECT 4.89 2.11 5.02 2.24 ;
 RECT 8.175 2.07 8.305 2.2 ;
 RECT 1.965 1.495 2.095 1.625 ;
 RECT 1.915 0.745 2.045 0.875 ;
 RECT 0.98 2.41 1.11 2.54 ;
 RECT 9.78 2.295 9.91 2.425 ;
 RECT 5.51 2.48 5.64 2.61 ;
 RECT 5.375 0.575 5.505 0.705 ;
 RECT 16.825 1.285 16.955 1.415 ;
 RECT 14.645 0.43 14.775 0.56 ;
 RECT 16.265 0.6 16.395 0.73 ;
 RECT 16.81 0.26 16.94 0.39 ;
 RECT 5.03 2.485 5.16 2.615 ;
 RECT 15.285 2.075 15.415 2.205 ;
 RECT 6.705 1.66 6.835 1.79 ;
 RECT 6 1.655 6.13 1.785 ;
 RECT 22.455 0.26 22.585 0.39 ;
 RECT 27.395 1.03 27.525 1.16 ;
 RECT 12.945 0.495 13.075 0.625 ;
 RECT 14.135 1.43 14.265 1.56 ;
 RECT 12.22 0.625 12.35 0.755 ;
 RECT 12.14 1.445 12.27 1.575 ;
 RECT 24.545 1.075 24.675 1.205 ;
 RECT 7.27 0.935 7.4 1.065 ;
 RECT 25.47 0.975 25.6 1.105 ;
 RECT 13.8 0.665 13.93 0.795 ;
 RECT 24.99 1.035 25.12 1.165 ;
 RECT 27.43 2.31 27.56 2.44 ;
 RECT 10.515 2.34 10.645 2.47 ;
 RECT 23.235 0.635 23.365 0.765 ;
 RECT 26.255 0.26 26.385 0.39 ;
 RECT 8.505 1.515 8.635 1.645 ;
 RECT 23.495 1.075 23.625 1.205 ;
 RECT 11.54 0.925 11.67 1.055 ;
 RECT 10.945 1.9 11.075 2.03 ;
 RECT 16.415 1.705 16.545 1.835 ;
 RECT 15.06 0.91 15.19 1.04 ;
 RECT 26.23 1.405 26.36 1.535 ;
 RECT 15.47 1.705 15.6 1.835 ;
 RECT 8.175 0.905 8.305 1.035 ;
 RECT 3.94 2.11 4.07 2.24 ;
 RECT 9.51 0.62 9.64 0.75 ;
 RECT 0.34 2.345 0.47 2.475 ;
 RECT 0.34 1.825 0.47 1.955 ;
 RECT 13.5 1.835 13.63 1.965 ;
 RECT 2.05 2.345 2.18 2.475 ;
 RECT 6.65 1.23 6.78 1.36 ;
 RECT 0.34 0.33 0.47 0.46 ;
 RECT 1.31 0.74 1.44 0.87 ;
 RECT 5.84 2.075 5.97 2.205 ;
 RECT 2.625 0.79 2.755 0.92 ;
 RECT 28.325 1.475 28.455 1.605 ;
 RECT 18.105 0.36 18.235 0.49 ;
 RECT 21.55 2.64 21.68 2.77 ;
 RECT 20.57 0.12 20.7 0.25 ;
 RECT 19.56 0.975 19.69 1.105 ;
 RECT 18.62 1.705 18.75 1.835 ;
 RECT 18.02 2.64 18.15 2.77 ;
 RECT 20.01 1.725 20.14 1.855 ;
 RECT 21.635 0.62 21.765 0.75 ;
 RECT 19.09 0.315 19.22 0.445 ;
 RECT 18.62 0.975 18.75 1.105 ;
 RECT 21.07 0.63 21.2 0.76 ;
 RECT 22.135 0.63 22.265 0.76 ;
 RECT 21.07 1.71 21.2 1.84 ;
 RECT 17.615 0.975 17.745 1.105 ;
 RECT 19.025 2.64 19.155 2.77 ;
 RECT 20.485 2.64 20.615 2.77 ;
 RECT 17.615 1.705 17.745 1.835 ;
 RECT 22.135 1.71 22.265 1.84 ;
 RECT 20.765 1.245 20.895 1.375 ;
 RECT 19.56 1.705 19.69 1.835 ;
 RECT 20.01 0.62 20.14 0.75 ;
 RECT 0.34 2.085 0.47 2.215 ;
 RECT 6.38 2.045 6.51 2.175 ;
 RECT 1.43 1.55 1.56 1.68 ;
 RECT 14.475 1.035 14.605 1.165 ;
 RECT 7.7 0.905 7.83 1.035 ;
 RECT 11.45 0.595 11.58 0.725 ;
 RECT 25.755 1.445 25.885 1.575 ;
 RECT 6.87 2.11 7 2.24 ;
 RECT 5.84 0.315 5.97 0.445 ;
 RECT 2.975 2.105 3.105 2.235 ;
 RECT 3.49 0.88 3.62 1.01 ;
 RECT 16.535 0.92 16.665 1.05 ;
 RECT 5.36 2.135 5.49 2.265 ;
 RECT 26.765 0.12 26.895 0.25 ;
 RECT 1.895 0.145 2.025 0.275 ;
 RECT 25.15 0.435 25.28 0.565 ;
 RECT 8.62 0.905 8.75 1.035 ;
 RECT 0.84 0.74 0.97 0.87 ;
 RECT 4.095 0.53 4.225 0.66 ;
 RECT 25.585 0.12 25.715 0.25 ;
 RECT 2.56 1.825 2.69 1.955 ;
 RECT 9.32 2.225 9.45 2.355 ;
 RECT 0.84 1.665 0.97 1.795 ;
 RECT 24.37 1.475 24.5 1.605 ;
 RECT 14.44 1.835 14.57 1.965 ;
 RECT 27.545 1.465 27.675 1.595 ;
 RECT 12.345 2.38 12.475 2.51 ;
 RECT 23.9 1.425 24.03 1.555 ;
 RECT 13.37 0.765 13.5 0.895 ;
 RECT 23.65 0.505 23.78 0.635 ;
 RECT 10.42 0.875 10.55 1.005 ;
 RECT 25.15 1.485 25.28 1.615 ;
 RECT 3.47 2.07 3.6 2.2 ;
 RECT 15.94 1.705 16.07 1.835 ;
 RECT 4.42 1.825 4.55 1.955 ;
 RECT 10.42 1.945 10.55 2.075 ;
 RECT 26.6 1.49 26.73 1.62 ;
 RECT 7.695 2.015 7.825 2.145 ;
 RECT 4.705 0.32 4.835 0.45 ;
 RECT 26.09 0.595 26.22 0.725 ;
 RECT 27.545 0.595 27.675 0.725 ;
 RECT 10.945 0.595 11.075 0.725 ;
 RECT 1.785 1.995 1.915 2.125 ;
 RECT 1.31 2.05 1.44 2.18 ;
 RECT 3.02 0.88 3.15 1.01 ;
 RECT 24.37 0.135 24.5 0.265 ;
 RECT 3.77 1.525 3.9 1.655 ;
 RECT 2.74 1.49 2.87 1.62 ;
 LAYER M1 ;
 RECT 23.585 1.015 23.895 1.035 ;
 RECT 23.445 1.035 23.895 1.055 ;
 RECT 23.72 0.64 23.86 1.015 ;
 RECT 23.895 1.225 24.035 1.75 ;
 RECT 23.6 0.5 23.86 0.64 ;
 RECT 24.495 1.035 24.725 1.055 ;
 RECT 24.495 1.195 24.725 1.245 ;
 RECT 23.445 1.055 24.725 1.195 ;
 RECT 25.465 1.145 25.605 1.345 ;
 RECT 25.145 1.485 25.285 1.76 ;
 RECT 25.465 0.73 25.605 0.935 ;
 RECT 25.145 0.355 25.285 0.59 ;
 RECT 25.145 1.345 25.605 1.485 ;
 RECT 25.42 0.935 25.65 1.145 ;
 RECT 25.145 0.59 25.605 0.73 ;
 RECT 22.405 0.36 22.635 0.43 ;
 RECT 24 0.36 24.14 0.565 ;
 RECT 22.405 0.22 24.14 0.36 ;
 RECT 24.74 0.705 24.88 0.75 ;
 RECT 24.865 0.995 25.17 1.205 ;
 RECT 24.865 0.89 25.005 0.995 ;
 RECT 24.74 0.75 25.005 0.89 ;
 RECT 24 0.565 24.88 0.705 ;
 RECT 13.75 0.57 13.98 0.95 ;
 RECT 16.76 0.22 16.99 0.28 ;
 RECT 16.76 0.42 16.99 0.43 ;
 RECT 14.595 0.28 16.99 0.42 ;
 RECT 14.595 0.42 14.825 0.6 ;
 RECT 15.49 0.775 15.63 1.405 ;
 RECT 16.215 0.56 16.445 0.635 ;
 RECT 14.47 1.405 15.63 1.545 ;
 RECT 14.47 1.545 14.61 1.83 ;
 RECT 13.425 1.83 14.675 1.97 ;
 RECT 14.47 1.17 14.61 1.405 ;
 RECT 14.4 1.03 14.68 1.17 ;
 RECT 19.605 0.36 19.745 0.635 ;
 RECT 15.49 0.635 19.745 0.775 ;
 RECT 20.285 0.36 20.425 0.68 ;
 RECT 19.605 0.22 20.425 0.36 ;
 RECT 20.76 0.675 20.9 0.68 ;
 RECT 20.76 0.82 20.9 1.445 ;
 RECT 20.285 0.68 20.9 0.82 ;
 RECT 12.17 0.585 13.125 0.63 ;
 RECT 12.895 0.63 13.125 0.665 ;
 RECT 12.895 0.455 13.125 0.49 ;
 RECT 12.195 0.49 13.125 0.585 ;
 RECT 12.17 0.63 12.4 0.795 ;
 RECT 11.445 0.525 11.585 0.885 ;
 RECT 11.445 1.095 11.585 2.065 ;
 RECT 11.445 0.885 11.72 1.095 ;
 RECT 8.17 1.04 8.31 2.34 ;
 RECT 8.17 0.895 8.31 0.9 ;
 RECT 8.965 2.055 9.105 2.34 ;
 RECT 8.1 0.9 8.375 1.04 ;
 RECT 8.17 2.34 9.105 2.48 ;
 RECT 9.49 1.66 9.63 1.915 ;
 RECT 8.965 1.915 9.63 2.055 ;
 RECT 9.49 1.52 11.08 1.66 ;
 RECT 10.415 0.765 10.555 1.52 ;
 RECT 10.415 1.66 10.555 2.145 ;
 RECT 10.94 0.525 11.08 1.52 ;
 RECT 10.94 1.66 11.08 2.11 ;
 RECT 3.765 0.895 7.45 1.035 ;
 RECT 7.22 1.035 7.45 1.105 ;
 RECT 3.305 0.52 3.905 0.66 ;
 RECT 3.765 0.66 3.905 0.895 ;
 RECT 3.31 1.82 4.89 1.96 ;
 RECT 4.75 1.79 4.89 1.82 ;
 RECT 3.395 1.96 3.675 2.215 ;
 RECT 3.485 0.805 3.625 1.22 ;
 RECT 3.31 1.22 3.625 1.36 ;
 RECT 3.31 1.36 3.45 1.82 ;
 RECT 5.95 1.615 6.18 1.65 ;
 RECT 5.95 1.79 6.18 1.825 ;
 RECT 4.75 1.65 6.185 1.79 ;
 RECT 13.74 1.23 13.88 1.42 ;
 RECT 11.89 1.09 13.88 1.23 ;
 RECT 11.89 0.385 12.03 1.09 ;
 RECT 9.88 0.385 10.02 0.895 ;
 RECT 9.875 0.255 12.03 0.385 ;
 RECT 9.875 0.245 12.025 0.255 ;
 RECT 8.965 0.895 10.02 1.035 ;
 RECT 8.965 0.745 9.105 0.895 ;
 RECT 4.045 0.605 9.105 0.745 ;
 RECT 5.325 0.535 5.555 0.605 ;
 RECT 4.045 0.485 4.36 0.605 ;
 RECT 14.085 1.39 14.315 1.42 ;
 RECT 13.74 1.42 14.315 1.56 ;
 RECT 14.085 1.56 14.315 1.6 ;
 RECT 0.615 1.335 0.755 1.66 ;
 RECT 0.615 0.875 0.755 1.195 ;
 RECT 0.615 1.66 1.02 1.8 ;
 RECT 0.615 0.735 1.04 0.875 ;
 RECT 0.615 1.195 1.725 1.335 ;
 RECT 1.585 0.6 1.725 1.195 ;
 RECT 3.015 0.36 3.155 2.035 ;
 RECT 2.33 0.22 3.155 0.36 ;
 RECT 2.33 0.36 2.47 0.46 ;
 RECT 2.97 2.17 3.11 2.305 ;
 RECT 2.97 2.035 3.155 2.17 ;
 RECT 1.585 0.46 2.47 0.6 ;
 RECT 1.865 0.88 2.005 1.475 ;
 RECT 1.825 1.63 1.965 1.99 ;
 RECT 1.825 1.475 2.17 1.63 ;
 RECT 1.715 1.99 1.965 2.13 ;
 RECT 1.865 0.74 2.185 0.88 ;
 RECT 2.62 1.67 2.76 1.82 ;
 RECT 2.62 1.96 2.76 2.51 ;
 RECT 4.98 2.445 5.21 2.51 ;
 RECT 4.98 2.65 5.21 2.655 ;
 RECT 2.62 0.5 2.76 1.44 ;
 RECT 2.62 1.44 2.875 1.67 ;
 RECT 2.49 1.82 2.76 1.96 ;
 RECT 2.62 2.51 5.21 2.65 ;
 RECT 12.86 1.895 13 2.39 ;
 RECT 17.005 2.205 17.145 2.39 ;
 RECT 12.86 2.39 17.145 2.53 ;
 RECT 11.735 1.755 13 1.895 ;
 RECT 11.735 1.895 11.875 2.34 ;
 RECT 10.465 2.3 10.695 2.34 ;
 RECT 10.465 2.48 10.695 2.51 ;
 RECT 10.465 2.34 11.875 2.48 ;
 RECT 17.005 2.065 23.18 2.205 ;
 RECT 23.04 2.205 23.18 2.52 ;
 RECT 27.38 2.48 27.52 2.52 ;
 RECT 23.04 2.52 27.52 2.66 ;
 RECT 27.38 2.27 27.61 2.48 ;
 RECT 15.41 1.7 15.745 1.84 ;
 RECT 15.605 1.84 15.745 2.075 ;
 RECT 16.3 1.84 16.44 2.075 ;
 RECT 16.3 1.7 16.595 1.84 ;
 RECT 15.605 2.075 16.44 2.215 ;
 RECT 15.935 1.385 16.075 1.625 ;
 RECT 16.495 1.055 16.635 1.245 ;
 RECT 15.935 1.245 17.005 1.385 ;
 RECT 16.775 1.385 17.005 1.455 ;
 RECT 16.465 0.915 16.765 1.055 ;
 RECT 15.905 1.625 16.16 1.92 ;
 RECT 13.14 1.56 13.28 2.11 ;
 RECT 12.09 1.405 12.32 1.42 ;
 RECT 12.09 1.42 13.28 1.56 ;
 RECT 12.09 1.56 12.32 1.615 ;
 RECT 13.14 2.11 15.465 2.245 ;
 RECT 15.235 2.035 15.465 2.11 ;
 RECT 13.14 2.245 15.46 2.25 ;
 RECT 8.615 1.685 9.34 1.775 ;
 RECT 8.615 1.775 8.755 2.18 ;
 RECT 8.455 1.635 9.34 1.685 ;
 RECT 9.2 1.205 9.34 1.635 ;
 RECT 8.615 1.04 8.755 1.475 ;
 RECT 8.455 1.475 8.755 1.635 ;
 RECT 8.545 0.9 8.82 1.04 ;
 RECT 3.87 2.105 5.09 2.245 ;
 RECT 4.43 1.225 7.08 1.25 ;
 RECT 6.375 1.365 6.515 2.25 ;
 RECT 4.43 1.365 4.57 1.5 ;
 RECT 3.6 1.64 4.105 1.675 ;
 RECT 3.6 1.5 4.57 1.64 ;
 RECT 7.69 1.04 7.83 1.25 ;
 RECT 7.69 1.39 7.83 2.215 ;
 RECT 7.69 0.885 7.83 0.9 ;
 RECT 4.43 1.25 7.83 1.365 ;
 RECT 6.94 1.365 7.83 1.39 ;
 RECT 7.625 0.9 7.9 1.04 ;
 RECT 26.085 0.73 26.225 1.04 ;
 RECT 26.225 1.18 26.365 1.605 ;
 RECT 26.02 0.59 26.295 0.73 ;
 RECT 27.345 0.99 27.575 1.04 ;
 RECT 26.085 1.04 27.575 1.18 ;
 RECT 27.345 1.18 27.575 1.2 ;
 RECT 26.205 0.29 26.575 0.43 ;
 RECT 26.435 0.43 26.575 0.71 ;
 RECT 26.205 0.22 26.435 0.29 ;
 RECT 27.855 0.85 27.995 1.385 ;
 RECT 27.54 1.525 27.68 1.73 ;
 RECT 26.435 0.71 27.995 0.85 ;
 RECT 27.54 0.51 27.68 0.71 ;
 RECT 27.54 1.385 27.995 1.525 ;
 RECT 23.445 1.225 23.675 1.245 ;
 RECT 23.445 1.195 24.035 1.225 ;
 END
END RDFFNSRASX2

MACRO RDFFNSRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 24.96 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 15.52 1.16 15.885 1.4 ;
 RECT 15.745 0.695 15.885 1.16 ;
 RECT 16.805 1.905 16.945 1.91 ;
 RECT 15.745 1.765 16.945 1.905 ;
 RECT 16.805 0.71 16.945 1.765 ;
 RECT 15.745 1.4 15.885 1.765 ;
 END
 ANTENNADIFFAREA 0.717 ;
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 24.96 0.08 ;
 RECT 14.655 0.28 14.92 0.44 ;
 RECT 8.335 0.615 8.605 0.755 ;
 RECT 2.18 0.08 2.32 1.055 ;
 RECT 21.785 0.08 22.025 0.31 ;
 RECT 5.525 0.08 5.76 0.595 ;
 RECT 20.65 0.08 20.79 0.325 ;
 RECT 0.68 0.08 0.82 0.775 ;
 RECT 19.435 0.08 19.575 0.31 ;
 RECT 11.575 0.08 11.715 1.155 ;
 RECT 2.925 0.08 3.065 0.39 ;
 RECT 16.305 0.08 16.445 0.965 ;
 RECT 12.65 0.08 12.79 0.525 ;
 RECT 14.71 0.08 14.85 0.28 ;
 RECT 8.4 0.08 8.54 0.615 ;
 END
 END VSS

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.005 0.57 18.485 0.78 ;
 RECT 18.005 0.78 18.375 0.865 ;
 RECT 18.005 0.565 18.375 0.57 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.625 2.305 9.08 2.52 ;
 RECT 8.83 2.12 9.08 2.305 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 23.345 1.41 23.685 1.775 ;
 RECT 21.665 1.965 23.53 2.105 ;
 RECT 19.435 2.195 21.805 2.335 ;
 RECT 21.665 1.41 21.805 1.965 ;
 RECT 23.39 1.775 23.53 1.965 ;
 RECT 19.435 1.365 19.575 2.195 ;
 RECT 20.82 1.345 20.96 2.195 ;
 RECT 21.665 2.105 21.805 2.195 ;
 END
 END VDDG

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.23 1.475 2.56 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 24.96 2.96 ;
 RECT 2.855 2.34 3.105 2.8 ;
 RECT 6.11 2.07 6.25 2.8 ;
 RECT 8.21 2.375 8.35 2.8 ;
 RECT 14.705 2.57 14.845 2.8 ;
 RECT 11.8 2.57 11.94 2.8 ;
 RECT 2.18 1.98 2.32 2.8 ;
 RECT 16.22 2.57 16.36 2.8 ;
 RECT 0.725 1.74 0.865 2.8 ;
 RECT 12.645 2.57 12.785 2.8 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.22 1.7 15.365 1.75 ;
 RECT 14.005 1.84 14.36 1.99 ;
 RECT 14.005 1.75 15.365 1.84 ;
 RECT 14.22 0.905 14.36 1.7 ;
 RECT 15.225 0.915 15.365 1.7 ;
 RECT 15.225 1.84 15.365 1.92 ;
 END
 ANTENNADIFFAREA 0.531 ;
 END QN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.675 0.22 2.04 0.615 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 19.22 0.73 19.79 0.77 ;
 RECT 21.92 1.125 22.02 2.175 ;
 RECT 18.26 0.78 19.79 0.83 ;
 RECT 18.26 0.83 19.32 0.87 ;
 RECT 19.69 0.19 19.79 0.73 ;
 RECT 19.22 0.185 19.32 0.73 ;
 RECT 18.255 0.57 18.485 0.77 ;
 RECT 19.22 2.175 22.02 2.275 ;
 RECT 22.395 0.37 22.495 1.01 ;
 RECT 22.395 1.01 22.645 1.22 ;
 RECT 22.395 1.22 22.495 2.245 ;
 RECT 22.395 2.245 22.68 2.455 ;
 RECT 12.055 0.64 12.155 1.26 ;
 RECT 11.85 1.26 12.155 1.47 ;
 RECT 12.055 1.47 12.155 2.21 ;
 RECT 19.56 1.01 19.795 1.22 ;
 RECT 19.695 1.22 19.795 1.995 ;
 RECT 13.865 0.84 13.965 1.3 ;
 RECT 13.175 1.25 13.435 1.3 ;
 RECT 13.175 1.3 13.965 1.4 ;
 RECT 13.175 1.4 13.435 1.46 ;
 RECT 13.335 0.61 13.435 1.25 ;
 RECT 13.335 1.46 13.435 2.56 ;
 RECT 13.85 0.63 14.08 0.84 ;
 RECT 20 0.19 20.1 0.97 ;
 RECT 20 0.97 20.24 1.18 ;
 RECT 20 1.18 20.1 1.975 ;
 RECT 12.9 1.635 13 1.66 ;
 RECT 12.9 1.66 13.155 1.87 ;
 RECT 12.9 1.87 13 2.565 ;
 RECT 6.2 1.61 6.465 1.82 ;
 RECT 6.365 1.82 6.465 2.49 ;
 RECT 5.995 0.66 6.095 1.51 ;
 RECT 5.995 1.51 6.465 1.61 ;
 RECT 2.44 0.57 2.54 1.495 ;
 RECT 2.245 1.495 2.54 1.745 ;
 RECT 2.44 1.745 2.54 2.37 ;
 RECT 1.965 0.52 2.065 2.465 ;
 RECT 1.725 0.27 2.065 0.52 ;
 RECT 8.66 0.655 8.76 1.235 ;
 RECT 8.08 1.335 8.31 1.475 ;
 RECT 8.08 1.235 8.76 1.335 ;
 RECT 4.635 1.475 4.945 1.71 ;
 RECT 4.635 0.65 4.735 1.475 ;
 RECT 4.635 1.71 4.735 2.475 ;
 RECT 18.46 1.175 18.745 1.305 ;
 RECT 18.46 1.305 18.56 2.64 ;
 RECT 23.095 0.19 23.195 2.64 ;
 RECT 22.085 0.09 23.195 0.19 ;
 RECT 22.085 0.19 22.185 0.94 ;
 RECT 18.46 1.075 18.79 1.175 ;
 RECT 18.46 2.64 23.195 2.74 ;
 RECT 9.055 2.69 10.705 2.695 ;
 RECT 10.53 2.54 10.705 2.69 ;
 RECT 9.845 2.695 10.705 2.79 ;
 RECT 9.055 0.655 9.155 2.595 ;
 RECT 9.055 2.595 9.945 2.69 ;
 RECT 10.53 2.33 10.76 2.54 ;
 RECT 20.91 0.355 21.01 0.985 ;
 RECT 20.91 0.255 21.645 0.355 ;
 RECT 21.415 0.355 21.645 0.465 ;
 RECT 21.08 1.215 21.18 1.815 ;
 RECT 20.52 1.115 21.18 1.215 ;
 RECT 20.52 0.985 21.01 1.115 ;
 RECT 14.485 0.39 14.585 1.4 ;
 RECT 13.48 0.225 13.71 0.29 ;
 RECT 13.48 0.39 13.71 0.435 ;
 RECT 13.48 0.29 14.585 0.39 ;
 RECT 14.485 1.5 14.585 2.35 ;
 RECT 14.975 0.505 15.075 1.4 ;
 RECT 14.975 1.5 15.075 2.35 ;
 RECT 14.485 1.4 15.075 1.5 ;
 RECT 4.145 0.705 4.245 1.17 ;
 RECT 4.145 0.47 4.43 0.705 ;
 RECT 3.56 1.27 3.805 1.46 ;
 RECT 3.56 1.17 4.245 1.27 ;
 RECT 5.895 1.79 5.995 2.465 ;
 RECT 5.68 2.465 5.995 2.71 ;
 RECT 11.29 0.19 11.39 1.795 ;
 RECT 11.29 0.09 13.005 0.19 ;
 RECT 6.385 0.47 6.57 0.5 ;
 RECT 10.595 1.71 10.695 1.795 ;
 RECT 12.905 0.19 13.005 1.18 ;
 RECT 10.595 1.795 11.39 1.895 ;
 RECT 9.575 0.47 9.675 1.61 ;
 RECT 10.125 1.71 10.225 2.445 ;
 RECT 6.34 0.5 6.57 0.71 ;
 RECT 6.385 0.37 9.675 0.47 ;
 RECT 9.575 1.61 10.695 1.71 ;
 RECT 15.99 1.285 16.685 1.385 ;
 RECT 16.585 0.38 16.685 1.285 ;
 RECT 15.99 1.385 16.2 1.435 ;
 RECT 15.99 1.2 16.2 1.285 ;
 RECT 16.005 0.47 16.105 1.2 ;
 RECT 16.005 1.435 16.105 2.645 ;
 RECT 16.585 1.385 16.685 2.645 ;
 RECT 17.255 0.22 17.485 0.28 ;
 RECT 17.255 0.38 17.485 0.435 ;
 RECT 16.585 0.28 17.485 0.38 ;
 RECT 3.215 1.62 3.315 2.375 ;
 RECT 3.28 0.185 10.19 0.19 ;
 RECT 3.28 0.19 5.435 0.285 ;
 RECT 3.28 0.285 3.38 1.52 ;
 RECT 10.09 1.29 11.11 1.39 ;
 RECT 10.09 0.19 10.19 1.29 ;
 RECT 4.1 1.565 4.2 2.375 ;
 RECT 2.78 1.44 3.025 1.52 ;
 RECT 2.78 1.62 3.025 1.69 ;
 RECT 2.78 1.52 3.38 1.62 ;
 RECT 5.335 0.285 5.435 1.24 ;
 RECT 5.335 0.09 10.19 0.185 ;
 RECT 10.88 1.285 11.11 1.29 ;
 RECT 10.88 1.39 11.11 1.615 ;
 RECT 3.215 2.375 4.2 2.475 ;
 RECT 7.765 0.655 7.865 1.13 ;
 RECT 7.765 1.23 7.865 1.655 ;
 RECT 6.85 0.66 6.95 1.13 ;
 RECT 7.765 1.655 8.725 1.755 ;
 RECT 8.625 1.755 8.725 2.31 ;
 RECT 7.765 1.755 7.865 2.57 ;
 RECT 6.85 1.13 7.865 1.23 ;
 RECT 8.625 2.31 8.855 2.52 ;
 RECT 6.84 1.575 6.94 2.485 ;
 RECT 7.35 1.41 7.58 1.475 ;
 RECT 7.35 1.575 7.58 1.62 ;
 RECT 6.84 1.475 7.58 1.575 ;
 RECT 19.22 0.87 19.32 2.175 ;
 RECT 18.255 0.77 19.79 0.78 ;
 LAYER CO ;
 RECT 2.93 0.21 3.06 0.34 ;
 RECT 21.465 0.295 21.595 0.425 ;
 RECT 6.39 0.54 6.52 0.67 ;
 RECT 22.465 1.05 22.595 1.18 ;
 RECT 13.9 0.67 14.03 0.8 ;
 RECT 7.4 1.45 7.53 1.58 ;
 RECT 18.305 0.61 18.435 0.74 ;
 RECT 18.565 1.135 18.695 1.265 ;
 RECT 22.5 2.285 22.63 2.415 ;
 RECT 17.305 0.265 17.435 0.395 ;
 RECT 11.9 1.3 12.03 1.43 ;
 RECT 3.615 1.265 3.745 1.395 ;
 RECT 19.61 1.05 19.74 1.18 ;
 RECT 10.93 1.445 11.06 1.575 ;
 RECT 20.57 1.025 20.7 1.155 ;
 RECT 13.225 1.29 13.355 1.42 ;
 RECT 10.58 2.37 10.71 2.5 ;
 RECT 13.53 0.265 13.66 0.395 ;
 RECT 20.06 1.01 20.19 1.14 ;
 RECT 12.975 1.7 13.105 1.83 ;
 RECT 1.715 2.115 1.845 2.245 ;
 RECT 10.345 0.595 10.475 0.725 ;
 RECT 7.515 0.88 7.645 1.01 ;
 RECT 8.13 1.28 8.26 1.41 ;
 RECT 12.655 0.33 12.785 0.46 ;
 RECT 2.79 0.88 2.92 1.01 ;
 RECT 12.275 1.705 12.405 1.835 ;
 RECT 4.25 0.525 4.38 0.655 ;
 RECT 16.225 2.64 16.355 2.77 ;
 RECT 1.715 0.79 1.845 0.92 ;
 RECT 8.405 0.62 8.535 0.75 ;
 RECT 16.31 0.77 16.44 0.9 ;
 RECT 13.555 1.78 13.685 1.91 ;
 RECT 5.575 0.455 5.705 0.585 ;
 RECT 14.225 0.975 14.355 1.105 ;
 RECT 9.315 0.875 9.445 1.005 ;
 RECT 3.85 2.105 3.98 2.235 ;
 RECT 3.435 1.825 3.565 1.955 ;
 RECT 2.185 0.79 2.315 0.92 ;
 RECT 2.925 2.345 3.055 2.475 ;
 RECT 13.555 0.83 13.685 0.96 ;
 RECT 15.75 0.77 15.88 0.9 ;
 RECT 14.225 1.72 14.355 1.85 ;
 RECT 15.75 1.725 15.88 1.855 ;
 RECT 2.84 1.495 2.97 1.625 ;
 RECT 3.895 0.88 4.025 1.01 ;
 RECT 16.03 1.25 16.16 1.38 ;
 RECT 11.805 2.64 11.935 2.77 ;
 RECT 0.685 0.33 0.815 0.46 ;
 RECT 0.73 2.345 0.86 2.475 ;
 RECT 22.615 0.59 22.745 0.72 ;
 RECT 6.585 2.015 6.715 2.145 ;
 RECT 20.655 0.11 20.785 0.24 ;
 RECT 4.365 0.88 4.495 1.01 ;
 RECT 4.345 2.07 4.475 2.2 ;
 RECT 12.65 2.64 12.78 2.77 ;
 RECT 14.71 2.64 14.84 2.77 ;
 RECT 9.315 1.945 9.445 2.075 ;
 RECT 7.515 1.885 7.645 2.015 ;
 RECT 18.72 0.505 18.85 0.635 ;
 RECT 0.73 1.825 0.86 1.955 ;
 RECT 19.44 1.45 19.57 1.58 ;
 RECT 5.645 2.125 5.775 2.255 ;
 RECT 15.23 1.72 15.36 1.85 ;
 RECT 9.84 0.595 9.97 0.725 ;
 RECT 7.07 2.07 7.2 2.2 ;
 RECT 1.785 0.325 1.915 0.455 ;
 RECT 6.255 1.63 6.385 1.76 ;
 RECT 21.135 0.59 21.265 0.72 ;
 RECT 21.67 1.465 21.8 1.595 ;
 RECT 2.305 1.55 2.435 1.68 ;
 RECT 0.73 2.085 0.86 2.215 ;
 RECT 6.115 2.135 6.245 2.265 ;
 RECT 6.585 0.93 6.715 1.06 ;
 RECT 2.185 2.05 2.315 2.18 ;
 RECT 10.345 1.87 10.475 2 ;
 RECT 16.81 0.78 16.94 0.91 ;
 RECT 21.3 1.38 21.43 1.51 ;
 RECT 7.07 0.88 7.2 1.01 ;
 RECT 21.835 0.115 21.965 0.245 ;
 RECT 23.395 1.45 23.525 1.58 ;
 RECT 20.22 0.41 20.35 0.54 ;
 RECT 3.5 0.905 3.63 1.035 ;
 RECT 15.23 0.975 15.36 1.105 ;
 RECT 9.84 1.9 9.97 2.03 ;
 RECT 4.765 1.525 4.895 1.655 ;
 RECT 20.825 1.42 20.955 1.55 ;
 RECT 4.855 2.125 4.985 2.255 ;
 RECT 16.81 1.71 16.94 1.84 ;
 RECT 18.97 1.4 19.1 1.53 ;
 RECT 14.715 0.305 14.845 0.435 ;
 RECT 20.22 1.46 20.35 1.59 ;
 RECT 8.215 2.445 8.345 2.575 ;
 RECT 11.58 0.955 11.71 1.085 ;
 RECT 0.685 0.59 0.815 0.72 ;
 RECT 19.44 0.11 19.57 0.24 ;
 RECT 5.72 2.515 5.85 2.645 ;
 RECT 22.615 1.44 22.745 1.57 ;
 RECT 12.275 0.96 12.405 1.09 ;
 RECT 2.66 1.995 2.79 2.125 ;
 RECT 8.675 2.35 8.805 2.48 ;
 LAYER M1 ;
 RECT 4.745 2.12 5.845 2.26 ;
 RECT 13.85 0.72 14.08 0.84 ;
 RECT 15.12 0.37 15.26 0.58 ;
 RECT 13.85 0.63 15.26 0.72 ;
 RECT 13.86 0.58 15.26 0.63 ;
 RECT 16.025 0.37 16.165 1.46 ;
 RECT 15.12 0.23 16.165 0.37 ;
 RECT 7.51 1.62 7.65 1.735 ;
 RECT 7.51 1.875 7.65 2.085 ;
 RECT 7.51 1.735 8.265 1.875 ;
 RECT 8.125 1.21 8.265 1.735 ;
 RECT 7.51 0.81 7.65 1.41 ;
 RECT 7.35 1.41 7.65 1.62 ;
 RECT 3.495 1.96 3.635 2.51 ;
 RECT 3.495 1.435 3.635 1.82 ;
 RECT 3.495 0.5 3.635 1.225 ;
 RECT 3.495 1.225 3.795 1.435 ;
 RECT 3.365 1.82 3.635 1.96 ;
 RECT 3.495 2.51 5.97 2.65 ;
 RECT 20.52 1.195 20.66 1.32 ;
 RECT 20.215 1.46 20.355 1.735 ;
 RECT 20.535 0.705 20.675 0.985 ;
 RECT 20.215 0.33 20.355 0.565 ;
 RECT 20.215 1.32 20.66 1.46 ;
 RECT 20.215 0.565 20.675 0.705 ;
 RECT 20.52 0.985 20.75 1.195 ;
 RECT 12.27 1.37 13.405 1.46 ;
 RECT 12.27 1.095 12.41 1.37 ;
 RECT 12.27 1.46 13.4 1.51 ;
 RECT 12.27 1.51 12.41 1.7 ;
 RECT 13.175 1.25 13.405 1.37 ;
 RECT 12.2 0.955 12.47 1.095 ;
 RECT 12.205 1.7 12.48 1.84 ;
 RECT 10.53 2.42 10.76 2.54 ;
 RECT 17.995 2.42 18.135 2.505 ;
 RECT 10.53 2.28 18.135 2.42 ;
 RECT 22.45 2.455 22.59 2.505 ;
 RECT 22.45 2.245 22.68 2.455 ;
 RECT 17.995 2.505 22.59 2.645 ;
 RECT 11.855 0.805 11.995 1.26 ;
 RECT 11.85 1.26 12.08 1.295 ;
 RECT 11.85 1.435 12.08 1.47 ;
 RECT 11.26 1.295 12.08 1.435 ;
 RECT 11.26 1.105 11.4 1.295 ;
 RECT 10.34 0.525 10.48 0.965 ;
 RECT 10.34 1.105 10.48 2.065 ;
 RECT 10.34 0.965 11.4 1.105 ;
 RECT 13.55 0.435 13.69 0.665 ;
 RECT 13.55 0.805 13.69 1.98 ;
 RECT 11.855 0.665 13.69 0.805 ;
 RECT 13.55 0.22 13.69 0.225 ;
 RECT 13.48 0.225 13.71 0.435 ;
 RECT 17.255 0.36 17.485 0.435 ;
 RECT 19.07 0.36 19.21 0.54 ;
 RECT 17.255 0.225 19.21 0.36 ;
 RECT 17.29 0.22 19.21 0.225 ;
 RECT 19.935 0.535 20.075 0.54 ;
 RECT 19.935 0.68 20.075 0.97 ;
 RECT 19.07 0.54 20.075 0.68 ;
 RECT 19.935 0.97 20.24 1.18 ;
 RECT 21.505 0.465 21.645 0.685 ;
 RECT 21.415 0.255 21.645 0.465 ;
 RECT 21.505 0.685 23.065 0.825 ;
 RECT 22.925 0.825 23.065 1.36 ;
 RECT 22.61 1.5 22.75 1.705 ;
 RECT 22.61 0.485 22.75 0.685 ;
 RECT 22.61 1.36 23.065 1.5 ;
 RECT 7.915 2.165 8.055 2.225 ;
 RECT 7.065 0.82 7.205 2.225 ;
 RECT 7.065 2.225 8.055 2.365 ;
 RECT 8.405 1.605 8.545 2.025 ;
 RECT 7.915 2.025 8.545 2.165 ;
 RECT 9.31 1.605 9.45 2.025 ;
 RECT 9.835 0.525 9.975 2.025 ;
 RECT 9.31 0.765 9.45 1.465 ;
 RECT 9.31 2.025 9.975 2.165 ;
 RECT 8.405 1.465 9.45 1.605 ;
 RECT 21.13 0.48 21.27 1.08 ;
 RECT 21.295 1.22 21.435 1.58 ;
 RECT 22.415 1.01 22.645 1.08 ;
 RECT 21.13 1.08 22.645 1.22 ;
 RECT 2.7 1.63 2.84 1.99 ;
 RECT 2.7 1.475 3.045 1.63 ;
 RECT 2.785 0.81 2.925 1.475 ;
 RECT 2.59 1.99 2.84 2.13 ;
 RECT 4.18 0.52 4.78 0.66 ;
 RECT 4.64 0.66 4.78 1.015 ;
 RECT 6.185 0.505 6.57 0.71 ;
 RECT 4.64 1.015 6.325 1.155 ;
 RECT 6.34 0.5 6.57 0.505 ;
 RECT 6.185 0.71 6.325 1.015 ;
 RECT 18.79 0.64 18.93 0.99 ;
 RECT 18.515 1.17 19.105 1.2 ;
 RECT 18.965 1.2 19.105 1.725 ;
 RECT 18.655 0.99 18.965 1.03 ;
 RECT 18.515 1.2 18.745 1.305 ;
 RECT 18.67 0.5 18.93 0.64 ;
 RECT 19.56 1.01 19.79 1.03 ;
 RECT 18.51 1.03 19.79 1.17 ;
 RECT 19.56 1.17 19.79 1.22 ;
 RECT 1.49 1.335 1.63 2.11 ;
 RECT 1.49 0.925 1.63 1.195 ;
 RECT 1.49 2.11 1.915 2.25 ;
 RECT 1.49 0.785 1.915 0.925 ;
 RECT 1.49 1.195 2.6 1.335 ;
 RECT 2.46 0.67 2.6 1.195 ;
 RECT 3.205 0.22 4.03 0.36 ;
 RECT 3.89 0.36 4.03 0.9 ;
 RECT 3.965 1.08 4.105 1.945 ;
 RECT 2.46 0.53 3.345 0.67 ;
 RECT 3.205 0.36 3.345 0.53 ;
 RECT 3.89 0.9 4.105 1.08 ;
 RECT 3.845 1.945 4.105 2.17 ;
 RECT 3.845 2.17 3.985 2.305 ;
 RECT 5.625 1.79 5.765 1.82 ;
 RECT 4.36 0.805 4.5 1.82 ;
 RECT 4.27 1.96 4.55 2.215 ;
 RECT 4.27 1.82 5.765 1.96 ;
 RECT 6.2 1.58 6.44 1.65 ;
 RECT 5.625 1.65 6.44 1.79 ;
 RECT 6.2 1.79 6.44 1.835 ;
 RECT 10.875 1.43 11.11 1.615 ;
 RECT 10.875 1.615 11.015 1.985 ;
 RECT 10.88 1.405 11.11 1.43 ;
 RECT 10.875 1.985 13.11 2.125 ;
 RECT 12.925 1.87 13.11 1.985 ;
 RECT 12.925 1.66 13.155 1.87 ;
 RECT 4.695 1.52 5.445 1.66 ;
 RECT 5.305 1.44 5.445 1.52 ;
 RECT 6.58 0.865 6.72 1.3 ;
 RECT 6.58 1.44 6.72 2.215 ;
 RECT 5.305 1.3 6.72 1.44 ;
 END
END RDFFNSRX1

MACRO RDFFNSRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 24.64 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.585 0.57 18.065 0.78 ;
 RECT 17.585 0.565 17.955 0.57 ;
 RECT 17.585 0.78 17.955 0.865 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 24.64 0.08 ;
 RECT 13.645 0.28 13.91 0.44 ;
 RECT 1.505 0.08 1.645 1.055 ;
 RECT 4.85 0.08 5.085 0.595 ;
 RECT 21.365 0.08 21.605 0.31 ;
 RECT 10.34 0.08 10.48 1.155 ;
 RECT 16.575 0.08 16.715 0.965 ;
 RECT 11.415 0.08 11.555 0.525 ;
 RECT 15.63 0.08 15.77 0.965 ;
 RECT 19.015 0.08 19.155 0.31 ;
 RECT 2.25 0.08 2.39 0.39 ;
 RECT 0.47 0.08 0.61 0.775 ;
 RECT 7.725 0.08 7.865 0.815 ;
 RECT 20.23 0.08 20.37 0.325 ;
 RECT 13.7 0.08 13.84 0.28 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.01 1.205 13.365 1.445 ;
 RECT 12.615 1.705 14.77 1.845 ;
 RECT 13.22 0.88 13.36 1.205 ;
 RECT 14.23 0.89 14.37 1.705 ;
 RECT 13.22 1.445 13.36 1.705 ;
 END
 ANTENNADIFFAREA 0.815 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.845 1.16 15.2 1.4 ;
 RECT 14.97 0.695 15.11 1.16 ;
 RECT 14.97 1.765 17.185 1.905 ;
 RECT 14.97 1.4 15.11 1.765 ;
 RECT 17.045 0.71 17.185 1.765 ;
 RECT 16.1 0.71 16.24 1.765 ;
 END
 ANTENNADIFFAREA 1.132 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 24.64 2.96 ;
 RECT 2.18 2.34 2.43 2.8 ;
 RECT 7.535 2.375 7.675 2.8 ;
 RECT 14.095 2.57 14.235 2.8 ;
 RECT 15.445 2.57 15.585 2.8 ;
 RECT 13.145 2.57 13.285 2.8 ;
 RECT 5.435 2.07 5.575 2.8 ;
 RECT 11.41 2.57 11.55 2.8 ;
 RECT 10.565 2.57 10.705 2.8 ;
 RECT 16.43 2.57 16.57 2.8 ;
 RECT 0.505 1.74 0.645 2.8 ;
 RECT 1.505 1.98 1.645 2.8 ;
 END
 END VDD

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.115 1.235 7.4 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 22.925 1.41 23.265 1.775 ;
 RECT 21.245 1.965 23.11 2.105 ;
 RECT 19.015 2.195 21.385 2.335 ;
 RECT 22.97 1.775 23.11 1.965 ;
 RECT 21.245 1.41 21.385 1.965 ;
 RECT 19.015 1.365 19.155 2.195 ;
 RECT 20.4 1.345 20.54 2.195 ;
 RECT 21.245 2.105 21.385 2.195 ;
 END
 END VDDG

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 1.475 1.885 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 0.22 1.365 0.615 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 19.58 1.18 19.68 1.975 ;
 RECT 1.57 1.495 1.865 1.745 ;
 RECT 1.765 1.745 1.865 2.37 ;
 RECT 5.525 1.61 5.79 1.82 ;
 RECT 5.69 1.82 5.79 2.49 ;
 RECT 5.32 0.66 5.42 1.51 ;
 RECT 5.32 1.51 5.79 1.61 ;
 RECT 3.96 1.475 4.27 1.71 ;
 RECT 3.96 0.65 4.06 1.475 ;
 RECT 3.96 1.71 4.06 2.475 ;
 RECT 5.005 2.465 5.32 2.71 ;
 RECT 5.22 1.79 5.32 2.465 ;
 RECT 1.05 0.27 1.39 0.52 ;
 RECT 1.29 0.52 1.39 2.465 ;
 RECT 9.955 0.09 11.77 0.19 ;
 RECT 11.67 0.19 11.77 1.18 ;
 RECT 9.955 0.19 10.185 0.45 ;
 RECT 8.765 0.47 9 0.59 ;
 RECT 8.9 0.59 9 1.61 ;
 RECT 5.71 0.47 5.895 0.5 ;
 RECT 9.45 1.71 9.55 2.445 ;
 RECT 8.9 1.61 9.55 1.71 ;
 RECT 5.71 0.37 9 0.47 ;
 RECT 5.665 0.5 5.895 0.71 ;
 RECT 18.8 0.87 18.9 2.175 ;
 RECT 17.835 0.77 19.37 0.78 ;
 RECT 18.8 0.73 19.37 0.77 ;
 RECT 21.5 1.125 21.6 2.175 ;
 RECT 17.84 0.78 19.37 0.83 ;
 RECT 17.84 0.83 18.9 0.87 ;
 RECT 19.27 0.19 19.37 0.73 ;
 RECT 18.8 0.185 18.9 0.73 ;
 RECT 17.835 0.57 18.065 0.77 ;
 RECT 18.8 2.175 21.6 2.275 ;
 RECT 15.225 1.2 15.525 1.285 ;
 RECT 15.225 0.525 15.325 1.2 ;
 RECT 15.225 1.285 16.935 1.385 ;
 RECT 16.83 0.38 16.93 1.285 ;
 RECT 15.225 1.435 15.325 2.625 ;
 RECT 15.225 1.385 15.525 1.435 ;
 RECT 16.21 1.385 16.31 2.625 ;
 RECT 16.355 0.525 16.455 1.285 ;
 RECT 15.715 1.385 15.815 2.625 ;
 RECT 16.685 1.385 16.785 2.625 ;
 RECT 15.885 0.52 15.985 1.285 ;
 RECT 17.125 0.22 17.355 0.28 ;
 RECT 17.125 0.38 17.355 0.435 ;
 RECT 16.83 0.28 17.355 0.38 ;
 RECT 13.885 1.5 13.985 2.275 ;
 RECT 13.475 0.39 13.575 1.4 ;
 RECT 13.955 0.37 14.055 1.4 ;
 RECT 12.935 1.4 14.45 1.5 ;
 RECT 12.935 1.5 13.035 2.275 ;
 RECT 14.35 1.5 14.45 2.275 ;
 RECT 13.41 1.5 13.51 2.275 ;
 RECT 12.605 0.29 13.575 0.39 ;
 RECT 12.605 0.22 12.835 0.29 ;
 RECT 12.605 0.39 12.835 0.43 ;
 RECT 20.49 0.355 20.59 0.985 ;
 RECT 20.66 1.215 20.76 1.815 ;
 RECT 20.1 1.115 20.76 1.215 ;
 RECT 20.1 0.985 20.59 1.115 ;
 RECT 20.995 0.355 21.225 0.465 ;
 RECT 20.49 0.255 21.225 0.355 ;
 RECT 19.14 1.01 19.375 1.22 ;
 RECT 19.275 1.22 19.375 1.995 ;
 RECT 21.975 0.37 22.075 1.01 ;
 RECT 21.975 1.01 22.225 1.22 ;
 RECT 21.975 1.22 22.075 2.245 ;
 RECT 21.975 2.245 22.26 2.455 ;
 RECT 18.04 1.075 18.325 1.305 ;
 RECT 22.675 0.19 22.775 2.64 ;
 RECT 21.665 0.09 22.775 0.19 ;
 RECT 18.04 1.305 18.14 2.64 ;
 RECT 21.665 0.19 21.765 0.94 ;
 RECT 18.04 2.64 22.775 2.74 ;
 RECT 8.38 2.69 10.03 2.695 ;
 RECT 9.855 2.54 10.03 2.69 ;
 RECT 9.17 2.695 10.03 2.79 ;
 RECT 8.38 0.655 8.48 2.595 ;
 RECT 8.38 2.595 9.27 2.69 ;
 RECT 9.855 2.33 10.085 2.54 ;
 RECT 10.82 0.64 10.92 1.26 ;
 RECT 10.615 1.26 10.92 1.47 ;
 RECT 10.82 1.47 10.92 2.21 ;
 RECT 2.54 1.62 2.64 2.375 ;
 RECT 2.605 0.185 9.515 0.19 ;
 RECT 2.605 0.19 4.76 0.285 ;
 RECT 2.605 0.285 2.705 1.52 ;
 RECT 9.415 1.29 10.32 1.39 ;
 RECT 9.415 0.19 9.515 1.29 ;
 RECT 3.425 1.565 3.525 2.375 ;
 RECT 2.105 1.44 2.35 1.52 ;
 RECT 2.105 1.62 2.35 1.69 ;
 RECT 2.105 1.52 2.705 1.62 ;
 RECT 4.66 0.285 4.76 1.24 ;
 RECT 4.66 0.09 9.515 0.185 ;
 RECT 10.09 1.39 10.32 1.82 ;
 RECT 2.54 2.375 3.525 2.475 ;
 RECT 3.47 0.705 3.57 1.17 ;
 RECT 3.47 0.47 3.755 0.705 ;
 RECT 2.885 1.17 3.57 1.27 ;
 RECT 2.885 1.27 3.13 1.46 ;
 RECT 11.665 1.635 11.765 1.66 ;
 RECT 11.665 1.66 11.92 1.87 ;
 RECT 11.665 1.87 11.765 2.565 ;
 RECT 6.165 1.575 6.265 2.485 ;
 RECT 6.675 1.41 6.905 1.475 ;
 RECT 6.675 1.575 6.905 1.62 ;
 RECT 6.165 1.475 6.905 1.575 ;
 RECT 7.09 1.45 7.19 1.655 ;
 RECT 7.09 1.755 7.19 2.57 ;
 RECT 7.09 1.655 8.05 1.755 ;
 RECT 7.95 1.755 8.05 2.355 ;
 RECT 7.09 0.655 7.19 1.13 ;
 RECT 7.09 1.23 7.19 1.24 ;
 RECT 6.175 0.66 6.275 1.13 ;
 RECT 7.09 1.24 7.345 1.45 ;
 RECT 6.175 1.13 7.19 1.23 ;
 RECT 12.1 1.195 12.2 1.25 ;
 RECT 11.945 1.25 12.2 1.46 ;
 RECT 12.1 1.46 12.2 2.56 ;
 RECT 12.63 0.84 12.73 1.095 ;
 RECT 12.1 0.61 12.2 1.095 ;
 RECT 12.1 1.095 12.73 1.195 ;
 RECT 12.615 0.63 12.845 0.84 ;
 RECT 19.58 0.19 19.68 0.97 ;
 RECT 19.58 0.97 19.82 1.18 ;
 RECT 7.985 0.655 8.085 1.24 ;
 RECT 7.855 1.24 8.085 1.475 ;
 RECT 1.765 0.57 1.865 1.495 ;
 LAYER CO ;
 RECT 22.195 0.59 22.325 0.72 ;
 RECT 13.705 0.305 13.835 0.435 ;
 RECT 8.64 1.945 8.77 2.075 ;
 RECT 14.975 1.725 15.105 1.855 ;
 RECT 9.67 1.87 9.8 2 ;
 RECT 14.975 0.77 15.105 0.9 ;
 RECT 2.825 0.905 2.955 1.035 ;
 RECT 17.05 0.78 17.18 0.91 ;
 RECT 8.64 0.875 8.77 1.005 ;
 RECT 15.45 2.64 15.58 2.77 ;
 RECT 9.165 1.9 9.295 2.03 ;
 RECT 16.58 0.78 16.71 0.91 ;
 RECT 22.195 1.44 22.325 1.57 ;
 RECT 3.575 0.525 3.705 0.655 ;
 RECT 15.95 1.77 16.08 1.9 ;
 RECT 9.165 0.595 9.295 0.725 ;
 RECT 11.04 0.96 11.17 1.09 ;
 RECT 13.15 2.64 13.28 2.77 ;
 RECT 20.235 0.11 20.365 0.24 ;
 RECT 15.355 1.25 15.485 1.38 ;
 RECT 19.02 0.11 19.15 0.24 ;
 RECT 0.475 0.33 0.605 0.46 ;
 RECT 3.175 2.105 3.305 2.235 ;
 RECT 7.73 0.62 7.86 0.75 ;
 RECT 21.25 1.465 21.38 1.595 ;
 RECT 16.105 0.79 16.235 0.92 ;
 RECT 5.91 2.015 6.04 2.145 ;
 RECT 5.91 0.93 6.04 1.06 ;
 RECT 16.435 2.64 16.565 2.77 ;
 RECT 4.09 1.525 4.22 1.655 ;
 RECT 1.04 2.115 1.17 2.245 ;
 RECT 6.84 1.885 6.97 2.015 ;
 RECT 6.395 0.88 6.525 1.01 ;
 RECT 11.04 1.705 11.17 1.835 ;
 RECT 1.985 1.995 2.115 2.125 ;
 RECT 16.91 1.77 17.04 1.9 ;
 RECT 20.715 0.59 20.845 0.72 ;
 RECT 11.415 2.64 11.545 2.77 ;
 RECT 15.635 0.77 15.765 0.9 ;
 RECT 3.22 0.88 3.35 1.01 ;
 RECT 22.975 1.45 23.105 1.58 ;
 RECT 2.25 2.345 2.38 2.475 ;
 RECT 1.11 0.325 1.24 0.455 ;
 RECT 2.255 0.21 2.385 0.34 ;
 RECT 19.8 1.46 19.93 1.59 ;
 RECT 5.44 2.135 5.57 2.265 ;
 RECT 19.8 0.41 19.93 0.54 ;
 RECT 10.57 2.64 10.7 2.77 ;
 RECT 11.42 0.33 11.55 0.46 ;
 RECT 10.345 0.955 10.475 1.085 ;
 RECT 14.235 0.96 14.365 1.09 ;
 RECT 7.54 2.445 7.67 2.575 ;
 RECT 4.18 2.125 4.31 2.255 ;
 RECT 5.045 2.515 5.175 2.645 ;
 RECT 1.04 0.79 1.17 0.92 ;
 RECT 12.32 0.83 12.45 0.96 ;
 RECT 20.88 1.38 21.01 1.51 ;
 RECT 13.635 1.71 13.765 1.84 ;
 RECT 2.165 1.495 2.295 1.625 ;
 RECT 13.225 0.95 13.355 1.08 ;
 RECT 4.9 0.455 5.03 0.585 ;
 RECT 18.3 0.505 18.43 0.635 ;
 RECT 1.51 2.05 1.64 2.18 ;
 RECT 20.405 1.42 20.535 1.55 ;
 RECT 6.84 0.88 6.97 1.01 ;
 RECT 3.67 2.07 3.8 2.2 ;
 RECT 0.51 2.085 0.64 2.215 ;
 RECT 9.67 0.595 9.8 0.725 ;
 RECT 12.685 1.71 12.815 1.84 ;
 RECT 14.57 1.71 14.7 1.84 ;
 RECT 12.32 1.78 12.45 1.91 ;
 RECT 0.51 2.345 0.64 2.475 ;
 RECT 7.905 1.28 8.035 1.41 ;
 RECT 18.55 1.4 18.68 1.53 ;
 RECT 5.58 1.63 5.71 1.76 ;
 RECT 19.02 1.45 19.15 1.58 ;
 RECT 21.415 0.115 21.545 0.245 ;
 RECT 2.115 0.88 2.245 1.01 ;
 RECT 4.97 2.125 5.1 2.255 ;
 RECT 14.1 2.64 14.23 2.77 ;
 RECT 6.395 2.07 6.525 2.2 ;
 RECT 0.475 0.59 0.605 0.72 ;
 RECT 1.63 1.55 1.76 1.68 ;
 RECT 0.51 1.825 0.64 1.955 ;
 RECT 2.76 1.825 2.89 1.955 ;
 RECT 1.51 0.79 1.64 0.92 ;
 RECT 3.69 0.88 3.82 1.01 ;
 RECT 8.815 0.42 8.945 0.55 ;
 RECT 10.005 0.28 10.135 0.41 ;
 RECT 5.715 0.54 5.845 0.67 ;
 RECT 17.885 0.61 18.015 0.74 ;
 RECT 17.175 0.265 17.305 0.395 ;
 RECT 12.655 0.26 12.785 0.39 ;
 RECT 20.15 1.025 20.28 1.155 ;
 RECT 22.045 1.05 22.175 1.18 ;
 RECT 21.045 0.295 21.175 0.425 ;
 RECT 19.19 1.05 19.32 1.18 ;
 RECT 22.08 2.285 22.21 2.415 ;
 RECT 18.145 1.135 18.275 1.265 ;
 RECT 9.905 2.37 10.035 2.5 ;
 RECT 10.665 1.3 10.795 1.43 ;
 RECT 10.14 1.65 10.27 1.78 ;
 RECT 11.995 1.29 12.125 1.42 ;
 RECT 2.94 1.265 3.07 1.395 ;
 RECT 11.74 1.7 11.87 1.83 ;
 RECT 6.725 1.45 6.855 1.58 ;
 RECT 7.165 1.28 7.295 1.41 ;
 RECT 12.665 0.67 12.795 0.8 ;
 RECT 19.64 1.01 19.77 1.14 ;
 LAYER M1 ;
 RECT 4.07 2.12 5.17 2.26 ;
 RECT 4.02 1.52 4.77 1.66 ;
 RECT 4.63 1.44 4.77 1.52 ;
 RECT 5.905 0.865 6.045 1.3 ;
 RECT 5.905 1.44 6.045 2.215 ;
 RECT 4.63 1.3 6.045 1.44 ;
 RECT 6.39 0.82 6.53 2.225 ;
 RECT 7.24 2.165 7.38 2.225 ;
 RECT 6.39 2.225 7.38 2.365 ;
 RECT 8.635 0.765 8.775 2.025 ;
 RECT 9.16 0.525 9.3 2.025 ;
 RECT 7.24 2.025 9.3 2.165 ;
 RECT 2.025 1.63 2.165 1.99 ;
 RECT 2.025 1.475 2.37 1.63 ;
 RECT 2.11 0.81 2.25 1.475 ;
 RECT 1.915 1.99 2.165 2.13 ;
 RECT 4.95 1.79 5.09 1.82 ;
 RECT 3.685 0.805 3.825 1.82 ;
 RECT 3.595 1.96 3.875 2.215 ;
 RECT 3.595 1.82 5.09 1.96 ;
 RECT 5.525 1.58 5.765 1.65 ;
 RECT 4.95 1.65 5.765 1.79 ;
 RECT 5.525 1.79 5.765 1.835 ;
 RECT 0.815 0.925 0.955 1.195 ;
 RECT 0.815 1.335 0.955 2.11 ;
 RECT 0.815 1.195 1.925 1.335 ;
 RECT 1.785 0.67 1.925 1.195 ;
 RECT 0.815 0.785 1.24 0.925 ;
 RECT 0.815 2.11 1.24 2.25 ;
 RECT 3.215 0.36 3.355 0.9 ;
 RECT 3.29 1.08 3.43 1.945 ;
 RECT 2.53 0.22 3.355 0.36 ;
 RECT 3.17 2.17 3.31 2.305 ;
 RECT 3.17 1.945 3.43 2.17 ;
 RECT 3.215 0.9 3.43 1.08 ;
 RECT 2.53 0.36 2.67 0.53 ;
 RECT 1.785 0.53 2.67 0.67 ;
 RECT 9.955 0.38 10.185 0.45 ;
 RECT 8.765 0.38 8.995 0.59 ;
 RECT 8.765 0.24 10.2 0.38 ;
 RECT 3.505 0.52 4.105 0.66 ;
 RECT 3.965 0.66 4.105 1.015 ;
 RECT 5.51 0.505 5.895 0.71 ;
 RECT 5.665 0.5 5.895 0.505 ;
 RECT 3.965 1.015 5.65 1.155 ;
 RECT 5.51 0.71 5.65 1.015 ;
 RECT 20.115 0.705 20.255 0.985 ;
 RECT 19.795 0.33 19.935 0.565 ;
 RECT 20.1 1.195 20.24 1.32 ;
 RECT 19.795 1.46 19.935 1.735 ;
 RECT 19.795 0.565 20.255 0.705 ;
 RECT 19.795 1.32 20.24 1.46 ;
 RECT 20.1 0.985 20.33 1.195 ;
 RECT 20.71 0.48 20.85 1.08 ;
 RECT 20.875 1.22 21.015 1.58 ;
 RECT 21.995 1.01 22.225 1.08 ;
 RECT 20.71 1.08 22.225 1.22 ;
 RECT 21.085 0.465 21.225 0.685 ;
 RECT 20.995 0.255 21.225 0.465 ;
 RECT 22.505 0.825 22.645 1.36 ;
 RECT 21.085 0.685 22.645 0.825 ;
 RECT 22.19 1.5 22.33 1.705 ;
 RECT 22.19 0.485 22.33 0.685 ;
 RECT 22.19 1.36 22.645 1.5 ;
 RECT 18.37 0.64 18.51 0.99 ;
 RECT 18.095 1.17 18.685 1.2 ;
 RECT 18.545 1.2 18.685 1.725 ;
 RECT 18.095 0.99 18.545 1.03 ;
 RECT 18.095 1.2 18.325 1.305 ;
 RECT 18.25 0.5 18.51 0.64 ;
 RECT 19.14 1.01 19.37 1.03 ;
 RECT 18.095 1.03 19.37 1.17 ;
 RECT 19.14 1.17 19.37 1.22 ;
 RECT 9.855 2.42 10.085 2.54 ;
 RECT 17.575 2.42 17.715 2.505 ;
 RECT 9.855 2.28 17.715 2.42 ;
 RECT 22.03 2.455 22.17 2.505 ;
 RECT 22.03 2.245 22.26 2.455 ;
 RECT 17.575 2.505 22.17 2.645 ;
 RECT 10.62 0.805 10.76 1.26 ;
 RECT 10.615 1.26 10.845 1.3 ;
 RECT 10.615 1.44 10.845 1.47 ;
 RECT 9.665 1.3 10.845 1.44 ;
 RECT 9.665 0.525 9.805 1.3 ;
 RECT 9.665 1.44 9.805 2.065 ;
 RECT 12.315 0.43 12.455 0.665 ;
 RECT 10.62 0.665 12.455 0.805 ;
 RECT 12.315 0.805 12.455 1.98 ;
 RECT 12.315 0.22 12.835 0.43 ;
 RECT 11.035 1.095 11.175 1.255 ;
 RECT 11.035 1.255 12.175 1.395 ;
 RECT 11.035 1.395 11.175 1.7 ;
 RECT 11.945 1.25 12.175 1.255 ;
 RECT 11.945 1.395 12.175 1.46 ;
 RECT 10.97 1.7 11.245 1.84 ;
 RECT 10.965 0.955 11.235 1.095 ;
 RECT 2.82 1.96 2.96 2.51 ;
 RECT 2.82 1.435 2.96 1.82 ;
 RECT 2.82 0.5 2.96 1.225 ;
 RECT 2.82 1.225 3.12 1.435 ;
 RECT 2.69 1.82 2.96 1.96 ;
 RECT 2.82 2.51 5.295 2.65 ;
 RECT 10.12 1.82 10.26 1.985 ;
 RECT 10.12 1.985 11.875 2.125 ;
 RECT 11.69 1.87 11.875 1.985 ;
 RECT 10.09 1.61 10.32 1.82 ;
 RECT 11.69 1.66 11.92 1.87 ;
 RECT 6.835 1.62 6.975 1.735 ;
 RECT 6.835 1.875 6.975 2.085 ;
 RECT 6.835 0.81 6.975 1.41 ;
 RECT 6.675 1.41 6.975 1.62 ;
 RECT 7.585 1.415 7.725 1.735 ;
 RECT 6.835 1.735 7.725 1.875 ;
 RECT 7.585 1.275 8.105 1.415 ;
 RECT 12.615 0.72 12.845 0.84 ;
 RECT 14.11 0.37 14.25 0.58 ;
 RECT 12.615 0.58 14.25 0.72 ;
 RECT 15.35 0.37 15.49 1.46 ;
 RECT 14.11 0.23 15.49 0.37 ;
 RECT 17.125 0.36 17.355 0.435 ;
 RECT 17.115 0.22 18.79 0.36 ;
 RECT 18.65 0.36 18.79 0.54 ;
 RECT 19.515 0.535 19.655 0.54 ;
 RECT 19.515 0.68 19.655 0.97 ;
 RECT 18.65 0.54 19.655 0.68 ;
 RECT 19.515 0.97 19.82 1.18 ;
 END
END RDFFNSRX2

MACRO RDFFSRARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 25.6 BY 2.88 ;
 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.01 0.465 4.25 0.695 ;
 RECT 4.055 0.735 5.13 0.875 ;
 RECT 9.875 1.09 12.245 1.23 ;
 RECT 4.055 0.695 4.25 0.735 ;
 RECT 4.99 0.22 6.625 0.36 ;
 RECT 4.99 0.36 5.13 0.735 ;
 RECT 6.485 0.525 7.03 0.665 ;
 RECT 6.89 0.905 8.005 1.045 ;
 RECT 7.86 0.245 10.01 0.255 ;
 RECT 7.86 0.255 10.015 0.385 ;
 RECT 9.875 0.385 10.015 1.09 ;
 RECT 12.105 0.81 12.245 1.09 ;
 RECT 12.105 0.6 12.395 0.81 ;
 RECT 6.485 0.36 6.625 0.525 ;
 RECT 6.89 0.665 7.03 0.905 ;
 RECT 7.865 0.385 8.005 0.905 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 25.6 0.08 ;
 RECT 22.515 0.08 22.755 0.26 ;
 RECT 7.425 0.615 7.695 0.755 ;
 RECT 15.105 0.335 15.37 0.495 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 2.015 0.08 2.155 0.39 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.615 0.08 4.85 0.595 ;
 RECT 11.35 0.08 11.49 0.945 ;
 RECT 12.855 0.08 12.995 0.525 ;
 RECT 20.165 0.08 20.305 0.36 ;
 RECT 16.875 0.08 17.015 0.82 ;
 RECT 21.38 0.08 21.52 0.35 ;
 RECT 7.49 0.08 7.63 0.615 ;
 RECT 15.16 0.08 15.3 0.335 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 25.6 2.96 ;
 RECT 1.945 2.34 2.195 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.27 1.98 1.41 2.8 ;
 RECT 5.2 2.07 5.34 2.8 ;
 RECT 7.3 2.375 7.44 2.8 ;
 RECT 11.95 2.57 12.09 2.8 ;
 RECT 15.075 2.57 15.215 2.8 ;
 RECT 12.85 2.57 12.99 2.8 ;
 RECT 16.79 2.57 16.93 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.475 1.65 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.765 0.22 1.13 0.615 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.57 1.185 14.81 1.425 ;
 RECT 14.67 0.915 14.81 1.185 ;
 RECT 15.665 1.84 15.805 1.9 ;
 RECT 14.67 1.7 15.805 1.84 ;
 RECT 15.665 0.915 15.805 1.7 ;
 RECT 14.67 1.84 14.81 1.9 ;
 RECT 14.67 1.425 14.81 1.7 ;
 END
 ANTENNADIFFAREA 0.961 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 16.215 1.185 16.455 1.425 ;
 RECT 16.315 0.55 16.455 1.185 ;
 RECT 17.375 1.905 17.515 1.91 ;
 RECT 16.315 1.765 17.515 1.905 ;
 RECT 17.375 0.56 17.515 1.765 ;
 RECT 16.315 1.905 16.455 1.915 ;
 RECT 16.315 1.425 16.455 1.765 ;
 END
 ANTENNADIFFAREA 0.725 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.715 2.33 8.12 2.54 ;
 RECT 7.78 2.54 8.12 2.545 ;
 RECT 7.78 2.12 8.12 2.33 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.845 0.59 19.215 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 24.075 1.435 24.415 1.8 ;
 RECT 22.395 1.99 24.26 2.13 ;
 RECT 20.165 2.22 22.535 2.36 ;
 RECT 22.395 1.435 22.535 1.99 ;
 RECT 24.12 1.8 24.26 1.99 ;
 RECT 20.165 1.39 20.305 2.22 ;
 RECT 21.55 1.37 21.69 2.22 ;
 RECT 22.395 2.13 22.535 2.22 ;
 END
 END VDDG

 OBS
 LAYER PO ;
 RECT 6.855 1.655 7.815 1.755 ;
 RECT 7.715 1.755 7.815 2.33 ;
 RECT 6.855 1.755 6.955 2.57 ;
 RECT 5.94 1.13 6.955 1.23 ;
 RECT 7.715 2.33 7.945 2.54 ;
 RECT 20.425 1.245 20.525 2.02 ;
 RECT 20.295 1.035 20.525 1.245 ;
 RECT 21.64 0.38 21.74 0.96 ;
 RECT 21.64 1.06 21.74 1.14 ;
 RECT 21.22 0.935 21.45 0.96 ;
 RECT 21.22 0.96 21.74 1.06 ;
 RECT 21.22 1.06 21.45 1.145 ;
 RECT 21.64 1.14 21.91 1.24 ;
 RECT 21.81 1.24 21.91 1.84 ;
 RECT 22.005 0.22 22.235 0.28 ;
 RECT 22.005 0.38 22.235 0.43 ;
 RECT 21.64 0.28 22.235 0.38 ;
 RECT 19.19 1.2 19.475 1.245 ;
 RECT 23.825 0.195 23.925 2.665 ;
 RECT 22.815 0.095 23.925 0.195 ;
 RECT 22.815 0.195 22.915 0.945 ;
 RECT 19.19 1.245 19.29 2.665 ;
 RECT 19.245 1.035 19.475 1.1 ;
 RECT 19.19 2.665 23.925 2.765 ;
 RECT 19.19 1.1 19.52 1.2 ;
 RECT 20.73 0.215 20.83 0.995 ;
 RECT 20.73 0.995 20.97 1.205 ;
 RECT 20.73 1.205 20.83 2 ;
 RECT 23.125 2.27 23.41 2.48 ;
 RECT 23.125 1.2 23.225 2.27 ;
 RECT 23.125 0.375 23.225 0.99 ;
 RECT 23.125 0.99 23.375 1.2 ;
 RECT 19.95 0.21 20.05 0.755 ;
 RECT 19.95 0.855 20.05 2.2 ;
 RECT 22.815 1.125 22.915 2.2 ;
 RECT 18.985 0.755 20.52 0.84 ;
 RECT 18.985 0.84 20.515 0.855 ;
 RECT 20.42 0.215 20.52 0.755 ;
 RECT 18.985 0.595 19.215 0.755 ;
 RECT 19.95 2.2 22.915 2.3 ;
 RECT 17.155 0.19 17.255 1.33 ;
 RECT 18.405 0.19 18.505 0.22 ;
 RECT 16.56 1.2 16.77 1.33 ;
 RECT 16.56 1.43 16.77 1.435 ;
 RECT 16.56 1.33 17.255 1.43 ;
 RECT 16.575 0.4 16.675 1.2 ;
 RECT 16.575 1.435 16.675 2.585 ;
 RECT 17.155 1.43 17.255 2.58 ;
 RECT 17.155 0.09 18.505 0.19 ;
 RECT 18.405 0.22 18.635 0.43 ;
 RECT 10.155 0.795 10.32 0.925 ;
 RECT 9.475 0.885 9.705 0.925 ;
 RECT 9.475 1.025 9.705 1.095 ;
 RECT 9.475 0.925 10.32 1.025 ;
 RECT 10.155 0.585 10.385 0.795 ;
 RECT 13.105 1.635 13.205 1.66 ;
 RECT 13.105 1.66 13.36 1.87 ;
 RECT 13.105 1.87 13.205 2.565 ;
 RECT 13.685 0.29 15.035 0.39 ;
 RECT 14.935 0.39 15.035 1.17 ;
 RECT 14.935 1.27 15.035 2.375 ;
 RECT 15.45 0.38 15.55 1.17 ;
 RECT 15.45 1.27 15.55 2.375 ;
 RECT 13.685 0.225 13.915 0.29 ;
 RECT 13.685 0.39 13.915 0.435 ;
 RECT 14.935 1.17 15.55 1.27 ;
 RECT 13.38 1.25 13.64 1.3 ;
 RECT 13.54 0.61 13.64 1.25 ;
 RECT 13.38 1.4 13.64 1.46 ;
 RECT 13.54 1.46 13.64 2.56 ;
 RECT 14.07 0.84 14.17 1.3 ;
 RECT 13.38 1.3 14.17 1.4 ;
 RECT 14.055 0.63 14.285 0.84 ;
 RECT 12.205 0.81 12.305 2.21 ;
 RECT 12.165 0.6 12.395 0.81 ;
 RECT 10.88 0.455 11.9 0.47 ;
 RECT 10.96 0.37 11.9 0.455 ;
 RECT 10.88 0.47 11.11 0.665 ;
 RECT 11.735 0.47 11.9 0.625 ;
 RECT 11.735 0.835 11.835 2.21 ;
 RECT 11.735 0.625 11.965 0.835 ;
 RECT 8.145 2.69 10.055 2.79 ;
 RECT 9.955 2.54 10.055 2.69 ;
 RECT 8.145 0.655 8.245 2.69 ;
 RECT 9.955 2.33 10.185 2.54 ;
 RECT 9.18 0.19 9.28 1.29 ;
 RECT 2.69 0.185 9.28 0.19 ;
 RECT 10.075 1.39 10.27 1.405 ;
 RECT 2.69 0.285 2.79 0.51 ;
 RECT 2.69 0.19 4.525 0.285 ;
 RECT 4.425 0.285 4.525 1.24 ;
 RECT 4.425 0.09 9.28 0.185 ;
 RECT 9.18 1.29 10.27 1.39 ;
 RECT 2.65 0.51 2.895 0.755 ;
 RECT 10.075 1.405 10.305 1.615 ;
 RECT 5.475 0.47 5.66 0.5 ;
 RECT 13.11 0.19 13.21 1.18 ;
 RECT 10.57 0.19 10.67 1.91 ;
 RECT 9.75 1.71 9.85 1.91 ;
 RECT 8.665 1.61 9.85 1.71 ;
 RECT 8.665 0.47 8.765 1.61 ;
 RECT 9.215 1.71 9.315 2.445 ;
 RECT 10.57 0.09 13.21 0.19 ;
 RECT 9.75 1.91 10.67 2.01 ;
 RECT 5.475 0.37 8.765 0.47 ;
 RECT 5.43 0.5 5.66 0.71 ;
 RECT 5.93 1.575 6.03 2.485 ;
 RECT 6.44 1.41 6.67 1.475 ;
 RECT 6.44 1.575 6.67 1.62 ;
 RECT 5.93 1.475 6.67 1.575 ;
 RECT 5.29 1.61 5.555 1.82 ;
 RECT 5.455 1.82 5.555 2.49 ;
 RECT 5.085 0.66 5.185 1.51 ;
 RECT 5.085 1.51 5.555 1.61 ;
 RECT 7.75 0.655 7.85 1.24 ;
 RECT 7.17 1.34 7.4 1.475 ;
 RECT 7.17 1.24 7.85 1.34 ;
 RECT 1.53 0.655 1.63 1.495 ;
 RECT 1.335 1.495 1.63 1.745 ;
 RECT 1.53 1.745 1.63 2.37 ;
 RECT 0.815 0.27 1.155 0.52 ;
 RECT 1.055 0.52 1.155 2.465 ;
 RECT 3.19 1.595 3.29 2.48 ;
 RECT 2.65 1.445 2.895 1.495 ;
 RECT 2.65 1.495 3.29 1.595 ;
 RECT 2.65 1.595 2.895 1.69 ;
 RECT 3.685 1.33 3.825 1.475 ;
 RECT 3.685 1.71 3.785 2.475 ;
 RECT 3.725 0.65 3.825 1.33 ;
 RECT 3.685 1.475 3.915 1.71 ;
 RECT 2.37 1.265 2.47 1.52 ;
 RECT 1.87 1.52 2.47 1.62 ;
 RECT 2.305 1.62 2.405 2.69 ;
 RECT 4.985 1.79 5.085 2.69 ;
 RECT 1.87 1.44 2.115 1.52 ;
 RECT 1.87 1.62 2.115 1.69 ;
 RECT 3.235 0.47 3.52 0.705 ;
 RECT 3.235 0.705 3.335 1.165 ;
 RECT 2.37 0.585 2.47 1.165 ;
 RECT 2.305 2.69 5.085 2.79 ;
 RECT 2.37 1.165 3.335 1.265 ;
 RECT 4.125 0.695 4.225 1.61 ;
 RECT 4.16 1.71 4.26 2.48 ;
 RECT 4.125 1.61 4.26 1.71 ;
 RECT 4.005 0.465 4.245 0.695 ;
 RECT 6.855 0.655 6.955 1.13 ;
 RECT 6.855 1.23 6.955 1.655 ;
 RECT 5.94 0.66 6.04 1.13 ;
 LAYER CO ;
 RECT 19.7 1.425 19.83 1.555 ;
 RECT 20.17 1.475 20.3 1.605 ;
 RECT 21.555 1.445 21.685 1.575 ;
 RECT 23.345 1.465 23.475 1.595 ;
 RECT 22.565 0.12 22.695 0.25 ;
 RECT 19.45 0.505 19.58 0.635 ;
 RECT 20.95 0.435 21.08 0.565 ;
 RECT 24.125 1.475 24.255 1.605 ;
 RECT 20.95 1.485 21.08 1.615 ;
 RECT 20.17 0.135 20.3 0.265 ;
 RECT 21.89 0.595 22.02 0.725 ;
 RECT 15.67 1.705 15.8 1.835 ;
 RECT 15.67 0.975 15.8 1.105 ;
 RECT 16.32 0.62 16.45 0.75 ;
 RECT 11.355 0.745 11.485 0.875 ;
 RECT 13.76 0.83 13.89 0.96 ;
 RECT 12.86 0.33 12.99 0.46 ;
 RECT 13.76 1.78 13.89 1.91 ;
 RECT 12.855 2.64 12.985 2.77 ;
 RECT 12.46 0.96 12.59 1.09 ;
 RECT 12.425 1.705 12.555 1.835 ;
 RECT 11.955 2.64 12.085 2.77 ;
 RECT 11.485 1.7 11.615 1.83 ;
 RECT 7.305 2.445 7.435 2.575 ;
 RECT 4.06 0.515 4.19 0.645 ;
 RECT 3.435 2.07 3.565 2.2 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 4.665 0.455 4.795 0.585 ;
 RECT 2.705 1.49 2.835 1.62 ;
 RECT 2.705 0.555 2.835 0.685 ;
 RECT 3.455 0.88 3.585 1.01 ;
 RECT 0.875 0.325 1.005 0.455 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 5.205 2.135 5.335 2.265 ;
 RECT 2.015 2.345 2.145 2.475 ;
 RECT 6.16 2.07 6.29 2.2 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.805 2.115 0.935 2.245 ;
 RECT 3.905 2.125 4.035 2.255 ;
 RECT 2.59 0.905 2.72 1.035 ;
 RECT 2.94 2.105 3.07 2.235 ;
 RECT 1.88 0.875 2.01 1.005 ;
 RECT 1.275 2.05 1.405 2.18 ;
 RECT 4.385 1.825 4.515 1.955 ;
 RECT 1.395 1.55 1.525 1.68 ;
 RECT 2.02 0.21 2.15 0.34 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 4.735 2.125 4.865 2.255 ;
 RECT 1.75 1.995 1.88 2.125 ;
 RECT 3.735 1.525 3.865 1.655 ;
 RECT 2.985 0.88 3.115 1.01 ;
 RECT 5.675 0.93 5.805 1.06 ;
 RECT 3.34 0.525 3.47 0.655 ;
 RECT 6.605 1.995 6.735 2.125 ;
 RECT 6.16 0.88 6.29 1.01 ;
 RECT 1.93 1.495 2.06 1.625 ;
 RECT 8.405 0.875 8.535 1.005 ;
 RECT 2.525 1.825 2.655 1.955 ;
 RECT 7.22 1.28 7.35 1.41 ;
 RECT 5.675 2.015 5.805 2.145 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 6.605 0.88 6.735 1.01 ;
 RECT 8.405 1.945 8.535 2.075 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 7.495 0.62 7.625 0.75 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 7.765 2.37 7.895 2.5 ;
 RECT 20.345 1.075 20.475 1.205 ;
 RECT 21.27 0.975 21.4 1.105 ;
 RECT 22.055 0.26 22.185 0.39 ;
 RECT 23.23 2.31 23.36 2.44 ;
 RECT 19.295 1.075 19.425 1.205 ;
 RECT 20.79 1.035 20.92 1.165 ;
 RECT 23.195 1.03 23.325 1.16 ;
 RECT 19.035 0.635 19.165 0.765 ;
 RECT 18.455 0.26 18.585 0.39 ;
 RECT 10.93 0.495 11.06 0.625 ;
 RECT 10.205 0.625 10.335 0.755 ;
 RECT 9.525 0.925 9.655 1.055 ;
 RECT 14.105 0.67 14.235 0.8 ;
 RECT 13.18 1.7 13.31 1.83 ;
 RECT 13.735 0.265 13.865 0.395 ;
 RECT 13.43 1.29 13.56 1.42 ;
 RECT 12.215 0.64 12.345 0.77 ;
 RECT 11.785 0.665 11.915 0.795 ;
 RECT 10.005 2.37 10.135 2.5 ;
 RECT 10.125 1.445 10.255 1.575 ;
 RECT 5.48 0.54 5.61 0.67 ;
 RECT 6.49 1.45 6.62 1.58 ;
 RECT 5.345 1.63 5.475 1.76 ;
 RECT 14.675 0.975 14.805 1.105 ;
 RECT 9.435 0.595 9.565 0.725 ;
 RECT 9.435 1.87 9.565 2 ;
 RECT 8.93 0.595 9.06 0.725 ;
 RECT 8.93 1.9 9.06 2.03 ;
 RECT 17.38 0.63 17.51 0.76 ;
 RECT 17.38 1.71 17.51 1.84 ;
 RECT 16.795 2.64 16.925 2.77 ;
 RECT 15.165 0.36 15.295 0.49 ;
 RECT 15.08 2.64 15.21 2.77 ;
 RECT 14.675 1.705 14.805 1.835 ;
 RECT 16.32 1.725 16.45 1.855 ;
 RECT 16.6 1.25 16.73 1.38 ;
 RECT 16.88 0.62 17.01 0.75 ;
 RECT 23.345 0.595 23.475 0.725 ;
 RECT 21.385 0.12 21.515 0.25 ;
 RECT 22.4 1.49 22.53 1.62 ;
 RECT 22.03 1.405 22.16 1.535 ;
 LAYER M1 ;
 RECT 3.835 2.12 4.935 2.26 ;
 RECT 4.395 1.44 4.535 1.52 ;
 RECT 3.665 1.52 4.535 1.66 ;
 RECT 5.67 0.865 5.81 1.3 ;
 RECT 4.395 1.3 5.81 1.44 ;
 RECT 5.67 1.44 5.81 2.215 ;
 RECT 3.275 1.22 3.59 1.36 ;
 RECT 3.45 0.805 3.59 1.22 ;
 RECT 3.36 1.96 3.64 2.215 ;
 RECT 3.275 1.36 3.415 1.82 ;
 RECT 3.275 1.82 4.855 1.96 ;
 RECT 4.715 1.79 4.855 1.82 ;
 RECT 5.29 1.58 5.53 1.65 ;
 RECT 5.29 1.79 5.53 1.835 ;
 RECT 4.715 1.65 5.53 1.79 ;
 RECT 6.6 1.62 6.74 1.735 ;
 RECT 6.6 1.875 6.74 2.18 ;
 RECT 6.6 0.81 6.74 1.41 ;
 RECT 6.44 1.41 6.74 1.62 ;
 RECT 6.6 1.735 7.355 1.875 ;
 RECT 7.215 1.21 7.355 1.735 ;
 RECT 1.79 1.63 1.93 1.99 ;
 RECT 1.79 1.475 2.135 1.63 ;
 RECT 1.875 0.825 2.015 1.475 ;
 RECT 1.68 1.99 1.93 2.13 ;
 RECT 21.885 0.73 22.025 1.04 ;
 RECT 22.025 1.18 22.165 1.605 ;
 RECT 21.82 0.59 22.095 0.73 ;
 RECT 23.145 0.99 23.375 1.04 ;
 RECT 21.885 1.04 23.375 1.18 ;
 RECT 23.145 1.18 23.375 1.2 ;
 RECT 22.005 0.29 22.375 0.43 ;
 RECT 22.235 0.43 22.375 0.71 ;
 RECT 22.005 0.22 22.235 0.29 ;
 RECT 23.655 0.85 23.795 1.385 ;
 RECT 23.34 1.525 23.48 1.73 ;
 RECT 22.235 0.71 23.795 0.85 ;
 RECT 23.34 0.51 23.48 0.71 ;
 RECT 23.34 1.385 23.795 1.525 ;
 RECT 21.265 1.145 21.405 1.345 ;
 RECT 20.945 1.485 21.085 1.76 ;
 RECT 21.265 0.73 21.405 0.935 ;
 RECT 20.945 0.355 21.085 0.59 ;
 RECT 20.945 1.345 21.405 1.485 ;
 RECT 21.22 0.935 21.45 1.145 ;
 RECT 20.945 0.59 21.405 0.73 ;
 RECT 19.245 1.225 19.475 1.245 ;
 RECT 19.245 1.195 19.835 1.225 ;
 RECT 19.385 1.015 19.695 1.035 ;
 RECT 19.245 1.035 19.695 1.055 ;
 RECT 19.52 0.64 19.66 1.015 ;
 RECT 19.695 1.225 19.835 1.75 ;
 RECT 19.4 0.5 19.66 0.64 ;
 RECT 20.295 1.035 20.525 1.055 ;
 RECT 20.295 1.195 20.525 1.245 ;
 RECT 19.245 1.055 20.525 1.195 ;
 RECT 18.405 0.36 18.635 0.43 ;
 RECT 19.8 0.36 19.94 0.565 ;
 RECT 18.405 0.22 19.94 0.36 ;
 RECT 20.54 0.705 20.68 0.75 ;
 RECT 20.665 0.995 20.97 1.205 ;
 RECT 20.665 0.89 20.805 0.995 ;
 RECT 20.54 0.75 20.805 0.89 ;
 RECT 19.8 0.565 20.68 0.705 ;
 RECT 14.055 0.63 14.285 0.635 ;
 RECT 14.055 0.775 14.285 0.84 ;
 RECT 15.57 0.37 15.71 0.635 ;
 RECT 14.05 0.635 15.71 0.775 ;
 RECT 16.595 0.37 16.735 1.46 ;
 RECT 15.565 0.23 16.735 0.37 ;
 RECT 9.43 0.525 9.57 0.885 ;
 RECT 9.43 1.095 9.57 2.065 ;
 RECT 9.43 0.885 9.705 1.095 ;
 RECT 7.005 2.165 7.145 2.33 ;
 RECT 6.155 2.33 7.145 2.47 ;
 RECT 7.495 1.515 7.635 2.025 ;
 RECT 7.005 2.025 7.635 2.165 ;
 RECT 6.155 0.82 6.295 2.33 ;
 RECT 8.4 0.765 8.54 1.375 ;
 RECT 8.4 1.515 8.54 2.14 ;
 RECT 8.925 0.525 9.065 1.375 ;
 RECT 8.925 1.515 9.065 2.1 ;
 RECT 7.495 1.375 9.065 1.515 ;
 RECT 10.155 0.585 11.11 0.63 ;
 RECT 10.88 0.63 11.11 0.665 ;
 RECT 10.88 0.455 11.11 0.49 ;
 RECT 10.18 0.49 11.11 0.585 ;
 RECT 10.155 0.63 10.385 0.795 ;
 RECT 11.735 0.36 11.965 0.835 ;
 RECT 12.535 0.36 12.675 0.665 ;
 RECT 11.735 0.22 12.68 0.36 ;
 RECT 13.755 0.22 13.895 0.225 ;
 RECT 13.755 0.435 13.895 0.665 ;
 RECT 12.535 0.665 13.895 0.805 ;
 RECT 13.755 0.805 13.895 1.98 ;
 RECT 13.685 0.225 13.915 0.435 ;
 RECT 3.27 0.52 3.87 0.66 ;
 RECT 3.73 0.66 3.87 1.015 ;
 RECT 5.275 0.505 5.66 0.71 ;
 RECT 5.43 0.5 5.66 0.505 ;
 RECT 3.73 1.015 5.415 1.155 ;
 RECT 5.275 0.71 5.415 1.015 ;
 RECT 2.585 0.5 2.84 0.965 ;
 RECT 2.585 1.67 2.725 1.82 ;
 RECT 2.585 1.96 2.725 2.65 ;
 RECT 2.585 0.965 2.725 1.44 ;
 RECT 2.585 1.44 2.84 1.67 ;
 RECT 2.455 1.82 2.725 1.96 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.11 ;
 RECT 0.58 2.25 0.72 2.255 ;
 RECT 0.58 0.87 1.005 1.01 ;
 RECT 0.58 2.11 1.005 2.25 ;
 RECT 0.58 1.195 1.69 1.335 ;
 RECT 1.55 0.67 1.69 1.195 ;
 RECT 2.98 0.36 3.12 2.035 ;
 RECT 2.295 0.22 3.12 0.36 ;
 RECT 1.55 0.53 2.435 0.67 ;
 RECT 2.935 2.17 3.075 2.305 ;
 RECT 2.935 2.035 3.12 2.17 ;
 RECT 2.295 0.36 2.435 0.53 ;
 RECT 9.955 2.42 10.185 2.54 ;
 RECT 18.84 2.42 18.98 2.52 ;
 RECT 9.955 2.28 18.98 2.42 ;
 RECT 23.18 2.48 23.32 2.52 ;
 RECT 18.84 2.52 23.32 2.66 ;
 RECT 23.18 2.27 23.41 2.48 ;
 RECT 11.48 1.51 11.62 1.695 ;
 RECT 11.41 1.695 11.69 1.835 ;
 RECT 12.455 1.095 12.595 1.37 ;
 RECT 12.42 1.51 12.56 1.7 ;
 RECT 13.38 1.25 13.61 1.37 ;
 RECT 11.48 1.37 13.61 1.51 ;
 RECT 12.385 0.955 12.665 1.095 ;
 RECT 12.355 1.7 12.63 1.84 ;
 RECT 10.09 2.05 10.23 2.055 ;
 RECT 10.09 1.915 11.265 1.985 ;
 RECT 10.09 1.91 11.26 1.915 ;
 RECT 10.09 1.615 10.23 1.91 ;
 RECT 13.13 1.87 13.315 1.985 ;
 RECT 10.09 1.985 13.315 2.05 ;
 RECT 11.12 2.05 13.315 2.125 ;
 RECT 13.13 1.66 13.36 1.87 ;
 RECT 10.075 1.405 10.305 1.615 ;
 END
END RDFFSRARX1

MACRO RDFFSRARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 29.44 BY 2.88 ;
 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.02 0.465 4.245 0.695 ;
 RECT 4.055 0.735 5.13 0.875 ;
 RECT 9.875 1.09 12.245 1.23 ;
 RECT 4.055 0.445 4.195 0.465 ;
 RECT 4.055 0.695 4.245 0.735 ;
 RECT 4.99 0.22 6.625 0.36 ;
 RECT 4.99 0.36 5.13 0.735 ;
 RECT 6.485 0.525 7.03 0.665 ;
 RECT 6.89 0.925 8.005 1.065 ;
 RECT 7.86 0.245 10.01 0.255 ;
 RECT 7.86 0.255 10.015 0.385 ;
 RECT 9.875 0.385 10.015 1.09 ;
 RECT 12.105 0.81 12.245 1.09 ;
 RECT 12.105 0.6 12.395 0.81 ;
 RECT 6.485 0.36 6.625 0.525 ;
 RECT 6.89 0.665 7.03 0.925 ;
 RECT 7.865 0.385 8.005 0.925 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 29.44 0.08 ;
 RECT 26.175 0.08 26.415 0.26 ;
 RECT 7.425 0.615 7.695 0.755 ;
 RECT 15.105 0.335 15.37 0.495 ;
 RECT 16.295 0.335 16.56 0.495 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 4.615 0.08 4.85 0.595 ;
 RECT 2.015 0.08 2.155 0.39 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 11.35 0.08 11.49 0.945 ;
 RECT 12.855 0.08 12.995 0.525 ;
 RECT 18.03 0.08 18.17 0.82 ;
 RECT 23.825 0.08 23.965 0.36 ;
 RECT 25.04 0.08 25.18 0.35 ;
 RECT 7.49 0.08 7.63 0.615 ;
 RECT 15.16 0.08 15.3 0.335 ;
 RECT 16.35 0.08 16.49 0.335 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 29.44 2.96 ;
 RECT 11.88 2.52 12.155 2.66 ;
 RECT 1.945 2.34 2.195 2.8 ;
 RECT 5.2 2.07 5.34 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.27 1.98 1.41 2.8 ;
 RECT 7.3 2.375 7.44 2.8 ;
 RECT 17.865 2.5 18.005 2.8 ;
 RECT 12.85 2.5 12.99 2.8 ;
 RECT 15.075 2.5 15.215 2.8 ;
 RECT 16.305 2.5 16.445 2.8 ;
 RECT 19.07 2.5 19.21 2.8 ;
 RECT 11.95 2.66 12.09 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.475 1.65 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.765 0.22 1.13 0.615 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 15.65 1.25 15.89 1.49 ;
 RECT 15.65 0.915 15.79 1.25 ;
 RECT 14.67 0.915 14.81 1.765 ;
 RECT 16.91 1.905 17.05 1.91 ;
 RECT 14.67 1.765 17.05 1.905 ;
 RECT 16.91 0.915 17.05 1.765 ;
 RECT 15.65 1.905 15.79 1.91 ;
 RECT 15.65 1.49 15.79 1.765 ;
 END
 ANTENNADIFFAREA 1.311 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.29 1.25 17.53 1.49 ;
 RECT 17.39 1.765 20.005 1.905 ;
 RECT 17.32 0.94 17.6 1.08 ;
 RECT 17.39 1.905 17.53 1.915 ;
 RECT 17.39 1.49 17.53 1.765 ;
 RECT 17.39 1.08 17.53 1.25 ;
 RECT 17.39 0.915 17.53 0.94 ;
 RECT 18.505 1.905 18.645 1.91 ;
 RECT 18.505 0.56 18.645 1.765 ;
 END
 ANTENNADIFFAREA 1.473 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.71 2.31 8.12 2.52 ;
 RECT 7.88 2.12 8.12 2.31 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 27.735 1.435 28.075 1.8 ;
 RECT 26.055 1.99 27.92 2.13 ;
 RECT 23.825 2.22 26.195 2.36 ;
 RECT 26.055 1.435 26.195 1.99 ;
 RECT 27.78 1.8 27.92 1.99 ;
 RECT 23.825 1.39 23.965 2.22 ;
 RECT 25.21 1.37 25.35 2.22 ;
 RECT 26.055 2.13 26.195 2.22 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.505 0.59 22.875 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 OBS
 LAYER PO ;
 RECT 21.85 0.19 21.95 0.235 ;
 RECT 19.475 1.43 19.575 2.565 ;
 RECT 18.785 1.43 18.885 2.565 ;
 RECT 17.65 1.43 17.92 1.435 ;
 RECT 17.65 1.435 17.75 2.57 ;
 RECT 17.65 1.33 19.575 1.43 ;
 RECT 18.29 1.43 18.39 2.565 ;
 RECT 21.94 0.36 22.17 0.445 ;
 RECT 18.29 0.09 21.95 0.19 ;
 RECT 26.785 2.27 27.07 2.48 ;
 RECT 26.785 1.2 26.885 2.27 ;
 RECT 26.785 0.375 26.885 0.99 ;
 RECT 26.785 0.99 27.035 1.2 ;
 RECT 25.3 0.38 25.4 0.96 ;
 RECT 25.3 1.06 25.4 1.14 ;
 RECT 24.88 0.935 25.11 0.96 ;
 RECT 24.88 0.96 25.4 1.06 ;
 RECT 24.88 1.06 25.11 1.145 ;
 RECT 25.3 1.14 25.57 1.24 ;
 RECT 25.47 1.24 25.57 1.84 ;
 RECT 25.665 0.22 25.895 0.28 ;
 RECT 25.665 0.38 25.895 0.43 ;
 RECT 25.3 0.28 25.895 0.38 ;
 RECT 24.39 0.215 24.49 0.995 ;
 RECT 24.39 0.995 24.63 1.205 ;
 RECT 24.39 1.205 24.49 2 ;
 RECT 27.485 0.195 27.585 2.665 ;
 RECT 26.475 0.095 27.585 0.195 ;
 RECT 22.85 1.245 22.95 2.665 ;
 RECT 22.85 1.2 23.135 1.245 ;
 RECT 26.475 0.195 26.575 0.945 ;
 RECT 22.905 1.035 23.135 1.1 ;
 RECT 22.85 2.665 27.585 2.765 ;
 RECT 22.85 1.1 23.18 1.2 ;
 RECT 23.61 0.21 23.71 0.755 ;
 RECT 23.61 0.855 23.71 2.2 ;
 RECT 26.475 1.125 26.575 2.2 ;
 RECT 22.645 0.755 24.18 0.84 ;
 RECT 22.645 0.84 24.175 0.855 ;
 RECT 24.08 0.215 24.18 0.755 ;
 RECT 22.645 0.595 22.875 0.755 ;
 RECT 23.61 2.2 26.575 2.3 ;
 RECT 24.085 1.245 24.185 2.02 ;
 RECT 23.955 1.035 24.185 1.245 ;
 RECT 10.155 0.795 10.32 0.925 ;
 RECT 9.475 0.885 9.705 0.925 ;
 RECT 9.475 1.025 9.705 1.095 ;
 RECT 9.475 0.925 10.32 1.025 ;
 RECT 10.155 0.585 10.385 0.795 ;
 RECT 13.105 1.635 13.205 1.66 ;
 RECT 13.105 1.66 13.36 1.87 ;
 RECT 13.105 1.87 13.205 2.565 ;
 RECT 14.935 0.39 15.035 1.31 ;
 RECT 14.935 1.41 15.035 2.27 ;
 RECT 15.415 0.395 15.515 1.31 ;
 RECT 15.415 1.41 15.515 2.27 ;
 RECT 13.685 0.29 15.035 0.39 ;
 RECT 16.64 0.395 16.74 1.31 ;
 RECT 16.09 0.395 16.19 1.31 ;
 RECT 14.935 1.31 16.74 1.41 ;
 RECT 16.64 1.41 16.74 2.27 ;
 RECT 16.09 1.41 16.19 2.27 ;
 RECT 13.685 0.225 13.915 0.29 ;
 RECT 13.685 0.39 13.915 0.435 ;
 RECT 13.38 1.25 13.64 1.3 ;
 RECT 13.54 0.61 13.64 1.25 ;
 RECT 13.38 1.4 13.64 1.46 ;
 RECT 13.54 1.46 13.64 2.56 ;
 RECT 14.07 0.84 14.17 1.3 ;
 RECT 13.38 1.3 14.17 1.4 ;
 RECT 14.055 0.63 14.285 0.84 ;
 RECT 12.205 0.81 12.305 2.21 ;
 RECT 12.165 0.6 12.395 0.81 ;
 RECT 10.88 0.455 11.9 0.47 ;
 RECT 10.96 0.37 11.9 0.455 ;
 RECT 10.88 0.47 11.11 0.665 ;
 RECT 11.735 0.47 11.9 0.625 ;
 RECT 11.735 0.835 11.835 2.21 ;
 RECT 11.735 0.625 11.965 0.835 ;
 RECT 8.145 2.69 10.055 2.695 ;
 RECT 9.955 2.54 10.055 2.69 ;
 RECT 8.935 2.695 10.055 2.79 ;
 RECT 8.145 0.655 8.245 2.595 ;
 RECT 8.145 2.595 9.035 2.69 ;
 RECT 9.955 2.33 10.185 2.54 ;
 RECT 9.18 0.19 9.28 1.29 ;
 RECT 2.69 0.185 9.28 0.19 ;
 RECT 10.075 1.39 10.27 1.405 ;
 RECT 2.69 0.285 2.79 0.51 ;
 RECT 2.69 0.19 4.525 0.285 ;
 RECT 4.425 0.285 4.525 1.24 ;
 RECT 4.425 0.09 9.28 0.185 ;
 RECT 9.18 1.29 10.27 1.39 ;
 RECT 2.65 0.51 2.895 0.755 ;
 RECT 10.075 1.405 10.305 1.615 ;
 RECT 5.475 0.475 5.66 0.5 ;
 RECT 13.11 0.19 13.21 1.18 ;
 RECT 10.57 0.09 13.21 0.19 ;
 RECT 10.57 0.19 10.67 1.91 ;
 RECT 9.75 1.71 9.85 1.91 ;
 RECT 8.665 0.475 8.765 1.61 ;
 RECT 8.665 1.61 9.85 1.71 ;
 RECT 8.665 1.71 8.765 1.725 ;
 RECT 9.215 1.71 9.315 2.445 ;
 RECT 9.75 1.91 10.67 2.01 ;
 RECT 5.475 0.375 8.765 0.475 ;
 RECT 5.43 0.5 5.66 0.71 ;
 RECT 5.93 1.575 6.03 2.485 ;
 RECT 6.44 1.41 6.67 1.475 ;
 RECT 6.44 1.575 6.67 1.62 ;
 RECT 5.93 1.475 6.67 1.575 ;
 RECT 7.75 0.655 7.85 1.24 ;
 RECT 7.14 1.34 7.37 1.475 ;
 RECT 7.14 1.24 7.85 1.34 ;
 RECT 1.53 0.655 1.63 1.495 ;
 RECT 1.335 1.495 1.63 1.745 ;
 RECT 1.53 1.745 1.63 2.37 ;
 RECT 0.815 0.27 1.155 0.52 ;
 RECT 1.055 0.52 1.155 2.465 ;
 RECT 3.19 1.595 3.29 2.48 ;
 RECT 2.65 1.445 2.895 1.495 ;
 RECT 2.65 1.495 3.29 1.595 ;
 RECT 2.65 1.595 2.895 1.69 ;
 RECT 3.685 1.33 3.825 1.475 ;
 RECT 3.685 1.71 3.785 2.475 ;
 RECT 3.725 0.65 3.825 1.33 ;
 RECT 3.685 1.475 3.915 1.71 ;
 RECT 2.37 1.265 2.47 1.52 ;
 RECT 1.87 1.52 2.47 1.62 ;
 RECT 2.305 1.62 2.405 2.69 ;
 RECT 4.985 1.79 5.085 2.69 ;
 RECT 1.87 1.44 2.115 1.52 ;
 RECT 1.87 1.62 2.115 1.69 ;
 RECT 3.235 0.47 3.52 0.705 ;
 RECT 3.235 0.705 3.335 1.165 ;
 RECT 2.37 0.585 2.47 1.165 ;
 RECT 2.305 2.69 5.085 2.79 ;
 RECT 2.37 1.165 3.335 1.265 ;
 RECT 4.125 0.695 4.225 1.61 ;
 RECT 4.16 1.71 4.26 2.48 ;
 RECT 4.125 1.61 4.26 1.71 ;
 RECT 4.005 0.465 4.245 0.695 ;
 RECT 5.29 1.61 5.555 1.82 ;
 RECT 5.455 1.82 5.555 2.49 ;
 RECT 5.085 0.66 5.185 1.51 ;
 RECT 5.085 1.51 5.555 1.61 ;
 RECT 6.855 0.655 6.955 1.13 ;
 RECT 6.855 1.23 6.955 1.655 ;
 RECT 5.94 0.66 6.04 1.13 ;
 RECT 6.855 1.655 7.815 1.755 ;
 RECT 7.715 1.755 7.815 2.31 ;
 RECT 6.855 1.755 6.955 2.57 ;
 RECT 5.94 1.13 6.955 1.23 ;
 RECT 7.71 2.31 7.94 2.52 ;
 RECT 21.85 0.235 22.17 0.36 ;
 RECT 17.65 0.4 17.75 1.2 ;
 RECT 17.65 1.2 17.92 1.33 ;
 RECT 18.29 0.19 18.39 1.33 ;
 LAYER CO ;
 RECT 13.76 0.83 13.89 0.96 ;
 RECT 12.86 0.33 12.99 0.46 ;
 RECT 13.76 1.78 13.89 1.91 ;
 RECT 12.855 2.57 12.985 2.7 ;
 RECT 12.46 0.96 12.59 1.09 ;
 RECT 12.425 1.665 12.555 1.795 ;
 RECT 11.955 2.525 12.085 2.655 ;
 RECT 11.485 1.665 11.615 1.795 ;
 RECT 7.305 2.445 7.435 2.575 ;
 RECT 2.015 2.345 2.145 2.475 ;
 RECT 6.16 2.07 6.29 2.2 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.805 2.115 0.935 2.245 ;
 RECT 3.905 2.125 4.035 2.255 ;
 RECT 2.59 0.905 2.72 1.035 ;
 RECT 2.94 2.105 3.07 2.235 ;
 RECT 1.88 0.875 2.01 1.005 ;
 RECT 1.275 2.05 1.405 2.18 ;
 RECT 4.385 1.825 4.515 1.955 ;
 RECT 1.395 1.55 1.525 1.68 ;
 RECT 2.02 0.21 2.15 0.34 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 4.735 2.125 4.865 2.255 ;
 RECT 1.75 1.995 1.88 2.125 ;
 RECT 3.735 1.525 3.865 1.655 ;
 RECT 2.985 0.88 3.115 1.01 ;
 RECT 5.675 0.93 5.805 1.06 ;
 RECT 3.34 0.525 3.47 0.655 ;
 RECT 6.605 1.995 6.735 2.125 ;
 RECT 6.16 0.88 6.29 1.01 ;
 RECT 1.93 1.495 2.06 1.625 ;
 RECT 8.405 0.875 8.535 1.005 ;
 RECT 5.345 1.63 5.475 1.76 ;
 RECT 14.675 0.975 14.805 1.105 ;
 RECT 9.435 0.595 9.565 0.725 ;
 RECT 9.435 1.87 9.565 2 ;
 RECT 8.93 0.595 9.06 0.725 ;
 RECT 8.93 1.9 9.06 2.03 ;
 RECT 2.525 1.825 2.655 1.955 ;
 RECT 7.19 1.28 7.32 1.41 ;
 RECT 5.675 2.015 5.805 2.145 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 6.605 0.88 6.735 1.01 ;
 RECT 8.405 1.945 8.535 2.075 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 7.495 0.62 7.625 0.75 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 4.06 0.515 4.19 0.645 ;
 RECT 3.435 2.07 3.565 2.2 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 4.665 0.455 4.795 0.585 ;
 RECT 2.705 1.49 2.835 1.62 ;
 RECT 2.705 0.555 2.835 0.685 ;
 RECT 3.455 0.88 3.585 1.01 ;
 RECT 0.875 0.325 1.005 0.455 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 5.205 2.135 5.335 2.265 ;
 RECT 7.76 2.35 7.89 2.48 ;
 RECT 21.99 0.275 22.12 0.405 ;
 RECT 26.89 2.31 27.02 2.44 ;
 RECT 24.93 0.975 25.06 1.105 ;
 RECT 26.855 1.03 26.985 1.16 ;
 RECT 25.715 0.26 25.845 0.39 ;
 RECT 24.45 1.035 24.58 1.165 ;
 RECT 22.955 1.075 23.085 1.205 ;
 RECT 22.695 0.635 22.825 0.765 ;
 RECT 24.005 1.075 24.135 1.205 ;
 RECT 10.93 0.495 11.06 0.625 ;
 RECT 10.205 0.625 10.335 0.755 ;
 RECT 9.525 0.925 9.655 1.055 ;
 RECT 14.105 0.67 14.235 0.8 ;
 RECT 13.18 1.7 13.31 1.83 ;
 RECT 13.735 0.265 13.865 0.395 ;
 RECT 13.43 1.29 13.56 1.42 ;
 RECT 12.215 0.64 12.345 0.77 ;
 RECT 11.785 0.665 11.915 0.795 ;
 RECT 10.005 2.37 10.135 2.5 ;
 RECT 10.125 1.445 10.255 1.575 ;
 RECT 5.48 0.54 5.61 0.67 ;
 RECT 6.49 1.45 6.62 1.58 ;
 RECT 23.36 1.425 23.49 1.555 ;
 RECT 25.69 1.405 25.82 1.535 ;
 RECT 27.785 1.475 27.915 1.605 ;
 RECT 27.005 0.595 27.135 0.725 ;
 RECT 23.83 1.475 23.96 1.605 ;
 RECT 26.225 0.12 26.355 0.25 ;
 RECT 27.005 1.465 27.135 1.595 ;
 RECT 26.06 1.49 26.19 1.62 ;
 RECT 25.55 0.595 25.68 0.725 ;
 RECT 23.83 0.135 23.96 0.265 ;
 RECT 25.215 1.445 25.345 1.575 ;
 RECT 24.61 1.485 24.74 1.615 ;
 RECT 24.61 0.435 24.74 0.565 ;
 RECT 23.11 0.505 23.24 0.635 ;
 RECT 25.045 0.12 25.175 0.25 ;
 RECT 18.51 0.63 18.64 0.76 ;
 RECT 18.51 1.71 18.64 1.84 ;
 RECT 17.87 2.57 18 2.7 ;
 RECT 15.165 0.36 15.295 0.49 ;
 RECT 15.655 0.97 15.785 1.1 ;
 RECT 15.655 1.705 15.785 1.835 ;
 RECT 14.675 1.705 14.805 1.835 ;
 RECT 17.395 1.725 17.525 1.855 ;
 RECT 17.75 1.25 17.88 1.38 ;
 RECT 18.035 0.62 18.165 0.75 ;
 RECT 19.79 1.77 19.92 1.9 ;
 RECT 16.915 0.97 17.045 1.1 ;
 RECT 16.915 1.705 17.045 1.835 ;
 RECT 19.075 2.57 19.205 2.7 ;
 RECT 16.355 0.36 16.485 0.49 ;
 RECT 16.31 2.57 16.44 2.7 ;
 RECT 15.08 2.57 15.21 2.7 ;
 RECT 17.395 0.95 17.525 1.08 ;
 RECT 11.355 0.745 11.485 0.875 ;
 LAYER M1 ;
 RECT 4.395 1.44 4.535 1.52 ;
 RECT 3.665 1.52 4.535 1.66 ;
 RECT 5.67 0.865 5.81 1.3 ;
 RECT 4.395 1.3 5.81 1.44 ;
 RECT 5.67 1.44 5.81 2.215 ;
 RECT 1.79 1.63 1.93 1.99 ;
 RECT 1.79 1.475 2.135 1.63 ;
 RECT 1.875 0.825 2.015 1.475 ;
 RECT 1.68 1.99 1.93 2.13 ;
 RECT 3.275 1.22 3.59 1.36 ;
 RECT 3.45 0.805 3.59 1.22 ;
 RECT 3.36 1.96 3.64 2.215 ;
 RECT 3.275 1.36 3.415 1.82 ;
 RECT 3.275 1.82 4.855 1.96 ;
 RECT 4.715 1.79 4.855 1.82 ;
 RECT 5.29 1.58 5.53 1.65 ;
 RECT 5.29 1.79 5.53 1.835 ;
 RECT 4.715 1.65 5.53 1.79 ;
 RECT 6.6 1.62 6.74 1.735 ;
 RECT 6.6 1.875 6.74 2.18 ;
 RECT 6.6 0.81 6.74 1.41 ;
 RECT 6.44 1.41 6.74 1.62 ;
 RECT 6.6 1.735 7.325 1.875 ;
 RECT 7.185 1.21 7.325 1.735 ;
 RECT 25.545 0.73 25.685 1.04 ;
 RECT 25.685 1.18 25.825 1.605 ;
 RECT 25.48 0.59 25.755 0.73 ;
 RECT 26.805 0.99 27.035 1.04 ;
 RECT 25.545 1.04 27.035 1.18 ;
 RECT 26.805 1.18 27.035 1.2 ;
 RECT 24.925 1.145 25.065 1.345 ;
 RECT 24.605 1.485 24.745 1.76 ;
 RECT 24.925 0.73 25.065 0.935 ;
 RECT 24.605 0.355 24.745 0.59 ;
 RECT 24.605 1.345 25.065 1.485 ;
 RECT 24.88 0.935 25.11 1.145 ;
 RECT 24.605 0.59 25.065 0.73 ;
 RECT 22.905 1.225 23.135 1.245 ;
 RECT 22.905 1.195 23.495 1.225 ;
 RECT 23.045 1.015 23.355 1.035 ;
 RECT 22.905 1.035 23.355 1.055 ;
 RECT 23.18 0.64 23.32 1.015 ;
 RECT 23.355 1.225 23.495 1.75 ;
 RECT 23.06 0.5 23.32 0.64 ;
 RECT 23.955 1.035 24.185 1.055 ;
 RECT 23.955 1.195 24.185 1.245 ;
 RECT 22.905 1.055 24.185 1.195 ;
 RECT 21.94 0.36 22.17 0.445 ;
 RECT 23.46 0.36 23.6 0.565 ;
 RECT 21.94 0.235 23.6 0.36 ;
 RECT 22.065 0.22 23.6 0.235 ;
 RECT 24.2 0.705 24.34 0.75 ;
 RECT 24.325 0.995 24.63 1.205 ;
 RECT 24.325 0.89 24.465 0.995 ;
 RECT 24.2 0.75 24.465 0.89 ;
 RECT 23.46 0.565 24.34 0.705 ;
 RECT 25.665 0.29 26.035 0.43 ;
 RECT 25.895 0.43 26.035 0.71 ;
 RECT 25.665 0.22 25.895 0.29 ;
 RECT 27.315 0.85 27.455 1.385 ;
 RECT 27 1.525 27.14 1.73 ;
 RECT 25.895 0.71 27.455 0.85 ;
 RECT 27 0.51 27.14 0.71 ;
 RECT 27 1.385 27.455 1.525 ;
 RECT 10.155 0.585 11.11 0.63 ;
 RECT 10.88 0.63 11.11 0.665 ;
 RECT 10.88 0.455 11.11 0.49 ;
 RECT 10.18 0.49 11.11 0.585 ;
 RECT 10.155 0.63 10.385 0.795 ;
 RECT 14.055 0.63 14.285 0.635 ;
 RECT 14.055 0.775 14.285 0.84 ;
 RECT 17.745 0.775 17.885 1.46 ;
 RECT 14.05 0.635 17.885 0.775 ;
 RECT 11.735 0.36 11.965 0.835 ;
 RECT 12.535 0.36 12.675 0.665 ;
 RECT 11.735 0.22 12.68 0.36 ;
 RECT 13.755 0.22 13.895 0.225 ;
 RECT 13.755 0.435 13.895 0.665 ;
 RECT 12.535 0.665 13.895 0.805 ;
 RECT 13.755 0.805 13.895 1.98 ;
 RECT 13.685 0.225 13.915 0.435 ;
 RECT 7.005 2.165 7.145 2.33 ;
 RECT 7.005 2.47 7.145 2.475 ;
 RECT 6.155 2.33 7.145 2.47 ;
 RECT 7.465 1.65 7.605 2.025 ;
 RECT 7.005 2.025 7.605 2.165 ;
 RECT 6.155 0.82 6.295 2.33 ;
 RECT 6.155 2.47 6.295 2.475 ;
 RECT 8.4 0.765 8.54 1.51 ;
 RECT 8.4 1.65 8.54 2.145 ;
 RECT 8.925 0.525 9.065 1.51 ;
 RECT 8.925 1.65 9.065 2.1 ;
 RECT 7.465 1.51 9.065 1.65 ;
 RECT 2.585 0.5 2.84 0.965 ;
 RECT 2.585 1.67 2.725 1.82 ;
 RECT 2.585 1.96 2.725 2.65 ;
 RECT 2.585 0.965 2.725 1.44 ;
 RECT 2.585 1.44 2.84 1.67 ;
 RECT 2.455 1.82 2.725 1.96 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.11 ;
 RECT 0.58 2.25 0.72 2.255 ;
 RECT 0.58 0.87 1.005 1.01 ;
 RECT 0.58 2.11 1.005 2.25 ;
 RECT 0.58 1.195 1.69 1.335 ;
 RECT 1.55 0.67 1.69 1.195 ;
 RECT 2.98 0.36 3.12 2.035 ;
 RECT 2.295 0.22 3.12 0.36 ;
 RECT 1.55 0.53 2.435 0.67 ;
 RECT 2.935 2.17 3.075 2.305 ;
 RECT 2.935 2.035 3.12 2.17 ;
 RECT 2.295 0.36 2.435 0.53 ;
 RECT 9.43 0.525 9.57 0.885 ;
 RECT 9.43 1.095 9.57 2.065 ;
 RECT 9.43 0.885 9.705 1.095 ;
 RECT 3.27 0.52 3.87 0.66 ;
 RECT 3.73 0.66 3.87 1.015 ;
 RECT 5.275 0.505 5.66 0.71 ;
 RECT 5.43 0.5 5.66 0.505 ;
 RECT 3.73 1.015 5.415 1.155 ;
 RECT 5.275 0.71 5.415 1.015 ;
 RECT 9.955 2.36 10.185 2.54 ;
 RECT 22.5 2.36 22.64 2.52 ;
 RECT 9.955 2.22 22.64 2.36 ;
 RECT 26.84 2.48 26.98 2.52 ;
 RECT 22.5 2.52 26.98 2.66 ;
 RECT 26.84 2.27 27.07 2.48 ;
 RECT 11.48 1.51 11.62 1.66 ;
 RECT 11.41 1.66 11.69 1.8 ;
 RECT 12.455 1.095 12.595 1.37 ;
 RECT 12.42 1.51 12.56 1.66 ;
 RECT 11.48 1.37 13.61 1.51 ;
 RECT 13.38 1.25 13.61 1.37 ;
 RECT 12.385 0.955 12.665 1.095 ;
 RECT 12.355 1.66 12.63 1.8 ;
 RECT 13.13 1.87 13.315 1.94 ;
 RECT 10.09 1.615 10.23 1.91 ;
 RECT 10.09 1.94 13.315 2.05 ;
 RECT 10.09 1.91 11.26 1.94 ;
 RECT 11.125 2.05 13.315 2.08 ;
 RECT 13.13 1.66 13.36 1.87 ;
 RECT 10.075 1.405 10.305 1.615 ;
 RECT 3.835 2.12 4.935 2.26 ;
 END
END RDFFSRARX2

MACRO RDFFSRASRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.84 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.93 0.59 21.3 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.16 1.435 26.5 1.8 ;
 RECT 24.48 1.99 26.345 2.13 ;
 RECT 22.25 2.22 24.62 2.36 ;
 RECT 26.205 1.8 26.345 1.99 ;
 RECT 24.48 1.435 24.62 1.99 ;
 RECT 22.25 1.39 22.39 2.22 ;
 RECT 23.635 1.37 23.775 2.22 ;
 RECT 24.48 2.13 24.62 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.77 0.22 1.135 0.525 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.86 0.08 2.14 0.295 ;
 RECT 24.6 0.08 24.84 0.26 ;
 RECT 5.79 0.31 6.08 0.45 ;
 RECT 9.475 0.615 9.745 0.755 ;
 RECT 13.4 0.275 14.425 0.415 ;
 RECT 17.76 0.335 18.025 0.495 ;
 RECT 14.285 0.75 15.23 0.89 ;
 RECT 0 -0.08 27.84 0.08 ;
 RECT 1.275 0.08 1.415 0.97 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.685 0.08 4.92 0.46 ;
 RECT 19.405 0.08 19.545 0.82 ;
 RECT 22.25 0.08 22.39 0.36 ;
 RECT 23.465 0.08 23.605 0.35 ;
 RECT 5.87 0.08 6.01 0.31 ;
 RECT 9.54 0.08 9.68 0.615 ;
 RECT 13.4 0.415 13.54 0.945 ;
 RECT 13.4 0.08 13.54 0.275 ;
 RECT 17.815 0.08 17.955 0.335 ;
 RECT 15.09 0.89 15.23 1.11 ;
 RECT 14.285 0.415 14.425 0.75 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.215 1.205 17.465 1.445 ;
 RECT 17.325 0.915 17.465 1.205 ;
 RECT 18.33 1.84 18.47 1.885 ;
 RECT 18.33 0.915 18.47 1.7 ;
 RECT 17.325 1.84 17.465 1.885 ;
 RECT 17.325 1.7 18.47 1.84 ;
 RECT 17.325 1.445 17.465 1.7 ;
 END
 ANTENNADIFFAREA 0.7 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 17.67 2.6 17.935 2.8 ;
 RECT 19.26 2.6 19.525 2.8 ;
 RECT 9.285 2.215 9.56 2.355 ;
 RECT 0 2.8 27.84 2.96 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.275 1.98 1.415 2.8 ;
 RECT 2.015 2.34 2.265 2.8 ;
 RECT 5.87 1.98 6.01 2.8 ;
 RECT 5.39 2.07 5.53 2.8 ;
 RECT 6.9 2 7.04 2.8 ;
 RECT 12.31 2.335 12.58 2.8 ;
 RECT 9.35 2.355 9.49 2.8 ;
 RECT 9.35 2.195 9.49 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.325 1.475 1.655 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.725 1.095 18.985 1.335 ;
 RECT 18.845 0.51 18.985 1.095 ;
 RECT 19.905 1.905 20.045 1.91 ;
 RECT 18.845 1.765 20.045 1.905 ;
 RECT 19.905 0.56 20.045 1.765 ;
 RECT 18.845 1.905 18.985 1.915 ;
 RECT 18.845 1.335 18.985 1.765 ;
 END
 ANTENNADIFFAREA 0.568 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.765 2.255 10.09 2.465 ;
 RECT 9.82 2.12 10.09 2.255 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.08 0.485 4.395 0.605 ;
 RECT 9 0.905 10.055 1.045 ;
 RECT 9.915 0.245 12.06 0.255 ;
 RECT 9.915 0.255 12.065 0.385 ;
 RECT 11.925 1.09 13.915 1.23 ;
 RECT 14.12 1.56 14.35 1.6 ;
 RECT 13.775 1.42 14.35 1.56 ;
 RECT 14.12 1.39 14.35 1.42 ;
 RECT 4.08 0.605 9.14 0.745 ;
 RECT 9 0.745 9.14 0.905 ;
 RECT 9.915 0.385 10.055 0.905 ;
 RECT 11.925 0.385 12.065 1.09 ;
 RECT 13.775 1.23 13.915 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.24 1.795 7.48 2.04 ;
 RECT 6.69 1.795 6.92 1.83 ;
 RECT 6.69 1.655 7.48 1.795 ;
 RECT 6.69 1.62 6.92 1.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 OBS
 LAYER PO ;
 RECT 19.105 0.385 19.205 1.25 ;
 RECT 19.105 1.46 19.205 2.575 ;
 RECT 19.685 1.43 19.785 2.575 ;
 RECT 20.29 0.22 20.52 0.275 ;
 RECT 20.29 0.375 20.52 0.43 ;
 RECT 19.685 0.275 20.52 0.375 ;
 RECT 14.255 0.73 14.355 1.39 ;
 RECT 14.12 1.39 14.355 1.6 ;
 RECT 14.255 1.6 14.355 2.39 ;
 RECT 11.23 0.195 11.33 1.29 ;
 RECT 12.125 1.39 12.32 1.405 ;
 RECT 2.785 0.285 2.885 0.505 ;
 RECT 4.495 0.285 4.595 1.24 ;
 RECT 2.785 0.185 11.33 0.195 ;
 RECT 2.785 0.195 4.595 0.285 ;
 RECT 4.495 0.095 11.33 0.185 ;
 RECT 11.23 1.29 12.32 1.39 ;
 RECT 2.67 0.505 2.9 0.715 ;
 RECT 12.125 1.405 12.355 1.615 ;
 RECT 22.51 1.245 22.61 2.02 ;
 RECT 22.38 1.035 22.61 1.245 ;
 RECT 12.62 0.105 15.445 0.205 ;
 RECT 12.62 0.205 12.72 1.91 ;
 RECT 15.345 0.205 15.445 1.265 ;
 RECT 11.8 1.71 11.9 1.91 ;
 RECT 10.715 1.61 11.9 1.71 ;
 RECT 10.715 0.475 10.815 1.61 ;
 RECT 11.265 1.71 11.365 2.425 ;
 RECT 7.38 0.475 7.48 0.885 ;
 RECT 11.8 1.91 12.72 2.01 ;
 RECT 7.38 0.375 10.815 0.475 ;
 RECT 7.255 0.885 7.485 1.095 ;
 RECT 12.93 0.455 14.86 0.535 ;
 RECT 14.63 0.535 14.86 0.6 ;
 RECT 14.63 0.39 14.86 0.435 ;
 RECT 13.01 0.435 14.86 0.455 ;
 RECT 12.93 0.535 13.16 0.665 ;
 RECT 13.785 0.535 14.015 0.835 ;
 RECT 13.785 0.835 13.885 2.39 ;
 RECT 22.815 0.215 22.915 0.995 ;
 RECT 22.815 0.995 23.055 1.205 ;
 RECT 22.815 1.205 22.915 2 ;
 RECT 25.21 0.375 25.31 0.99 ;
 RECT 25.21 0.99 25.46 1.2 ;
 RECT 25.21 1.2 25.31 2.27 ;
 RECT 25.21 2.27 25.495 2.48 ;
 RECT 10.195 0.655 10.295 2.305 ;
 RECT 10.5 2.3 10.73 2.305 ;
 RECT 10.5 2.405 10.73 2.51 ;
 RECT 10.195 2.305 10.73 2.405 ;
 RECT 22.035 0.21 22.135 0.755 ;
 RECT 22.035 0.855 22.135 2.2 ;
 RECT 24.9 1.125 25 2.2 ;
 RECT 21.07 0.755 22.605 0.84 ;
 RECT 21.07 0.84 22.6 0.855 ;
 RECT 22.505 0.215 22.605 0.755 ;
 RECT 21.07 0.595 21.3 0.755 ;
 RECT 22.035 2.2 25 2.3 ;
 RECT 23.725 1.06 23.825 1.14 ;
 RECT 23.725 0.38 23.825 0.96 ;
 RECT 23.725 1.14 23.995 1.24 ;
 RECT 23.895 1.24 23.995 1.84 ;
 RECT 23.305 0.935 23.535 0.96 ;
 RECT 23.305 0.96 23.825 1.06 ;
 RECT 23.305 1.06 23.535 1.145 ;
 RECT 24.09 0.22 24.32 0.28 ;
 RECT 24.09 0.38 24.32 0.43 ;
 RECT 23.725 0.28 24.32 0.38 ;
 RECT 7.98 1.575 8.08 2.485 ;
 RECT 8.49 1.575 8.72 1.685 ;
 RECT 7.98 1.475 8.72 1.575 ;
 RECT 25.91 0.195 26.01 2.665 ;
 RECT 24.9 0.095 26.01 0.195 ;
 RECT 21.275 1.245 21.375 2.665 ;
 RECT 24.9 0.195 25 0.945 ;
 RECT 21.275 1.2 21.56 1.245 ;
 RECT 21.33 1.035 21.56 1.1 ;
 RECT 21.275 2.665 26.01 2.765 ;
 RECT 21.275 1.1 21.605 1.2 ;
 RECT 12.205 0.795 12.37 0.925 ;
 RECT 11.525 0.885 11.755 0.925 ;
 RECT 11.525 1.025 11.755 1.095 ;
 RECT 11.525 0.925 12.37 1.025 ;
 RECT 12.205 0.585 12.435 0.795 ;
 RECT 4.195 0.715 4.295 1.61 ;
 RECT 4.23 1.71 4.33 2.48 ;
 RECT 4.195 1.61 4.33 1.71 ;
 RECT 4.075 0.485 4.315 0.715 ;
 RECT 3.26 1.665 3.36 2.49 ;
 RECT 2.72 1.445 2.965 1.565 ;
 RECT 2.72 1.565 3.36 1.665 ;
 RECT 2.72 1.665 2.965 1.69 ;
 RECT 2.375 1.62 2.475 2.675 ;
 RECT 3.305 0.47 3.59 0.705 ;
 RECT 3.305 0.705 3.405 1.155 ;
 RECT 2.39 0.715 2.49 1.155 ;
 RECT 2.39 1.155 3.405 1.255 ;
 RECT 2.39 1.255 2.49 1.52 ;
 RECT 1.815 1.44 2.06 1.52 ;
 RECT 1.815 1.52 2.49 1.62 ;
 RECT 1.815 1.62 2.06 1.69 ;
 RECT 5.175 1.79 5.275 2.675 ;
 RECT 2.375 2.675 5.275 2.775 ;
 RECT 9.8 0.655 9.9 1.24 ;
 RECT 9.185 1.34 9.415 1.475 ;
 RECT 9.185 1.24 9.9 1.34 ;
 RECT 1.535 0.49 1.635 1.495 ;
 RECT 1.34 1.495 1.635 1.745 ;
 RECT 1.535 1.745 1.635 2.37 ;
 RECT 3.755 1.33 3.895 1.475 ;
 RECT 3.755 1.71 3.855 2.475 ;
 RECT 3.795 0.65 3.895 1.33 ;
 RECT 3.755 1.475 3.985 1.71 ;
 RECT 1.06 0.52 1.16 2.465 ;
 RECT 0.82 0.27 1.16 0.52 ;
 RECT 8.905 0.655 9.005 1.18 ;
 RECT 8.905 1.28 9.005 1.655 ;
 RECT 7.99 0.66 8.09 1.18 ;
 RECT 8.905 1.655 9.865 1.755 ;
 RECT 9.765 1.755 9.865 2.255 ;
 RECT 8.905 1.755 9.005 2.51 ;
 RECT 7.99 1.18 9.005 1.28 ;
 RECT 9.765 2.255 9.995 2.465 ;
 RECT 16.225 0.77 16.325 2.155 ;
 RECT 16.225 0.55 16.325 0.56 ;
 RECT 16.225 0.56 16.48 0.77 ;
 RECT 16.86 0.43 16.96 1.245 ;
 RECT 17.59 0.39 17.69 1.4 ;
 RECT 17.59 1.5 17.69 2.37 ;
 RECT 18.08 0.51 18.18 1.4 ;
 RECT 18.08 1.5 18.18 2.37 ;
 RECT 16.795 0.22 17.025 0.29 ;
 RECT 16.795 0.39 17.025 0.43 ;
 RECT 16.795 0.29 17.69 0.39 ;
 RECT 17.59 1.4 18.18 1.5 ;
 RECT 16.81 1.245 17.04 1.455 ;
 RECT 15.285 1.445 15.385 2.035 ;
 RECT 15.27 2.035 15.5 2.245 ;
 RECT 15.755 0.55 15.855 2.69 ;
 RECT 6.685 1.58 6.785 1.62 ;
 RECT 6.425 1.01 6.525 1.48 ;
 RECT 6.685 1.83 6.785 2.69 ;
 RECT 6.685 1.62 6.92 1.83 ;
 RECT 6.425 1.48 6.785 1.58 ;
 RECT 6.685 2.69 15.855 2.79 ;
 RECT 6.125 0.98 6.225 1.615 ;
 RECT 5.985 1.615 6.225 1.825 ;
 RECT 6.125 1.825 6.225 2.51 ;
 RECT 19.105 1.33 19.785 1.43 ;
 RECT 19.105 1.43 19.355 1.46 ;
 RECT 19.105 1.25 19.355 1.33 ;
 RECT 19.685 0.27 19.785 0.275 ;
 RECT 19.685 0.375 19.785 1.33 ;
 LAYER CO ;
 RECT 16.45 1.705 16.58 1.835 ;
 RECT 17.735 2.64 17.865 2.77 ;
 RECT 24.115 1.405 24.245 1.535 ;
 RECT 7.735 0.905 7.865 1.035 ;
 RECT 0.88 0.325 1.01 0.455 ;
 RECT 5.875 0.315 6.005 0.445 ;
 RECT 8.21 0.905 8.34 1.035 ;
 RECT 11.485 0.595 11.615 0.725 ;
 RECT 9.545 0.62 9.675 0.75 ;
 RECT 23.64 1.445 23.77 1.575 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 14.51 1.035 14.64 1.165 ;
 RECT 15.095 0.91 15.225 1.04 ;
 RECT 6.905 2.11 7.035 2.24 ;
 RECT 19.41 0.62 19.54 0.75 ;
 RECT 5.395 2.135 5.525 2.265 ;
 RECT 3.01 2.105 3.14 2.235 ;
 RECT 3.975 2.11 4.105 2.24 ;
 RECT 1.95 0.145 2.08 0.275 ;
 RECT 10.98 1.9 11.11 2.03 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 2.085 2.345 2.215 2.475 ;
 RECT 23.035 0.435 23.165 0.565 ;
 RECT 17.33 1.705 17.46 1.835 ;
 RECT 6.755 1.23 6.885 1.36 ;
 RECT 15.505 1.705 15.635 1.835 ;
 RECT 5.875 2.075 6.005 2.205 ;
 RECT 3.525 0.88 3.655 1.01 ;
 RECT 13.535 1.835 13.665 1.965 ;
 RECT 13.405 0.765 13.535 0.895 ;
 RECT 9.815 2.295 9.945 2.425 ;
 RECT 2.72 0.545 2.85 0.675 ;
 RECT 19.175 1.29 19.305 1.42 ;
 RECT 16.86 1.285 16.99 1.415 ;
 RECT 14.68 0.43 14.81 0.56 ;
 RECT 16.3 0.6 16.43 0.73 ;
 RECT 16.845 0.26 16.975 0.39 ;
 RECT 15.32 2.075 15.45 2.205 ;
 RECT 6.74 1.66 6.87 1.79 ;
 RECT 6.035 1.655 6.165 1.785 ;
 RECT 20.34 0.26 20.47 0.39 ;
 RECT 25.28 1.03 25.41 1.16 ;
 RECT 12.98 0.495 13.11 0.625 ;
 RECT 14.17 1.43 14.3 1.56 ;
 RECT 12.255 0.625 12.385 0.755 ;
 RECT 12.175 1.445 12.305 1.575 ;
 RECT 22.43 1.075 22.56 1.205 ;
 RECT 7.305 0.925 7.435 1.055 ;
 RECT 23.355 0.975 23.485 1.105 ;
 RECT 13.835 0.665 13.965 0.795 ;
 RECT 22.875 1.035 23.005 1.165 ;
 RECT 25.315 2.31 25.445 2.44 ;
 RECT 10.55 2.34 10.68 2.47 ;
 RECT 21.12 0.635 21.25 0.765 ;
 RECT 24.14 0.26 24.27 0.39 ;
 RECT 8.54 1.515 8.67 1.645 ;
 RECT 21.38 1.075 21.51 1.205 ;
 RECT 11.575 0.925 11.705 1.055 ;
 RECT 3.055 0.88 3.185 1.01 ;
 RECT 11.485 1.87 11.615 2 ;
 RECT 4.925 2.11 5.055 2.24 ;
 RECT 4.74 0.32 4.87 0.45 ;
 RECT 22.255 0.135 22.385 0.265 ;
 RECT 1.875 1.495 2.005 1.625 ;
 RECT 1.88 0.975 2.01 1.105 ;
 RECT 1.755 1.995 1.885 2.125 ;
 RECT 8.655 1.995 8.785 2.125 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 8.21 2.07 8.34 2.2 ;
 RECT 10.98 0.595 11.11 0.725 ;
 RECT 2.775 1.49 2.905 1.62 ;
 RECT 9.235 1.28 9.365 1.41 ;
 RECT 18.85 1.725 18.98 1.855 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 6.415 2.045 6.545 2.175 ;
 RECT 1.4 1.55 1.53 1.68 ;
 RECT 1.28 0.74 1.41 0.87 ;
 RECT 24.65 0.12 24.78 0.25 ;
 RECT 4.13 0.53 4.26 0.66 ;
 RECT 18.85 0.62 18.98 0.75 ;
 RECT 12.38 2.38 12.51 2.51 ;
 RECT 8.655 0.905 8.785 1.035 ;
 RECT 21.785 1.425 21.915 1.555 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 16.57 0.92 16.7 1.05 ;
 RECT 22.255 1.475 22.385 1.605 ;
 RECT 10.455 0.875 10.585 1.005 ;
 RECT 2.66 0.935 2.79 1.065 ;
 RECT 14.475 1.835 14.605 1.965 ;
 RECT 3.505 2.07 3.635 2.2 ;
 RECT 26.21 1.475 26.34 1.605 ;
 RECT 18.335 1.705 18.465 1.835 ;
 RECT 19.91 1.71 20.04 1.84 ;
 RECT 17.33 0.975 17.46 1.105 ;
 RECT 0.81 0.74 0.94 0.87 ;
 RECT 2.595 1.825 2.725 1.955 ;
 RECT 10.455 1.945 10.585 2.075 ;
 RECT 1.28 2.05 1.41 2.18 ;
 RECT 21.535 0.505 21.665 0.635 ;
 RECT 7.73 2.015 7.86 2.145 ;
 RECT 23.47 0.12 23.6 0.25 ;
 RECT 23.035 1.485 23.165 1.615 ;
 RECT 25.43 1.465 25.56 1.595 ;
 RECT 15.975 1.705 16.105 1.835 ;
 RECT 25.43 0.595 25.56 0.725 ;
 RECT 3.805 1.525 3.935 1.655 ;
 RECT 9.355 2.225 9.485 2.355 ;
 RECT 18.335 0.975 18.465 1.105 ;
 RECT 19.325 2.64 19.455 2.77 ;
 RECT 0.81 2.115 0.94 2.245 ;
 RECT 17.82 0.36 17.95 0.49 ;
 RECT 19.91 0.63 20.04 0.76 ;
 RECT 23.975 0.595 24.105 0.725 ;
 RECT 3.41 0.525 3.54 0.655 ;
 RECT 4.455 1.825 4.585 1.955 ;
 RECT 24.485 1.49 24.615 1.62 ;
 LAYER M1 ;
 RECT 1.685 1.99 1.935 2.13 ;
 RECT 23.97 0.73 24.11 1.04 ;
 RECT 24.11 1.18 24.25 1.605 ;
 RECT 23.905 0.59 24.18 0.73 ;
 RECT 25.23 0.99 25.46 1.04 ;
 RECT 23.97 1.04 25.46 1.18 ;
 RECT 25.23 1.18 25.46 1.2 ;
 RECT 24.09 0.29 24.46 0.43 ;
 RECT 24.32 0.43 24.46 0.71 ;
 RECT 24.09 0.22 24.32 0.29 ;
 RECT 25.74 0.85 25.88 1.385 ;
 RECT 25.425 1.525 25.565 1.73 ;
 RECT 24.32 0.71 25.88 0.85 ;
 RECT 25.425 0.51 25.565 0.71 ;
 RECT 25.425 1.385 25.88 1.525 ;
 RECT 21.33 1.225 21.56 1.245 ;
 RECT 21.33 1.195 21.92 1.225 ;
 RECT 21.47 1.015 21.78 1.035 ;
 RECT 21.33 1.035 21.78 1.055 ;
 RECT 21.605 0.64 21.745 1.015 ;
 RECT 21.78 1.225 21.92 1.75 ;
 RECT 21.485 0.5 21.745 0.64 ;
 RECT 22.38 1.035 22.61 1.055 ;
 RECT 22.38 1.195 22.61 1.245 ;
 RECT 21.33 1.055 22.61 1.195 ;
 RECT 23.35 1.145 23.49 1.345 ;
 RECT 23.03 1.485 23.17 1.76 ;
 RECT 23.35 0.73 23.49 0.935 ;
 RECT 23.03 0.355 23.17 0.59 ;
 RECT 23.03 1.345 23.49 1.485 ;
 RECT 23.305 0.935 23.535 1.145 ;
 RECT 23.03 0.59 23.49 0.73 ;
 RECT 20.29 0.36 20.52 0.43 ;
 RECT 21.885 0.36 22.025 0.565 ;
 RECT 20.29 0.22 22.025 0.36 ;
 RECT 22.625 0.705 22.765 0.75 ;
 RECT 22.75 0.995 23.055 1.205 ;
 RECT 22.75 0.89 22.89 0.995 ;
 RECT 22.625 0.75 22.89 0.89 ;
 RECT 21.885 0.565 22.765 0.705 ;
 RECT 15.525 0.775 15.665 1.405 ;
 RECT 16.25 0.56 16.48 0.635 ;
 RECT 14.505 1.405 15.665 1.545 ;
 RECT 14.505 1.545 14.645 1.83 ;
 RECT 13.46 1.83 14.71 1.97 ;
 RECT 14.505 1.17 14.645 1.405 ;
 RECT 14.435 1.03 14.715 1.17 ;
 RECT 18.445 0.36 18.585 0.635 ;
 RECT 15.525 0.635 18.585 0.775 ;
 RECT 19.125 0.36 19.265 1.25 ;
 RECT 19.125 1.25 19.355 1.46 ;
 RECT 18.445 0.22 19.265 0.36 ;
 RECT 11.48 0.525 11.62 0.885 ;
 RECT 11.48 1.095 11.62 2.065 ;
 RECT 11.48 0.885 11.755 1.095 ;
 RECT 9 2.055 9.14 2.34 ;
 RECT 8.205 2.34 9.14 2.48 ;
 RECT 9.535 1.66 9.675 1.915 ;
 RECT 9 1.915 9.675 2.055 ;
 RECT 8.205 1.04 8.345 2.34 ;
 RECT 8.205 0.895 8.345 0.9 ;
 RECT 8.135 0.9 8.41 1.04 ;
 RECT 9.535 1.52 11.115 1.66 ;
 RECT 10.975 0.525 11.115 1.52 ;
 RECT 10.975 1.66 11.115 2.11 ;
 RECT 10.45 0.765 10.59 1.52 ;
 RECT 10.45 1.66 10.59 2.145 ;
 RECT 12.205 0.585 13.16 0.63 ;
 RECT 12.93 0.63 13.16 0.665 ;
 RECT 12.93 0.455 13.16 0.49 ;
 RECT 12.23 0.49 13.16 0.585 ;
 RECT 12.205 0.63 12.435 0.795 ;
 RECT 13.785 0.57 14.015 0.95 ;
 RECT 16.795 0.22 17.025 0.28 ;
 RECT 16.795 0.42 17.025 0.43 ;
 RECT 14.63 0.28 17.025 0.42 ;
 RECT 14.63 0.42 14.86 0.6 ;
 RECT 3.8 0.66 3.94 0.895 ;
 RECT 3.34 0.52 3.94 0.66 ;
 RECT 4.72 1.035 4.86 1.09 ;
 RECT 5.4 1.035 5.54 1.09 ;
 RECT 7.255 0.885 7.485 0.895 ;
 RECT 7.255 1.035 7.485 1.095 ;
 RECT 3.8 0.895 4.86 1.035 ;
 RECT 5.4 0.895 7.485 1.035 ;
 RECT 4.72 1.09 5.54 1.23 ;
 RECT 3.345 1.82 4.925 1.96 ;
 RECT 4.785 1.79 4.925 1.82 ;
 RECT 3.43 1.96 3.71 2.215 ;
 RECT 3.52 0.805 3.66 1.22 ;
 RECT 3.345 1.22 3.66 1.36 ;
 RECT 3.345 1.36 3.485 1.82 ;
 RECT 5.985 1.615 6.215 1.65 ;
 RECT 5.985 1.79 6.215 1.825 ;
 RECT 4.785 1.65 6.22 1.79 ;
 RECT 2.655 1.67 2.795 1.82 ;
 RECT 2.655 1.96 2.795 2.25 ;
 RECT 2.655 0.715 2.795 1.44 ;
 RECT 2.655 1.44 2.91 1.67 ;
 RECT 2.655 0.505 2.9 0.715 ;
 RECT 2.525 1.82 2.795 1.96 ;
 RECT 0.585 1.335 0.725 2.11 ;
 RECT 0.585 2.25 0.725 2.255 ;
 RECT 0.585 0.875 0.725 1.195 ;
 RECT 0.585 2.11 1.01 2.25 ;
 RECT 0.585 0.735 1.01 0.875 ;
 RECT 0.585 1.195 1.695 1.335 ;
 RECT 1.555 0.6 1.695 1.195 ;
 RECT 3.05 0.36 3.19 2.035 ;
 RECT 2.285 0.36 2.425 0.46 ;
 RECT 3.005 2.17 3.145 2.305 ;
 RECT 3.005 2.035 3.19 2.17 ;
 RECT 2.285 0.22 3.19 0.36 ;
 RECT 1.555 0.46 2.425 0.6 ;
 RECT 12.895 1.895 13.035 2.39 ;
 RECT 17.04 2.205 17.18 2.39 ;
 RECT 12.895 2.39 17.18 2.53 ;
 RECT 11.77 1.755 13.035 1.895 ;
 RECT 11.77 1.895 11.91 2.34 ;
 RECT 10.5 2.3 10.73 2.34 ;
 RECT 10.5 2.48 10.73 2.51 ;
 RECT 10.5 2.34 11.91 2.48 ;
 RECT 20.925 2.205 21.065 2.52 ;
 RECT 17.04 2.065 21.065 2.205 ;
 RECT 25.265 2.48 25.405 2.52 ;
 RECT 20.925 2.52 25.405 2.66 ;
 RECT 25.265 2.27 25.495 2.48 ;
 RECT 16.335 1.7 16.63 1.84 ;
 RECT 16.335 1.84 16.475 2.075 ;
 RECT 15.64 1.84 15.78 2.075 ;
 RECT 15.445 1.7 15.78 1.84 ;
 RECT 15.64 2.075 16.475 2.215 ;
 RECT 16.53 1.055 16.67 1.245 ;
 RECT 15.97 1.385 16.11 1.625 ;
 RECT 16.81 1.385 17.04 1.455 ;
 RECT 15.97 1.245 17.04 1.385 ;
 RECT 16.5 0.915 16.8 1.055 ;
 RECT 15.94 1.625 16.195 1.92 ;
 RECT 13.175 1.56 13.315 2.11 ;
 RECT 12.125 1.405 12.355 1.42 ;
 RECT 12.125 1.56 12.355 1.615 ;
 RECT 12.125 1.42 13.315 1.56 ;
 RECT 13.175 2.11 15.5 2.245 ;
 RECT 13.175 2.245 15.495 2.25 ;
 RECT 15.27 2.035 15.5 2.11 ;
 RECT 8.65 1.775 8.79 2.18 ;
 RECT 8.65 1.04 8.79 1.475 ;
 RECT 8.49 1.475 8.79 1.635 ;
 RECT 8.58 0.9 8.855 1.04 ;
 RECT 8.65 1.685 9.37 1.775 ;
 RECT 8.49 1.635 9.37 1.685 ;
 RECT 9.23 1.21 9.37 1.635 ;
 RECT 3.905 2.105 5.125 2.245 ;
 RECT 5.705 1.225 6.945 1.255 ;
 RECT 6.695 1.205 6.945 1.225 ;
 RECT 6.41 1.365 6.55 2.25 ;
 RECT 5.705 1.365 5.845 1.37 ;
 RECT 3.635 1.5 5.845 1.51 ;
 RECT 4.445 1.37 5.845 1.5 ;
 RECT 3.635 1.51 4.605 1.64 ;
 RECT 3.635 1.64 4.14 1.675 ;
 RECT 5.705 1.255 7.865 1.365 ;
 RECT 6.695 1.365 7.865 1.395 ;
 RECT 7.725 0.885 7.865 0.9 ;
 RECT 7.725 1.04 7.865 1.255 ;
 RECT 7.725 1.395 7.865 2.215 ;
 RECT 7.66 0.9 7.935 1.04 ;
 RECT 1.795 1.63 1.935 1.99 ;
 RECT 1.795 1.475 2.1 1.63 ;
 RECT 1.875 0.905 2.015 1.475 ;
 END
END RDFFSRASRX1

MACRO CGLPPSX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.52 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.52 2.96 ;
 RECT 4.53 1.525 4.76 1.665 ;
 RECT 1.51 2.625 1.74 2.8 ;
 RECT 3.22 2.625 3.45 2.8 ;
 RECT 9.78 1.43 9.92 2.8 ;
 RECT 6.96 1.43 7.1 2.8 ;
 RECT 7.9 1.43 8.04 2.8 ;
 RECT 10.72 1.43 10.86 2.8 ;
 RECT 0.715 1.585 0.855 2.8 ;
 RECT 5.64 2.095 5.78 2.8 ;
 RECT 6.59 1.44 6.73 2.8 ;
 RECT 8.84 1.43 8.98 2.8 ;
 RECT 11.12 1.5 11.26 2.8 ;
 RECT 4.575 1.665 4.715 2.8 ;
 END
 END VDD

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.415 0.84 4.76 1.08 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END SE

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.43 1.12 10.39 1.26 ;
 RECT 10.25 1.47 10.39 2.45 ;
 RECT 7.43 1.26 7.57 2.45 ;
 RECT 7.43 0.475 7.57 1.12 ;
 RECT 9.31 1.26 9.45 2.45 ;
 RECT 9.31 0.475 9.45 1.12 ;
 RECT 8.37 1.26 8.51 2.45 ;
 RECT 8.37 0.475 8.51 1.12 ;
 RECT 10.08 1.26 10.39 1.47 ;
 RECT 10.25 0.475 10.39 1.12 ;
 END
 ANTENNADIFFAREA 2.472 ;
 END GCLK

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.525 1.16 0.92 1.4 ;
 END
 ANTENNAGATEAREA 0.063 ;
 END CLK

 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.575 1.13 1.88 1.43 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.52 0.08 ;
 RECT 1.505 0.585 1.76 0.725 ;
 RECT 4.53 0.515 4.76 0.655 ;
 RECT 3.265 0.08 3.405 0.74 ;
 RECT 5.82 0.08 5.96 0.7 ;
 RECT 9.78 0.08 9.92 0.975 ;
 RECT 6.96 0.08 7.1 0.94 ;
 RECT 0.715 0.08 0.855 0.985 ;
 RECT 8.84 0.08 8.98 0.975 ;
 RECT 1.62 0.08 1.76 0.585 ;
 RECT 10.72 0.08 10.86 0.975 ;
 RECT 7.9 0.08 8.04 0.975 ;
 RECT 11.12 0.08 11.26 0.85 ;
 RECT 4.575 0.08 4.715 0.515 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 2.75 1.56 2.85 2.35 ;
 RECT 2.69 2.35 2.9 2.58 ;
 RECT 3.365 0.89 3.62 1.1 ;
 RECT 4.83 0.285 4.93 2.06 ;
 RECT 3.52 0.34 3.62 0.89 ;
 RECT 3.52 1.1 3.62 2.06 ;
 RECT 3.52 2.06 4.93 2.16 ;
 RECT 4.36 0.865 4.65 1.075 ;
 RECT 4.36 0.285 4.46 0.865 ;
 RECT 4.36 1.075 4.46 1.88 ;
 RECT 1.81 0.37 1.91 1.19 ;
 RECT 1.81 1.4 1.91 2.14 ;
 RECT 1.61 1.19 1.91 1.4 ;
 RECT 0.5 1.17 0.755 1.38 ;
 RECT 0.5 1.38 0.6 2.08 ;
 RECT 0.5 0.57 0.6 1.17 ;
 RECT 0.97 0.19 1.07 2.31 ;
 RECT 0.97 2.31 1.24 2.365 ;
 RECT 0.34 2.365 1.24 2.465 ;
 RECT 0.97 2.465 1.24 2.52 ;
 RECT 2.28 0.19 2.38 0.885 ;
 RECT 0.34 2.31 0.57 2.365 ;
 RECT 0.34 2.465 0.57 2.52 ;
 RECT 0.97 0.09 2.38 0.19 ;
 RECT 6.075 0.09 6.175 1.09 ;
 RECT 5.905 1.19 6.005 2.43 ;
 RECT 4.04 2.34 4.27 2.43 ;
 RECT 4.04 2.53 4.27 2.55 ;
 RECT 4.04 2.43 6.005 2.53 ;
 RECT 5.905 1.09 6.175 1.19 ;
 RECT 5.13 1.2 5.365 1.23 ;
 RECT 5.13 0.29 5.23 1.2 ;
 RECT 5.135 1.33 5.4 1.41 ;
 RECT 5.3 1.41 5.4 2.155 ;
 RECT 5.13 1.23 5.4 1.33 ;
 RECT 3.05 0.315 3.15 1.17 ;
 RECT 3.05 1.38 3.15 2.14 ;
 RECT 2.95 1.17 3.18 1.38 ;
 RECT 2.75 0.315 2.85 0.89 ;
 RECT 2.28 1.26 2.38 2.03 ;
 RECT 2.67 0.89 2.85 0.99 ;
 RECT 2.67 0.99 2.77 1.16 ;
 RECT 2.28 1.16 2.77 1.26 ;
 RECT 2.205 2.03 2.435 2.24 ;
 RECT 6.375 0.09 6.475 2.215 ;
 RECT 6.245 2.215 6.475 2.445 ;
 RECT 7.05 1.25 7.315 1.29 ;
 RECT 7.215 1.29 7.315 2.74 ;
 RECT 7.05 1.08 7.315 1.15 ;
 RECT 7.215 0.225 7.315 1.08 ;
 RECT 8.625 0.225 8.725 1.15 ;
 RECT 8.625 1.25 8.725 2.74 ;
 RECT 9.565 0.225 9.665 1.15 ;
 RECT 9.565 1.25 9.665 2.74 ;
 RECT 9.095 0.225 9.195 1.15 ;
 RECT 9.095 1.25 9.195 2.74 ;
 RECT 10.035 0.225 10.135 1.15 ;
 RECT 10.035 1.25 10.135 2.74 ;
 RECT 8.155 0.225 8.255 1.15 ;
 RECT 8.155 1.25 8.255 2.74 ;
 RECT 10.505 0.225 10.605 1.15 ;
 RECT 10.505 1.25 10.605 2.74 ;
 RECT 7.685 0.225 7.785 1.15 ;
 RECT 7.685 1.25 7.785 2.74 ;
 RECT 7.05 1.15 10.605 1.25 ;
 LAYER CO ;
 RECT 11.125 0.41 11.255 0.54 ;
 RECT 1.56 0.59 1.69 0.72 ;
 RECT 5.825 0.5 5.955 0.63 ;
 RECT 7.905 1.745 8.035 1.875 ;
 RECT 7.435 2.27 7.565 2.4 ;
 RECT 6.595 0.5 6.725 0.63 ;
 RECT 2.03 1.78 2.16 1.91 ;
 RECT 7.435 1.48 7.565 1.61 ;
 RECT 4.11 0.52 4.24 0.65 ;
 RECT 10.725 2.27 10.855 2.4 ;
 RECT 0.25 1.585 0.38 1.715 ;
 RECT 9.315 0.525 9.445 0.655 ;
 RECT 4.58 1.53 4.71 1.66 ;
 RECT 8.375 2.27 8.505 2.4 ;
 RECT 7.435 0.525 7.565 0.655 ;
 RECT 6.965 1.48 7.095 1.61 ;
 RECT 8.845 1.48 8.975 1.61 ;
 RECT 10.725 0.785 10.855 0.915 ;
 RECT 10.255 1.745 10.385 1.875 ;
 RECT 4.11 1.53 4.24 1.66 ;
 RECT 8.845 0.785 8.975 0.915 ;
 RECT 10.255 0.525 10.385 0.655 ;
 RECT 0.25 0.79 0.38 0.92 ;
 RECT 8.375 1.745 8.505 1.875 ;
 RECT 9.785 1.48 9.915 1.61 ;
 RECT 6.295 2.26 6.425 2.39 ;
 RECT 2.5 1.78 2.63 1.91 ;
 RECT 11.125 1.55 11.255 1.68 ;
 RECT 10.255 1.48 10.385 1.61 ;
 RECT 9.785 1.745 9.915 1.875 ;
 RECT 4.58 0.52 4.71 0.65 ;
 RECT 11.125 2.07 11.255 2.2 ;
 RECT 9.315 1.48 9.445 1.61 ;
 RECT 7.1 1.12 7.23 1.25 ;
 RECT 1.19 1.5 1.32 1.63 ;
 RECT 8.845 2.27 8.975 2.4 ;
 RECT 3.74 1.78 3.87 1.91 ;
 RECT 3.415 0.93 3.545 1.06 ;
 RECT 5.645 2.145 5.775 2.275 ;
 RECT 1.56 2.63 1.69 2.76 ;
 RECT 6.965 2.01 7.095 2.14 ;
 RECT 10.725 1.48 10.855 1.61 ;
 RECT 10.725 2.01 10.855 2.14 ;
 RECT 5.35 0.52 5.48 0.65 ;
 RECT 6.965 0.495 7.095 0.625 ;
 RECT 8.375 1.48 8.505 1.61 ;
 RECT 9.315 2.27 9.445 2.4 ;
 RECT 8.845 2.01 8.975 2.14 ;
 RECT 7.905 0.785 8.035 0.915 ;
 RECT 0.575 1.21 0.705 1.34 ;
 RECT 7.905 2.01 8.035 2.14 ;
 RECT 9.315 0.785 9.445 0.915 ;
 RECT 9.315 1.745 9.445 1.875 ;
 RECT 8.375 0.525 8.505 0.655 ;
 RECT 11.125 0.67 11.255 0.8 ;
 RECT 4.47 0.905 4.6 1.035 ;
 RECT 0.72 0.79 0.85 0.92 ;
 RECT 7.905 0.525 8.035 0.655 ;
 RECT 1.66 1.23 1.79 1.36 ;
 RECT 10.255 2.01 10.385 2.14 ;
 RECT 7.905 1.48 8.035 1.61 ;
 RECT 10.725 1.745 10.855 1.875 ;
 RECT 7.435 2.01 7.565 2.14 ;
 RECT 10.725 0.525 10.855 0.655 ;
 RECT 8.375 2.01 8.505 2.14 ;
 RECT 3 1.21 3.13 1.34 ;
 RECT 10.255 0.785 10.385 0.915 ;
 RECT 1.06 2.35 1.19 2.48 ;
 RECT 6.965 1.74 7.095 1.87 ;
 RECT 9.315 2.01 9.445 2.14 ;
 RECT 2.03 0.59 2.16 0.72 ;
 RECT 6.595 1.75 6.725 1.88 ;
 RECT 9.785 2.27 9.915 2.4 ;
 RECT 3.27 0.535 3.4 0.665 ;
 RECT 2.5 0.535 2.63 0.665 ;
 RECT 6.125 1.49 6.255 1.62 ;
 RECT 11.125 1.81 11.255 1.94 ;
 RECT 7.905 2.27 8.035 2.4 ;
 RECT 9.785 0.525 9.915 0.655 ;
 RECT 2.73 2.4 2.86 2.53 ;
 RECT 3.74 0.6 3.87 0.73 ;
 RECT 8.845 1.745 8.975 1.875 ;
 RECT 3.27 2.63 3.4 2.76 ;
 RECT 10.255 2.27 10.385 2.4 ;
 RECT 2.255 2.07 2.385 2.2 ;
 RECT 4.09 2.38 4.22 2.51 ;
 RECT 8.845 0.525 8.975 0.655 ;
 RECT 6.595 1.49 6.725 1.62 ;
 RECT 8.375 0.785 8.505 0.915 ;
 RECT 0.72 1.635 0.85 1.765 ;
 RECT 9.785 0.785 9.915 0.915 ;
 RECT 5.185 1.24 5.315 1.37 ;
 RECT 5.05 1.53 5.18 1.66 ;
 RECT 7.435 0.785 7.565 0.915 ;
 RECT 7.435 1.745 7.565 1.875 ;
 RECT 0.39 2.35 0.52 2.48 ;
 RECT 6.965 0.76 7.095 0.89 ;
 RECT 6.965 2.27 7.095 2.4 ;
 RECT 1.19 0.79 1.32 0.92 ;
 RECT 9.785 2.01 9.915 2.14 ;
 LAYER M1 ;
 RECT 2.025 0.53 2.165 1.775 ;
 RECT 1.98 1.775 2.21 1.915 ;
 RECT 6.12 1.05 6.73 1.115 ;
 RECT 6.59 0.45 6.73 1.05 ;
 RECT 6.12 1.19 6.26 1.67 ;
 RECT 6.12 1.115 7.28 1.19 ;
 RECT 6.58 1.19 7.28 1.255 ;
 RECT 2.495 0.455 2.635 0.925 ;
 RECT 2.495 1.065 2.635 1.775 ;
 RECT 2.45 1.775 2.68 1.915 ;
 RECT 2.495 0.925 3.595 1.065 ;
 RECT 3.735 0.455 3.875 1.205 ;
 RECT 3.735 1.345 3.875 1.775 ;
 RECT 2.95 1.205 3.875 1.345 ;
 RECT 3.69 1.775 3.92 1.915 ;
 RECT 5.51 0.655 5.65 1.525 ;
 RECT 5.3 0.515 5.65 0.655 ;
 RECT 5 1.525 5.97 1.665 ;
 RECT 5.83 1.665 5.97 1.815 ;
 RECT 6.29 1.955 6.43 2.445 ;
 RECT 5.83 1.815 6.43 1.955 ;
 RECT 1.01 2.35 2.865 2.485 ;
 RECT 1.01 2.345 2.86 2.35 ;
 RECT 2.725 2.485 2.865 2.58 ;
 RECT 0.245 0.73 0.385 2.335 ;
 RECT 0.245 2.345 0.57 2.475 ;
 RECT 0.245 2.335 0.535 2.345 ;
 RECT 0.34 2.475 0.57 2.485 ;
 RECT 4.105 0.465 4.245 1.245 ;
 RECT 4.105 1.385 4.245 1.71 ;
 RECT 4.105 1.245 5.365 1.375 ;
 RECT 5.135 1.235 5.365 1.245 ;
 RECT 4.105 1.375 5.315 1.385 ;
 RECT 1.185 0.715 1.325 2.065 ;
 RECT 4.13 2.205 4.27 2.375 ;
 RECT 4.04 2.375 4.27 2.515 ;
 RECT 1.185 2.065 4.27 2.205 ;
 END
END CGLPPSX8

MACRO DELLN1X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 0.99 0.845 1.67 0.985 ;
 RECT 1.525 1.58 1.755 1.79 ;
 RECT 4.65 0.08 4.81 0.755 ;
 RECT 3.205 0.08 3.345 0.85 ;
 RECT 4.155 0.08 4.295 0.85 ;
 RECT 0.99 0.08 1.13 0.845 ;
 RECT 1.53 0.985 1.67 1.58 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 4.155 1.77 4.295 2.8 ;
 RECT 3.205 1.52 3.345 2.8 ;
 RECT 4.665 1.855 4.825 2.8 ;
 RECT 0.99 1.725 1.13 2.8 ;
 RECT 0.99 1.515 1.285 1.725 ;
 END
 END VDD

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.68 1.12 4.525 1.26 ;
 RECT 4.12 1.26 4.525 1.45 ;
 RECT 3.68 1.26 3.82 2.575 ;
 RECT 3.68 0.62 3.82 1.12 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END Z

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.505 1.28 0.825 1.61 ;
 END
 ANTENNAGATEAREA 0.035 ;
 END INP

 OBS
 LAYER PO ;
 RECT 2.99 0.985 3.09 1.51 ;
 RECT 2.23 1.51 3.09 1.61 ;
 RECT 2.99 1.61 3.09 2.745 ;
 RECT 2.23 1.4 2.46 1.51 ;
 RECT 2.89 0.485 3.09 0.985 ;
 RECT 1.245 1.905 1.625 2.005 ;
 RECT 1.525 1.79 1.625 1.905 ;
 RECT 1.245 2.005 1.345 2.79 ;
 RECT 1.525 1.58 1.755 1.79 ;
 RECT 3.935 0.305 4.035 2.745 ;
 RECT 3.46 0.305 3.56 2.745 ;
 RECT 2.38 0.205 4.035 0.305 ;
 RECT 2.38 0.305 2.61 0.43 ;
 RECT 1.745 0.28 1.845 0.465 ;
 RECT 1.945 1.04 2.045 2.2 ;
 RECT 1.545 2.3 1.645 2.775 ;
 RECT 0.365 0.28 0.595 0.455 ;
 RECT 1.645 0.465 1.845 0.94 ;
 RECT 1.545 2.2 2.045 2.3 ;
 RECT 0.365 0.18 1.845 0.28 ;
 RECT 1.645 0.94 2.045 1.04 ;
 RECT 1.245 0.965 1.345 1.515 ;
 RECT 1.055 1.515 1.345 1.725 ;
 RECT 1.245 0.465 1.445 0.965 ;
 RECT 0.775 0.46 0.875 1.39 ;
 RECT 0.595 1.39 0.875 1.6 ;
 RECT 0.775 1.6 0.875 2.78 ;
 LAYER CO ;
 RECT 3.685 1.845 3.815 1.975 ;
 RECT 3.685 1.57 3.815 1.7 ;
 RECT 4.16 2.395 4.29 2.525 ;
 RECT 4.16 2.12 4.29 2.25 ;
 RECT 4.16 1.845 4.29 1.975 ;
 RECT 3.685 2.395 3.815 2.525 ;
 RECT 3.21 1.855 3.34 1.985 ;
 RECT 3.21 2.125 3.34 2.255 ;
 RECT 3.21 2.395 3.34 2.525 ;
 RECT 4.665 0.305 4.795 0.435 ;
 RECT 4.665 0.575 4.795 0.705 ;
 RECT 4.68 1.905 4.81 2.035 ;
 RECT 4.68 2.175 4.81 2.305 ;
 RECT 3.21 1.57 3.34 1.7 ;
 RECT 2.64 0.67 2.77 0.8 ;
 RECT 3.685 2.12 3.815 2.25 ;
 RECT 2.43 0.26 2.56 0.39 ;
 RECT 2.28 1.44 2.41 1.57 ;
 RECT 1.575 1.62 1.705 1.75 ;
 RECT 1.105 1.555 1.235 1.685 ;
 RECT 0.525 2.43 0.655 2.56 ;
 RECT 1.775 2.43 1.905 2.56 ;
 RECT 0.415 0.285 0.545 0.415 ;
 RECT 3.685 1.57 3.815 1.7 ;
 RECT 3.685 1.845 3.815 1.975 ;
 RECT 3.685 2.12 3.815 2.25 ;
 RECT 4.16 1.845 4.29 1.975 ;
 RECT 4.16 2.12 4.29 2.25 ;
 RECT 4.16 2.395 4.29 2.525 ;
 RECT 3.685 2.395 3.815 2.525 ;
 RECT 4.16 0.67 4.29 0.8 ;
 RECT 3.685 0.67 3.815 0.8 ;
 RECT 2.74 2.395 2.87 2.525 ;
 RECT 3.21 0.67 3.34 0.8 ;
 RECT 1.965 0.65 2.095 0.78 ;
 RECT 0.525 0.65 0.655 0.78 ;
 RECT 0.995 0.65 1.125 0.78 ;
 RECT 0.995 2.43 1.125 2.56 ;
 RECT 4.68 2.175 4.81 2.305 ;
 RECT 4.665 0.305 4.795 0.435 ;
 RECT 4.665 0.575 4.795 0.705 ;
 RECT 0.645 1.43 0.775 1.56 ;
 LAYER M1 ;
 RECT 0.22 0.905 0.36 2.04 ;
 RECT 0.365 0.245 0.66 0.455 ;
 RECT 0.52 0.455 0.66 0.765 ;
 RECT 0.52 2.18 0.66 2.61 ;
 RECT 0.22 2.04 0.66 2.18 ;
 RECT 0.22 0.765 0.66 0.905 ;
 RECT 2.49 0.43 2.63 0.665 ;
 RECT 2.735 0.805 2.875 2.575 ;
 RECT 2.38 0.22 2.63 0.43 ;
 RECT 2.49 0.665 2.875 0.805 ;
 RECT 2.12 0.785 2.26 1.4 ;
 RECT 2.12 1.4 2.46 1.61 ;
 RECT 2.12 1.61 2.26 2.425 ;
 RECT 1.915 0.645 2.26 0.785 ;
 RECT 1.715 2.425 2.26 2.565 ;
 END
END DELLN1X2

MACRO DELLN2X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 0.99 0.845 1.67 0.985 ;
 RECT 1.525 1.58 1.755 1.79 ;
 RECT 4.36 0.08 4.5 0.85 ;
 RECT 4.855 0.08 5.015 0.755 ;
 RECT 3.41 0.08 3.55 0.85 ;
 RECT 0.99 0.08 1.13 0.845 ;
 RECT 1.53 0.985 1.67 1.58 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 4.36 1.735 4.5 2.8 ;
 RECT 4.87 1.855 5.03 2.8 ;
 RECT 3.41 1.52 3.55 2.8 ;
 RECT 0.99 1.725 1.13 2.8 ;
 RECT 0.99 1.515 1.285 1.725 ;
 END
 END VDD

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.885 1.12 4.535 1.26 ;
 RECT 4.165 1.26 4.535 1.475 ;
 RECT 4.165 1.065 4.535 1.12 ;
 RECT 3.885 1.26 4.025 2.575 ;
 RECT 3.885 0.62 4.025 1.12 ;
 END
 ANTENNADIFFAREA 0.578 ;
 END Z

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.45 1.125 0.825 1.515 ;
 END
 ANTENNAGATEAREA 0.028 ;
 END INP

 OBS
 LAYER PO ;
 RECT 1.245 1.905 1.625 2.005 ;
 RECT 1.525 1.79 1.625 1.905 ;
 RECT 1.245 2.005 1.375 2.745 ;
 RECT 1.525 1.58 1.755 1.79 ;
 RECT 2.3 1.4 2.53 1.51 ;
 RECT 2.3 1.51 3.295 1.61 ;
 RECT 3.155 0.985 3.295 1.51 ;
 RECT 3.155 1.61 3.295 2.745 ;
 RECT 2.925 0.485 3.295 0.985 ;
 RECT 3.665 0.275 3.765 2.745 ;
 RECT 4.14 0.275 4.24 2.745 ;
 RECT 2.51 0.275 2.74 0.435 ;
 RECT 2.51 0.175 4.245 0.275 ;
 RECT 0.365 0.18 1.915 0.28 ;
 RECT 1.815 0.28 1.915 0.465 ;
 RECT 0.365 0.28 0.595 0.455 ;
 RECT 1.945 0.965 2.045 2.195 ;
 RECT 1.575 2.295 1.705 2.745 ;
 RECT 1.815 0.465 2.185 0.965 ;
 RECT 1.575 2.195 2.045 2.295 ;
 RECT 1.245 0.965 1.345 1.515 ;
 RECT 1.055 1.515 1.345 1.725 ;
 RECT 1.245 0.465 1.615 0.965 ;
 RECT 0.775 0.46 0.875 1.215 ;
 RECT 0.595 1.215 0.875 1.425 ;
 RECT 0.775 1.425 0.875 2.745 ;
 LAYER CO ;
 RECT 3.415 0.67 3.545 0.8 ;
 RECT 2.675 0.67 2.805 0.8 ;
 RECT 2.305 0.65 2.435 0.78 ;
 RECT 0.525 0.65 0.655 0.78 ;
 RECT 0.995 0.65 1.125 0.78 ;
 RECT 3.89 2.12 4.02 2.25 ;
 RECT 3.89 1.845 4.02 1.975 ;
 RECT 3.89 1.57 4.02 1.7 ;
 RECT 3.89 2.395 4.02 2.525 ;
 RECT 0.415 0.285 0.545 0.415 ;
 RECT 3.89 1.845 4.02 1.975 ;
 RECT 3.89 2.12 4.02 2.25 ;
 RECT 4.365 1.845 4.495 1.975 ;
 RECT 4.365 2.12 4.495 2.25 ;
 RECT 2.56 0.265 2.69 0.395 ;
 RECT 2.35 1.44 2.48 1.57 ;
 RECT 4.885 2.175 5.015 2.305 ;
 RECT 4.87 0.305 5 0.435 ;
 RECT 4.87 0.575 5 0.705 ;
 RECT 3.415 1.855 3.545 1.985 ;
 RECT 3.415 2.125 3.545 2.255 ;
 RECT 3.415 2.395 3.545 2.525 ;
 RECT 4.87 0.305 5 0.435 ;
 RECT 4.87 0.575 5 0.705 ;
 RECT 4.885 1.905 5.015 2.035 ;
 RECT 4.885 2.175 5.015 2.305 ;
 RECT 3.415 1.57 3.545 1.7 ;
 RECT 3.89 1.57 4.02 1.7 ;
 RECT 4.365 2.395 4.495 2.525 ;
 RECT 4.365 2.12 4.495 2.25 ;
 RECT 4.365 1.845 4.495 1.975 ;
 RECT 1.575 1.62 1.705 1.75 ;
 RECT 1.105 1.555 1.235 1.685 ;
 RECT 0.525 2.43 0.655 2.56 ;
 RECT 1.825 2.43 1.955 2.56 ;
 RECT 4.365 2.395 4.495 2.525 ;
 RECT 3.89 2.395 4.02 2.525 ;
 RECT 4.365 0.67 4.495 0.8 ;
 RECT 3.89 0.67 4.02 0.8 ;
 RECT 2.905 2.395 3.035 2.525 ;
 RECT 0.995 2.43 1.125 2.56 ;
 RECT 0.645 1.255 0.775 1.385 ;
 LAYER M1 ;
 RECT 0.12 0.905 0.26 1.935 ;
 RECT 0.365 0.245 0.66 0.455 ;
 RECT 0.52 0.455 0.66 0.765 ;
 RECT 0.12 0.765 0.66 0.905 ;
 RECT 0.12 1.935 0.66 2.075 ;
 RECT 0.52 2.075 0.66 2.61 ;
 RECT 2.3 0.6 2.44 1.4 ;
 RECT 2.3 1.61 2.44 2.425 ;
 RECT 1.765 2.425 2.44 2.565 ;
 RECT 2.3 1.4 2.53 1.61 ;
 RECT 2.51 0.225 2.81 0.435 ;
 RECT 2.67 0.435 2.81 2.39 ;
 RECT 2.67 2.39 3.09 2.53 ;
 END
END DELLN2X2

MACRO DELLN3X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.68 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.68 0.08 ;
 RECT 0.99 0.845 1.67 0.985 ;
 RECT 3.385 0.845 4.065 0.985 ;
 RECT 1.525 1.845 1.755 2.055 ;
 RECT 3.92 1.845 4.15 2.055 ;
 RECT 7.23 0.08 7.39 0.755 ;
 RECT 6.735 0.08 6.875 0.85 ;
 RECT 5.785 0.08 5.925 0.85 ;
 RECT 0.99 0.08 1.13 0.845 ;
 RECT 3.385 0.08 3.525 0.845 ;
 RECT 1.53 0.985 1.67 1.845 ;
 RECT 3.925 0.985 4.065 1.845 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.68 2.96 ;
 RECT 6.735 1.785 6.875 2.8 ;
 RECT 5.785 1.52 5.925 2.8 ;
 RECT 7.235 1.855 7.395 2.8 ;
 RECT 3.385 1.385 3.525 2.8 ;
 RECT 3.385 1.175 3.705 1.385 ;
 RECT 0.99 1.765 1.13 2.8 ;
 RECT 0.99 1.555 1.305 1.765 ;
 END
 END VDD

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.26 1.5 6.4 2.575 ;
 RECT 6.26 1.12 7.06 1.5 ;
 RECT 6.26 0.62 6.4 1.12 ;
 END
 ANTENNADIFFAREA 0.578 ;
 END Z

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.485 1.155 0.845 1.365 ;
 RECT 0.485 1.365 0.84 1.485 ;
 RECT 0.485 1.04 0.84 1.155 ;
 END
 ANTENNAGATEAREA 0.028 ;
 END INP

 OBS
 LAYER PO ;
 RECT 3.64 1.955 4.15 2.055 ;
 RECT 3.64 2.055 3.76 2.775 ;
 RECT 3.92 1.845 4.15 1.955 ;
 RECT 3.475 1.175 3.74 1.385 ;
 RECT 3.64 0.965 3.74 1.175 ;
 RECT 3.64 0.465 4 0.965 ;
 RECT 2.5 0.18 4.3 0.28 ;
 RECT 4.2 0.28 4.3 0.465 ;
 RECT 2.5 0.28 2.73 0.43 ;
 RECT 4.46 0.965 4.56 2.24 ;
 RECT 3.96 2.34 4.08 2.775 ;
 RECT 4.2 0.465 4.56 0.965 ;
 RECT 3.96 2.24 4.56 2.34 ;
 RECT 1.245 1.955 1.755 2.055 ;
 RECT 1.525 1.845 1.755 1.955 ;
 RECT 1.245 2.055 1.365 2.775 ;
 RECT 6.04 0.225 6.14 2.745 ;
 RECT 6.515 0.225 6.615 2.745 ;
 RECT 4.89 0.225 5.12 0.43 ;
 RECT 4.89 0.125 6.615 0.225 ;
 RECT 5.56 0.985 5.67 1.51 ;
 RECT 5.56 1.61 5.67 2.71 ;
 RECT 4.745 1.51 5.67 1.61 ;
 RECT 4.745 1.45 4.975 1.51 ;
 RECT 4.745 1.61 4.975 1.66 ;
 RECT 5.38 0.485 5.67 0.985 ;
 RECT 3.15 0.965 3.27 1.56 ;
 RECT 2.345 1.56 3.27 1.66 ;
 RECT 3.15 1.66 3.27 2.775 ;
 RECT 2.345 1.45 2.575 1.56 ;
 RECT 2.91 0.465 3.27 0.965 ;
 RECT 1.245 0.965 1.345 1.555 ;
 RECT 1.075 1.555 1.345 1.765 ;
 RECT 1.245 0.465 1.605 0.965 ;
 RECT 1.565 2.24 2.165 2.335 ;
 RECT 2.065 0.965 2.165 2.24 ;
 RECT 1.565 2.335 2.1 2.34 ;
 RECT 1.565 2.34 1.685 2.775 ;
 RECT 1.805 0.28 1.905 0.465 ;
 RECT 0.365 0.18 1.905 0.28 ;
 RECT 0.365 0.28 0.595 0.43 ;
 RECT 1.805 0.465 2.165 0.965 ;
 RECT 0.775 0.46 0.875 1.155 ;
 RECT 0.615 1.155 0.875 1.365 ;
 RECT 0.775 1.365 0.875 2.77 ;
 LAYER CO ;
 RECT 3.97 1.885 4.1 2.015 ;
 RECT 4.795 1.49 4.925 1.62 ;
 RECT 4.94 0.26 5.07 0.39 ;
 RECT 3.525 1.215 3.655 1.345 ;
 RECT 2.395 1.49 2.525 1.62 ;
 RECT 1.125 1.595 1.255 1.725 ;
 RECT 0.415 0.26 0.545 0.39 ;
 RECT 7.25 2.175 7.38 2.305 ;
 RECT 6.265 2.12 6.395 2.25 ;
 RECT 6.265 1.845 6.395 1.975 ;
 RECT 6.265 1.57 6.395 1.7 ;
 RECT 6.74 2.395 6.87 2.525 ;
 RECT 6.74 2.12 6.87 2.25 ;
 RECT 6.74 1.845 6.87 1.975 ;
 RECT 6.265 2.395 6.395 2.525 ;
 RECT 4.68 0.65 4.81 0.78 ;
 RECT 3.39 2.455 3.52 2.585 ;
 RECT 2.66 0.65 2.79 0.78 ;
 RECT 2.9 2.455 3.03 2.585 ;
 RECT 3.39 0.65 3.52 0.78 ;
 RECT 4.2 2.455 4.33 2.585 ;
 RECT 5.79 1.855 5.92 1.985 ;
 RECT 5.79 2.125 5.92 2.255 ;
 RECT 5.79 2.395 5.92 2.525 ;
 RECT 7.245 0.305 7.375 0.435 ;
 RECT 7.245 0.575 7.375 0.705 ;
 RECT 7.25 1.905 7.38 2.035 ;
 RECT 7.25 2.175 7.38 2.305 ;
 RECT 5.79 1.57 5.92 1.7 ;
 RECT 6.265 1.57 6.395 1.7 ;
 RECT 6.265 1.845 6.395 1.975 ;
 RECT 6.265 2.12 6.395 2.25 ;
 RECT 6.74 1.845 6.87 1.975 ;
 RECT 6.74 2.12 6.87 2.25 ;
 RECT 6.74 2.395 6.87 2.525 ;
 RECT 6.265 2.395 6.395 2.525 ;
 RECT 6.74 0.67 6.87 0.8 ;
 RECT 6.265 0.67 6.395 0.8 ;
 RECT 5.3 2.395 5.43 2.525 ;
 RECT 5.79 0.67 5.92 0.8 ;
 RECT 5.08 0.67 5.21 0.8 ;
 RECT 2.285 0.65 2.415 0.78 ;
 RECT 0.525 0.65 0.655 0.78 ;
 RECT 0.995 0.65 1.125 0.78 ;
 RECT 1.805 2.455 1.935 2.585 ;
 RECT 0.995 2.455 1.125 2.585 ;
 RECT 0.525 2.455 0.655 2.585 ;
 RECT 2.55 0.26 2.68 0.39 ;
 RECT 1.575 1.885 1.705 2.015 ;
 RECT 7.245 0.305 7.375 0.435 ;
 RECT 7.245 0.575 7.375 0.705 ;
 RECT 0.665 1.195 0.795 1.325 ;
 LAYER M1 ;
 RECT 2.65 0.43 2.79 0.645 ;
 RECT 2.5 0.28 2.79 0.43 ;
 RECT 2.5 0.22 2.73 0.28 ;
 RECT 2.895 0.785 3.035 2.635 ;
 RECT 2.61 0.645 3.035 0.785 ;
 RECT 4.675 1.66 4.815 2.45 ;
 RECT 4.675 0.6 4.815 1.45 ;
 RECT 4.675 1.45 4.975 1.66 ;
 RECT 4.15 2.45 4.815 2.59 ;
 RECT 0.16 0.895 0.3 1.84 ;
 RECT 0.52 0.43 0.66 0.755 ;
 RECT 0.52 0.895 0.66 0.9 ;
 RECT 0.16 1.84 0.66 1.98 ;
 RECT 0.52 1.98 0.66 2.635 ;
 RECT 0.16 0.755 0.66 0.895 ;
 RECT 0.365 0.22 0.66 0.43 ;
 RECT 4.89 0.22 5.16 0.43 ;
 RECT 5.02 0.43 5.16 0.665 ;
 RECT 5.02 0.665 5.435 0.805 ;
 RECT 5.295 0.805 5.435 2.575 ;
 RECT 2.28 0.6 2.42 1.45 ;
 RECT 2.28 1.45 2.575 1.66 ;
 RECT 2.28 1.66 2.42 2.45 ;
 RECT 1.74 2.45 2.42 2.59 ;
 END
END DELLN3X2

MACRO RDFFSRASRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 29.76 BY 2.88 ;
 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.325 1.475 1.655 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.75 2.12 10.08 2.47 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.92 0.59 23.29 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.86 0.08 2.14 0.295 ;
 RECT 26.59 0.08 26.83 0.26 ;
 RECT 5.79 0.31 6.08 0.45 ;
 RECT 9.475 0.615 9.745 0.755 ;
 RECT 13.4 0.275 14.425 0.415 ;
 RECT 18.985 0.335 19.25 0.495 ;
 RECT 17.98 0.335 18.245 0.495 ;
 RECT 14.285 0.75 15.23 0.89 ;
 RECT 0 -0.08 29.76 0.08 ;
 RECT 1.275 0.08 1.415 0.97 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.685 0.08 4.92 0.46 ;
 RECT 20.5 0.08 20.64 0.82 ;
 RECT 21.565 0.08 21.705 0.82 ;
 RECT 24.24 0.08 24.38 0.36 ;
 RECT 25.455 0.08 25.595 0.35 ;
 RECT 5.87 0.08 6.01 0.31 ;
 RECT 9.54 0.08 9.68 0.615 ;
 RECT 13.4 0.415 13.54 0.945 ;
 RECT 13.4 0.08 13.54 0.275 ;
 RECT 19.04 0.08 19.18 0.335 ;
 RECT 18.035 0.08 18.175 0.335 ;
 RECT 15.09 0.89 15.23 1.11 ;
 RECT 14.285 0.415 14.425 0.75 ;
 END
 END VSS

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.24 1.795 7.48 2.04 ;
 RECT 6.69 1.795 6.92 1.83 ;
 RECT 6.69 1.655 7.48 1.795 ;
 RECT 6.69 1.62 6.92 1.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 28.11 1.435 28.47 1.8 ;
 RECT 26.47 1.99 28.335 2.13 ;
 RECT 24.24 2.22 26.61 2.36 ;
 RECT 26.47 1.435 26.61 1.99 ;
 RECT 28.195 1.8 28.335 1.99 ;
 RECT 24.24 1.39 24.38 2.22 ;
 RECT 25.625 1.37 25.765 2.22 ;
 RECT 26.47 2.13 26.61 2.22 ;
 END
 END VDDG

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 9.285 2.215 9.56 2.355 ;
 RECT 0 2.8 29.76 2.96 ;
 RECT 2.015 2.34 2.265 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.275 1.98 1.415 2.8 ;
 RECT 6.9 2 7.04 2.8 ;
 RECT 5.87 1.98 6.01 2.8 ;
 RECT 5.39 2.07 5.53 2.8 ;
 RECT 9.35 2.195 9.49 2.215 ;
 RECT 12.31 2.335 12.58 2.8 ;
 RECT 20.415 2.57 20.555 2.8 ;
 RECT 17.95 2.57 18.09 2.8 ;
 RECT 18.955 2.57 19.095 2.8 ;
 RECT 21.48 2.57 21.62 2.8 ;
 RECT 9.35 2.355 9.49 2.8 ;
 END
 END VDD

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.08 0.485 4.395 0.605 ;
 RECT 9 0.895 10.055 1.035 ;
 RECT 9.91 0.245 12.06 0.255 ;
 RECT 9.91 0.255 12.065 0.385 ;
 RECT 11.925 1.09 13.915 1.23 ;
 RECT 14.12 1.56 14.35 1.6 ;
 RECT 13.775 1.42 14.35 1.56 ;
 RECT 14.12 1.39 14.35 1.42 ;
 RECT 4.08 0.605 9.14 0.745 ;
 RECT 9 0.745 9.14 0.895 ;
 RECT 9.915 0.385 10.055 0.895 ;
 RECT 11.925 0.385 12.065 1.09 ;
 RECT 13.775 1.23 13.915 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.77 0.22 1.135 0.525 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.34 1.205 17.685 1.445 ;
 RECT 17.545 0.915 17.685 1.205 ;
 RECT 17.545 1.84 17.685 1.885 ;
 RECT 17.545 1.445 17.685 1.7 ;
 RECT 18.55 1.84 18.69 1.885 ;
 RECT 18.55 0.915 18.69 1.7 ;
 RECT 19.525 1.84 19.665 1.885 ;
 RECT 19.525 0.915 19.665 1.7 ;
 RECT 17.545 1.7 19.665 1.84 ;
 END
 ANTENNADIFFAREA 1.145 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.82 1.095 20.08 1.335 ;
 RECT 19.94 0.51 20.08 1.095 ;
 RECT 21 1.905 21.14 1.91 ;
 RECT 21 0.56 21.14 1.765 ;
 RECT 22.065 1.905 22.205 1.91 ;
 RECT 22.065 0.56 22.205 1.765 ;
 RECT 19.94 1.905 20.08 1.915 ;
 RECT 19.94 1.335 20.08 1.765 ;
 RECT 19.94 1.765 22.205 1.905 ;
 END
 ANTENNADIFFAREA 0.937 ;
 END Q

 OBS
 LAYER PO ;
 RECT 11.525 1.025 11.755 1.095 ;
 RECT 12.205 0.795 12.37 0.925 ;
 RECT 12.205 0.585 12.435 0.795 ;
 RECT 25.715 0.38 25.815 0.96 ;
 RECT 25.715 1.06 25.815 1.14 ;
 RECT 25.295 0.935 25.525 0.96 ;
 RECT 25.295 0.96 25.815 1.06 ;
 RECT 25.295 1.06 25.525 1.145 ;
 RECT 25.715 1.14 25.985 1.24 ;
 RECT 25.885 1.24 25.985 1.84 ;
 RECT 26.08 0.22 26.31 0.28 ;
 RECT 26.08 0.38 26.31 0.43 ;
 RECT 25.715 0.28 26.31 0.38 ;
 RECT 24.025 0.21 24.125 0.755 ;
 RECT 24.025 0.855 24.125 2.2 ;
 RECT 26.89 1.125 26.99 2.2 ;
 RECT 23.06 0.755 24.595 0.84 ;
 RECT 23.06 0.84 24.59 0.855 ;
 RECT 24.495 0.215 24.595 0.755 ;
 RECT 23.06 0.595 23.29 0.755 ;
 RECT 24.025 2.2 26.99 2.3 ;
 RECT 10.195 0.655 10.295 2.305 ;
 RECT 10.5 2.3 10.73 2.305 ;
 RECT 10.5 2.405 10.73 2.51 ;
 RECT 10.195 2.305 10.73 2.405 ;
 RECT 20.185 1.33 21.945 1.43 ;
 RECT 21.845 0.375 21.945 1.33 ;
 RECT 20.185 1.2 20.395 1.33 ;
 RECT 20.185 1.43 20.395 1.435 ;
 RECT 20.2 0.385 20.3 1.2 ;
 RECT 20.2 1.435 20.3 2.455 ;
 RECT 20.78 0.385 20.88 1.33 ;
 RECT 20.78 1.43 20.88 2.46 ;
 RECT 21.265 0.385 21.365 1.33 ;
 RECT 21.265 1.43 21.365 2.455 ;
 RECT 21.845 1.43 21.945 2.465 ;
 RECT 22.475 0.22 22.705 0.275 ;
 RECT 22.475 0.375 22.705 0.43 ;
 RECT 21.845 0.275 22.705 0.375 ;
 RECT 14.255 0.73 14.355 1.39 ;
 RECT 14.12 1.39 14.355 1.6 ;
 RECT 14.255 1.6 14.355 2.39 ;
 RECT 12.93 0.455 14.86 0.535 ;
 RECT 14.63 0.535 14.86 0.6 ;
 RECT 13.785 0.535 14.015 0.835 ;
 RECT 13.785 0.835 13.885 2.39 ;
 RECT 14.63 0.39 14.86 0.435 ;
 RECT 13.01 0.435 14.86 0.455 ;
 RECT 12.93 0.535 13.16 0.665 ;
 RECT 15.285 1.445 15.385 2.035 ;
 RECT 15.27 2.035 15.5 2.245 ;
 RECT 17.81 0.39 17.91 1.4 ;
 RECT 17.81 1.5 17.91 2.37 ;
 RECT 16.86 0.43 16.96 1.245 ;
 RECT 16.795 0.29 17.91 0.39 ;
 RECT 19.305 0.51 19.405 1.4 ;
 RECT 19.305 1.5 19.405 2.37 ;
 RECT 18.815 0.515 18.915 1.4 ;
 RECT 18.815 1.5 18.915 2.37 ;
 RECT 17.81 1.4 19.405 1.5 ;
 RECT 18.3 0.51 18.4 1.4 ;
 RECT 18.3 1.5 18.4 2.37 ;
 RECT 16.795 0.22 17.025 0.29 ;
 RECT 16.795 0.39 17.025 0.43 ;
 RECT 16.81 1.245 17.04 1.455 ;
 RECT 16.225 0.77 16.325 2.155 ;
 RECT 16.225 0.55 16.325 0.56 ;
 RECT 16.225 0.56 16.48 0.77 ;
 RECT 27.2 0.375 27.3 0.99 ;
 RECT 27.2 0.99 27.45 1.2 ;
 RECT 27.2 1.2 27.3 2.27 ;
 RECT 27.2 2.27 27.485 2.48 ;
 RECT 24.805 0.215 24.905 0.995 ;
 RECT 24.805 0.995 25.045 1.205 ;
 RECT 24.805 1.205 24.905 2 ;
 RECT 15.755 0.55 15.855 2.69 ;
 RECT 6.685 1.58 6.785 1.62 ;
 RECT 6.425 1.01 6.525 1.48 ;
 RECT 6.685 1.83 6.785 2.69 ;
 RECT 6.685 1.62 6.92 1.83 ;
 RECT 6.425 1.48 6.785 1.58 ;
 RECT 6.685 2.69 15.855 2.79 ;
 RECT 11.23 0.195 11.33 1.29 ;
 RECT 12.125 1.39 12.32 1.405 ;
 RECT 2.785 0.285 2.885 0.505 ;
 RECT 4.495 0.285 4.595 1.24 ;
 RECT 2.785 0.185 11.33 0.195 ;
 RECT 2.785 0.195 4.595 0.285 ;
 RECT 4.495 0.095 11.33 0.185 ;
 RECT 11.23 1.29 12.32 1.39 ;
 RECT 2.67 0.505 2.9 0.715 ;
 RECT 12.125 1.405 12.355 1.615 ;
 RECT 3.755 1.33 3.895 1.475 ;
 RECT 3.755 1.71 3.855 2.475 ;
 RECT 3.795 0.65 3.895 1.33 ;
 RECT 3.755 1.475 3.985 1.71 ;
 RECT 9.8 0.655 9.9 1.24 ;
 RECT 9.205 1.155 9.435 1.24 ;
 RECT 9.205 1.34 9.435 1.39 ;
 RECT 9.205 1.24 9.9 1.34 ;
 RECT 1.535 0.49 1.635 1.495 ;
 RECT 1.34 1.495 1.635 1.745 ;
 RECT 1.535 1.745 1.635 2.37 ;
 RECT 1.06 0.52 1.16 2.465 ;
 RECT 0.82 0.27 1.16 0.52 ;
 RECT 3.26 1.665 3.36 2.49 ;
 RECT 2.72 1.445 2.965 1.565 ;
 RECT 2.72 1.565 3.36 1.665 ;
 RECT 2.72 1.665 2.965 1.69 ;
 RECT 2.375 1.62 2.475 2.675 ;
 RECT 3.305 0.47 3.59 0.705 ;
 RECT 3.305 0.705 3.405 1.155 ;
 RECT 2.39 0.715 2.49 1.155 ;
 RECT 2.39 1.155 3.405 1.255 ;
 RECT 2.39 1.255 2.49 1.52 ;
 RECT 2.375 2.675 5.275 2.775 ;
 RECT 5.175 1.79 5.275 2.675 ;
 RECT 1.815 1.44 2.06 1.52 ;
 RECT 1.815 1.62 2.06 1.69 ;
 RECT 1.815 1.52 2.49 1.62 ;
 RECT 4.195 0.715 4.295 1.61 ;
 RECT 4.23 1.71 4.33 2.48 ;
 RECT 4.195 1.61 4.33 1.71 ;
 RECT 4.075 0.485 4.315 0.715 ;
 RECT 8.905 0.655 9.005 1.18 ;
 RECT 8.905 1.28 9.005 1.655 ;
 RECT 7.99 0.66 8.09 1.18 ;
 RECT 8.905 1.655 9.865 1.755 ;
 RECT 9.765 1.755 9.865 2.255 ;
 RECT 8.905 1.755 9.005 2.51 ;
 RECT 7.99 1.18 9.005 1.28 ;
 RECT 9.765 2.255 9.995 2.465 ;
 RECT 27.9 0.195 28 2.665 ;
 RECT 26.89 0.095 28 0.195 ;
 RECT 23.265 1.245 23.365 2.665 ;
 RECT 26.89 0.195 26.99 0.945 ;
 RECT 23.265 1.2 23.55 1.245 ;
 RECT 23.32 1.035 23.55 1.1 ;
 RECT 23.265 2.665 28 2.765 ;
 RECT 23.265 1.1 23.595 1.2 ;
 RECT 6.125 0.98 6.225 1.615 ;
 RECT 5.985 1.615 6.225 1.825 ;
 RECT 6.125 1.825 6.225 2.51 ;
 RECT 12.62 0.105 15.445 0.205 ;
 RECT 12.62 0.205 12.72 1.91 ;
 RECT 15.345 0.205 15.445 1.265 ;
 RECT 11.8 1.71 11.9 1.91 ;
 RECT 10.715 1.61 11.9 1.71 ;
 RECT 10.715 0.475 10.815 1.61 ;
 RECT 11.265 1.71 11.365 2.425 ;
 RECT 7.38 0.475 7.48 0.895 ;
 RECT 11.8 1.91 12.72 2.01 ;
 RECT 7.38 0.375 10.815 0.475 ;
 RECT 7.255 0.895 7.485 1.105 ;
 RECT 7.98 1.575 8.08 2.485 ;
 RECT 8.49 1.575 8.72 1.685 ;
 RECT 7.98 1.475 8.72 1.575 ;
 RECT 24.5 1.245 24.6 2.02 ;
 RECT 24.37 1.035 24.6 1.245 ;
 RECT 11.525 0.885 11.755 0.925 ;
 RECT 11.525 0.925 12.37 1.025 ;
 LAYER CO ;
 RECT 3.505 2.07 3.635 2.2 ;
 RECT 18.555 0.975 18.685 1.105 ;
 RECT 2.085 2.345 2.215 2.475 ;
 RECT 10.455 1.945 10.585 2.075 ;
 RECT 28.2 1.475 28.33 1.605 ;
 RECT 0.81 0.74 0.94 0.87 ;
 RECT 20.42 2.64 20.55 2.77 ;
 RECT 6.685 1.23 6.815 1.36 ;
 RECT 1.95 0.145 2.08 0.275 ;
 RECT 21.57 0.62 21.7 0.75 ;
 RECT 19.045 0.36 19.175 0.49 ;
 RECT 8.655 0.905 8.785 1.035 ;
 RECT 10.455 0.875 10.585 1.005 ;
 RECT 26.64 0.12 26.77 0.25 ;
 RECT 3.41 0.525 3.54 0.655 ;
 RECT 17.55 1.705 17.68 1.835 ;
 RECT 8.655 1.995 8.785 2.125 ;
 RECT 20.225 1.25 20.355 1.38 ;
 RECT 5.875 2.075 6.005 2.205 ;
 RECT 10.98 0.595 11.11 0.725 ;
 RECT 2.595 1.825 2.725 1.955 ;
 RECT 21.485 2.64 21.615 2.77 ;
 RECT 19.945 1.725 20.075 1.855 ;
 RECT 13.405 0.765 13.535 0.895 ;
 RECT 18.04 0.36 18.17 0.49 ;
 RECT 15.975 1.705 16.105 1.835 ;
 RECT 19.945 0.62 20.075 0.75 ;
 RECT 19.53 0.975 19.66 1.105 ;
 RECT 24.245 1.475 24.375 1.605 ;
 RECT 6.905 2.11 7.035 2.24 ;
 RECT 21.005 0.63 21.135 0.76 ;
 RECT 9.815 2.295 9.945 2.425 ;
 RECT 25.345 0.975 25.475 1.105 ;
 RECT 13.835 0.665 13.965 0.795 ;
 RECT 16.86 1.285 16.99 1.415 ;
 RECT 14.68 0.43 14.81 0.56 ;
 RECT 23.37 1.075 23.5 1.205 ;
 RECT 6.035 1.655 6.165 1.785 ;
 RECT 7.305 0.935 7.435 1.065 ;
 RECT 11.575 0.925 11.705 1.055 ;
 RECT 2.72 0.545 2.85 0.675 ;
 RECT 8.54 1.515 8.67 1.645 ;
 RECT 24.42 1.075 24.55 1.205 ;
 RECT 12.255 0.625 12.385 0.755 ;
 RECT 26.13 0.26 26.26 0.39 ;
 RECT 23.11 0.635 23.24 0.765 ;
 RECT 10.55 2.34 10.68 2.47 ;
 RECT 22.525 0.26 22.655 0.39 ;
 RECT 14.17 1.43 14.3 1.56 ;
 RECT 27.27 1.03 27.4 1.16 ;
 RECT 12.98 0.495 13.11 0.625 ;
 RECT 15.32 2.075 15.45 2.205 ;
 RECT 16.845 0.26 16.975 0.39 ;
 RECT 16.3 0.6 16.43 0.73 ;
 RECT 27.305 2.31 27.435 2.44 ;
 RECT 24.865 1.035 24.995 1.165 ;
 RECT 6.74 1.66 6.87 1.79 ;
 RECT 12.175 1.445 12.305 1.575 ;
 RECT 1.28 2.05 1.41 2.18 ;
 RECT 1.755 1.995 1.885 2.125 ;
 RECT 14.475 1.835 14.605 1.965 ;
 RECT 9.545 0.62 9.675 0.75 ;
 RECT 13.535 1.835 13.665 1.965 ;
 RECT 16.45 1.705 16.58 1.835 ;
 RECT 11.485 0.595 11.615 0.725 ;
 RECT 18.96 2.64 19.09 2.77 ;
 RECT 3.805 1.525 3.935 1.655 ;
 RECT 11.485 1.87 11.615 2 ;
 RECT 5.875 0.315 6.005 0.445 ;
 RECT 25.965 0.595 26.095 0.725 ;
 RECT 4.925 2.11 5.055 2.24 ;
 RECT 6.415 2.045 6.545 2.175 ;
 RECT 0.81 2.115 0.94 2.245 ;
 RECT 7.73 2.015 7.86 2.145 ;
 RECT 25.025 0.435 25.155 0.565 ;
 RECT 1.28 0.74 1.41 0.87 ;
 RECT 9.355 2.225 9.485 2.355 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 25.025 1.485 25.155 1.615 ;
 RECT 26.475 1.49 26.605 1.62 ;
 RECT 22.07 0.63 22.2 0.76 ;
 RECT 3.525 0.88 3.655 1.01 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 9.255 1.195 9.385 1.325 ;
 RECT 1.88 0.975 2.01 1.105 ;
 RECT 25.46 0.12 25.59 0.25 ;
 RECT 4.13 0.53 4.26 0.66 ;
 RECT 0.88 0.325 1.01 0.455 ;
 RECT 23.525 0.505 23.655 0.635 ;
 RECT 18.555 1.705 18.685 1.835 ;
 RECT 8.21 0.905 8.34 1.035 ;
 RECT 17.955 2.64 18.085 2.77 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 3.055 0.88 3.185 1.01 ;
 RECT 3.01 2.105 3.14 2.235 ;
 RECT 2.775 1.49 2.905 1.62 ;
 RECT 1.875 1.495 2.005 1.625 ;
 RECT 3.975 2.11 4.105 2.24 ;
 RECT 12.38 2.38 12.51 2.51 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 15.505 1.705 15.635 1.835 ;
 RECT 24.245 0.135 24.375 0.265 ;
 RECT 10.98 1.9 11.11 2.03 ;
 RECT 27.42 0.595 27.55 0.725 ;
 RECT 25.63 1.445 25.76 1.575 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 26.105 1.405 26.235 1.535 ;
 RECT 4.455 1.825 4.585 1.955 ;
 RECT 5.395 2.135 5.525 2.265 ;
 RECT 7.735 0.905 7.865 1.035 ;
 RECT 8.21 2.07 8.34 2.2 ;
 RECT 27.42 1.465 27.55 1.595 ;
 RECT 21.005 1.71 21.135 1.84 ;
 RECT 14.51 1.035 14.64 1.165 ;
 RECT 1.4 1.55 1.53 1.68 ;
 RECT 2.66 0.935 2.79 1.065 ;
 RECT 17.55 0.975 17.68 1.105 ;
 RECT 16.57 0.92 16.7 1.05 ;
 RECT 15.095 0.91 15.225 1.04 ;
 RECT 22.07 1.71 22.2 1.84 ;
 RECT 19.53 1.705 19.66 1.835 ;
 RECT 23.775 1.425 23.905 1.555 ;
 RECT 20.505 0.62 20.635 0.75 ;
 RECT 4.74 0.32 4.87 0.45 ;
 LAYER M1 ;
 RECT 4.465 1.25 7.865 1.365 ;
 RECT 6.975 1.365 7.865 1.39 ;
 RECT 7.66 0.9 7.935 1.04 ;
 RECT 3.345 1.82 4.925 1.96 ;
 RECT 4.785 1.79 4.925 1.82 ;
 RECT 3.345 1.22 3.66 1.36 ;
 RECT 3.52 0.805 3.66 1.22 ;
 RECT 3.43 1.96 3.71 2.215 ;
 RECT 3.345 1.36 3.485 1.82 ;
 RECT 5.985 1.615 6.215 1.65 ;
 RECT 5.985 1.79 6.215 1.825 ;
 RECT 4.785 1.65 6.22 1.79 ;
 RECT 1.795 1.63 1.935 1.99 ;
 RECT 1.795 1.475 2.1 1.63 ;
 RECT 1.875 0.905 2.015 1.475 ;
 RECT 1.685 1.99 1.935 2.13 ;
 RECT 25.96 0.73 26.1 1.04 ;
 RECT 26.1 1.18 26.24 1.605 ;
 RECT 25.895 0.59 26.17 0.73 ;
 RECT 27.22 0.99 27.45 1.04 ;
 RECT 25.96 1.04 27.45 1.18 ;
 RECT 27.22 1.18 27.45 1.2 ;
 RECT 26.08 0.29 26.45 0.43 ;
 RECT 26.31 0.43 26.45 0.71 ;
 RECT 26.08 0.22 26.31 0.29 ;
 RECT 27.73 0.85 27.87 1.385 ;
 RECT 27.415 1.525 27.555 1.73 ;
 RECT 26.31 0.71 27.87 0.85 ;
 RECT 27.415 0.51 27.555 0.71 ;
 RECT 27.415 1.385 27.87 1.525 ;
 RECT 25.34 1.145 25.48 1.345 ;
 RECT 25.02 1.485 25.16 1.76 ;
 RECT 25.34 0.73 25.48 0.935 ;
 RECT 25.02 0.355 25.16 0.59 ;
 RECT 25.02 1.345 25.48 1.485 ;
 RECT 25.295 0.935 25.525 1.145 ;
 RECT 25.02 0.59 25.48 0.73 ;
 RECT 23.32 1.225 23.55 1.245 ;
 RECT 23.32 1.195 23.91 1.225 ;
 RECT 23.46 1.015 23.77 1.035 ;
 RECT 23.32 1.035 23.77 1.055 ;
 RECT 23.595 0.64 23.735 1.015 ;
 RECT 23.77 1.225 23.91 1.75 ;
 RECT 23.475 0.5 23.735 0.64 ;
 RECT 24.37 1.035 24.6 1.055 ;
 RECT 24.37 1.195 24.6 1.245 ;
 RECT 23.32 1.055 24.6 1.195 ;
 RECT 22.475 0.36 22.705 0.43 ;
 RECT 22.475 0.22 24.015 0.36 ;
 RECT 23.875 0.36 24.015 0.565 ;
 RECT 24.615 0.705 24.755 0.75 ;
 RECT 24.74 0.995 25.045 1.205 ;
 RECT 24.74 0.89 24.88 0.995 ;
 RECT 24.615 0.75 24.88 0.89 ;
 RECT 23.875 0.565 24.755 0.705 ;
 RECT 15.525 0.775 15.665 1.405 ;
 RECT 16.25 0.56 16.48 0.635 ;
 RECT 14.505 1.405 15.665 1.545 ;
 RECT 14.505 1.545 14.645 1.83 ;
 RECT 14.505 1.17 14.645 1.405 ;
 RECT 13.46 1.83 14.71 1.97 ;
 RECT 14.435 1.03 14.715 1.17 ;
 RECT 19.54 0.36 19.68 0.635 ;
 RECT 15.525 0.635 19.68 0.775 ;
 RECT 20.22 0.36 20.36 1.46 ;
 RECT 19.54 0.22 20.36 0.36 ;
 RECT 12.205 0.585 13.16 0.63 ;
 RECT 12.205 0.63 12.435 0.795 ;
 RECT 12.23 0.49 13.16 0.585 ;
 RECT 12.93 0.455 13.16 0.49 ;
 RECT 12.93 0.63 13.16 0.665 ;
 RECT 13.785 0.57 14.015 0.95 ;
 RECT 16.795 0.22 17.025 0.28 ;
 RECT 16.795 0.42 17.025 0.43 ;
 RECT 14.63 0.28 17.025 0.42 ;
 RECT 14.63 0.42 14.86 0.6 ;
 RECT 11.48 0.525 11.62 0.885 ;
 RECT 11.48 1.095 11.62 2.065 ;
 RECT 11.48 0.885 11.755 1.095 ;
 RECT 9 2.055 9.14 2.34 ;
 RECT 8.205 2.34 9.14 2.48 ;
 RECT 9.44 1.66 9.58 1.915 ;
 RECT 9 1.915 9.58 2.055 ;
 RECT 8.205 1.04 8.345 2.34 ;
 RECT 8.205 0.895 8.345 0.9 ;
 RECT 8.135 0.9 8.41 1.04 ;
 RECT 9.44 1.52 11.115 1.66 ;
 RECT 10.45 0.765 10.59 1.52 ;
 RECT 10.45 1.66 10.59 2.145 ;
 RECT 10.975 0.525 11.115 1.52 ;
 RECT 10.975 1.66 11.115 2.11 ;
 RECT 3.8 0.66 3.94 0.895 ;
 RECT 3.34 0.52 3.94 0.66 ;
 RECT 3.8 0.895 7.485 1.035 ;
 RECT 7.255 1.035 7.485 1.105 ;
 RECT 2.655 1.67 2.795 1.82 ;
 RECT 2.655 1.96 2.795 2.25 ;
 RECT 2.655 0.715 2.795 1.44 ;
 RECT 2.655 1.44 2.91 1.67 ;
 RECT 2.655 0.505 2.9 0.715 ;
 RECT 2.525 1.82 2.795 1.96 ;
 RECT 0.585 1.335 0.725 2.11 ;
 RECT 0.585 2.25 0.725 2.255 ;
 RECT 0.585 0.875 0.725 1.195 ;
 RECT 0.585 2.11 1.01 2.25 ;
 RECT 0.585 0.735 1.01 0.875 ;
 RECT 0.585 1.195 1.695 1.335 ;
 RECT 1.555 0.6 1.695 1.195 ;
 RECT 3.05 0.36 3.19 2.035 ;
 RECT 2.285 0.36 2.425 0.46 ;
 RECT 3.005 2.17 3.145 2.305 ;
 RECT 3.005 2.035 3.19 2.17 ;
 RECT 1.555 0.46 2.425 0.6 ;
 RECT 2.285 0.22 3.19 0.36 ;
 RECT 12.895 1.895 13.035 2.39 ;
 RECT 16.835 2.205 16.975 2.39 ;
 RECT 12.895 2.39 16.975 2.53 ;
 RECT 11.77 1.755 13.035 1.895 ;
 RECT 11.77 1.895 11.91 2.34 ;
 RECT 10.5 2.3 10.73 2.34 ;
 RECT 10.5 2.48 10.73 2.51 ;
 RECT 10.5 2.34 11.91 2.48 ;
 RECT 16.835 2.065 23.055 2.205 ;
 RECT 22.915 2.205 23.055 2.52 ;
 RECT 27.255 2.48 27.395 2.52 ;
 RECT 22.915 2.52 27.395 2.66 ;
 RECT 27.255 2.27 27.485 2.48 ;
 RECT 16.335 1.7 16.63 1.84 ;
 RECT 16.335 1.84 16.475 2.075 ;
 RECT 15.64 1.84 15.78 2.075 ;
 RECT 15.445 1.7 15.78 1.84 ;
 RECT 15.64 2.075 16.475 2.215 ;
 RECT 16.53 1.055 16.67 1.245 ;
 RECT 15.97 1.385 16.11 1.625 ;
 RECT 15.97 1.245 17.04 1.385 ;
 RECT 16.81 1.385 17.04 1.455 ;
 RECT 16.5 0.915 16.8 1.055 ;
 RECT 15.94 1.625 16.195 1.92 ;
 RECT 13.175 1.56 13.315 2.11 ;
 RECT 12.125 1.405 12.355 1.42 ;
 RECT 12.125 1.56 12.355 1.615 ;
 RECT 12.125 1.42 13.315 1.56 ;
 RECT 13.175 2.11 15.5 2.245 ;
 RECT 13.175 2.245 15.495 2.25 ;
 RECT 15.27 2.035 15.5 2.11 ;
 RECT 8.65 1.04 8.79 1.475 ;
 RECT 8.49 1.475 8.79 1.635 ;
 RECT 8.65 1.775 8.79 2.18 ;
 RECT 8.58 0.9 8.855 1.04 ;
 RECT 9.16 1.33 9.3 1.635 ;
 RECT 8.65 1.685 9.3 1.775 ;
 RECT 9.16 1.19 9.455 1.33 ;
 RECT 8.49 1.635 9.3 1.685 ;
 RECT 3.905 2.105 5.125 2.245 ;
 RECT 4.465 1.225 7.115 1.25 ;
 RECT 6.41 1.365 6.55 2.25 ;
 RECT 4.465 1.365 4.605 1.5 ;
 RECT 3.635 1.64 4.14 1.675 ;
 RECT 3.635 1.5 4.605 1.64 ;
 RECT 7.725 1.04 7.865 1.25 ;
 RECT 7.725 1.39 7.865 2.215 ;
 RECT 7.725 0.885 7.865 0.9 ;
 END
END RDFFSRASRX2

MACRO CGLNPRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8 BY 2.88 ;
 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.965 1.145 2.36 1.4 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.53 1.8 6.84 2.04 ;
 RECT 6.325 1.21 6.67 1.35 ;
 RECT 6.325 0.48 6.465 1.21 ;
 RECT 6.53 2.04 6.67 2.45 ;
 RECT 6.53 1.35 6.67 1.8 ;
 END
 ANTENNADIFFAREA 0.61 ;
 END GCLK

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.415 1.415 1.755 1.72 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END SE

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.185 2.05 0.445 2.36 ;
 END
 ANTENNAGATEAREA 0.063 ;
 END CLK

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8 2.96 ;
 RECT 1.55 2.625 1.78 2.8 ;
 RECT 0.585 1.635 0.725 2.8 ;
 RECT 7 1.43 7.14 2.8 ;
 RECT 6.06 1.695 6.2 2.8 ;
 RECT 7.48 2.25 7.62 2.8 ;
 RECT 7.495 1.5 7.635 2.065 ;
 RECT 7.48 2.065 7.635 2.25 ;
 RECT 3.605 1.71 3.745 1.945 ;
 RECT 3.605 1.945 5.055 2.085 ;
 RECT 4.915 2.085 5.055 2.8 ;
 RECT 4.915 1.44 5.055 1.945 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8 0.08 ;
 RECT 1.895 0.08 2.035 0.725 ;
 RECT 4.915 0.08 5.055 0.68 ;
 RECT 0.585 0.08 0.725 0.975 ;
 RECT 6.795 0.08 6.935 0.98 ;
 RECT 5.855 0.08 5.995 0.68 ;
 RECT 3.605 0.08 3.745 0.74 ;
 RECT 7.46 0.08 7.6 0.85 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 5.64 0.28 5.74 0.75 ;
 RECT 5.475 1.275 5.575 2.22 ;
 RECT 5.475 0.85 5.575 1.065 ;
 RECT 5.475 0.75 5.74 0.85 ;
 RECT 5.455 1.065 5.685 1.275 ;
 RECT 2.62 0.19 2.72 0.885 ;
 RECT 1.27 0.19 1.5 0.395 ;
 RECT 1.27 0.09 2.72 0.19 ;
 RECT 2.62 1.26 2.72 2.35 ;
 RECT 3.09 0.315 3.19 0.89 ;
 RECT 3.01 0.89 3.19 0.99 ;
 RECT 3.01 0.99 3.11 1.16 ;
 RECT 2.62 1.16 3.11 1.26 ;
 RECT 2.51 2.35 2.72 2.58 ;
 RECT 5.885 1.04 6.21 1.25 ;
 RECT 6.11 0.25 6.21 1.04 ;
 RECT 6.11 1.25 6.21 1.255 ;
 RECT 6.58 0.25 6.68 1.255 ;
 RECT 6.785 1.355 6.885 2.74 ;
 RECT 6.315 1.355 6.415 2.745 ;
 RECT 6.11 1.255 6.885 1.355 ;
 RECT 2.91 2.03 3.19 2.24 ;
 RECT 3.09 1.56 3.19 2.03 ;
 RECT 2.15 1.32 2.25 2.14 ;
 RECT 2.15 0.37 2.25 1.11 ;
 RECT 1.97 1.11 2.25 1.32 ;
 RECT 1.495 0.955 1.595 1.43 ;
 RECT 1.68 0.37 1.78 0.855 ;
 RECT 1.85 1.64 1.95 2.14 ;
 RECT 1.465 1.43 1.695 1.54 ;
 RECT 1.465 1.54 1.95 1.64 ;
 RECT 1.495 0.855 1.78 0.955 ;
 RECT 4.7 0.2 4.8 1.85 ;
 RECT 3.39 0.2 3.49 1.17 ;
 RECT 3.39 1.38 3.49 2.14 ;
 RECT 3.39 0.1 4.8 0.2 ;
 RECT 3.29 1.17 3.52 1.38 ;
 RECT 5.17 0.28 5.27 2.38 ;
 RECT 4.545 2.34 4.775 2.38 ;
 RECT 4.545 2.48 4.775 2.55 ;
 RECT 4.545 2.38 5.27 2.48 ;
 RECT 3.705 0.89 3.96 1.1 ;
 RECT 3.86 0.38 3.96 0.89 ;
 RECT 3.86 1.1 3.96 2.14 ;
 RECT 0.37 0.57 0.47 2.05 ;
 RECT 0.205 2.05 0.47 2.26 ;
 RECT 0.68 1.12 0.94 1.33 ;
 RECT 0.84 0.565 0.94 1.12 ;
 RECT 0.84 1.33 0.94 2.345 ;
 RECT 0.84 2.345 1.095 2.555 ;
 LAYER CO ;
 RECT 7.005 1.48 7.135 1.61 ;
 RECT 2.55 2.4 2.68 2.53 ;
 RECT 2.96 2.07 3.09 2.2 ;
 RECT 7.465 0.41 7.595 0.54 ;
 RECT 5.86 0.5 5.99 0.63 ;
 RECT 1.9 0.545 2.03 0.675 ;
 RECT 0.59 0.79 0.72 0.92 ;
 RECT 3.34 1.21 3.47 1.34 ;
 RECT 6.535 2.01 6.665 2.14 ;
 RECT 1.06 0.79 1.19 0.92 ;
 RECT 4.08 0.6 4.21 0.73 ;
 RECT 4.595 2.38 4.725 2.51 ;
 RECT 6.065 1.745 6.195 1.875 ;
 RECT 6.535 2.27 6.665 2.4 ;
 RECT 4.45 0.53 4.58 0.66 ;
 RECT 6.065 2.01 6.195 2.14 ;
 RECT 2.84 0.535 2.97 0.665 ;
 RECT 0.12 0.79 0.25 0.92 ;
 RECT 1.43 0.59 1.56 0.72 ;
 RECT 5.935 1.08 6.065 1.21 ;
 RECT 7.5 2.07 7.63 2.2 ;
 RECT 7.5 1.81 7.63 1.94 ;
 RECT 1.515 1.47 1.645 1.6 ;
 RECT 6.535 1.745 6.665 1.875 ;
 RECT 5.39 0.5 5.52 0.63 ;
 RECT 1.6 2.63 1.73 2.76 ;
 RECT 2.37 1.78 2.5 1.91 ;
 RECT 2.02 1.15 2.15 1.28 ;
 RECT 4.45 0.79 4.58 0.92 ;
 RECT 7.5 1.55 7.63 1.68 ;
 RECT 2.37 0.59 2.5 0.72 ;
 RECT 5.695 1.765 5.825 1.895 ;
 RECT 6.33 0.79 6.46 0.92 ;
 RECT 6.065 2.27 6.195 2.4 ;
 RECT 4.92 0.5 5.05 0.63 ;
 RECT 4.45 1.5 4.58 1.63 ;
 RECT 0.73 1.16 0.86 1.29 ;
 RECT 0.255 2.09 0.385 2.22 ;
 RECT 0.915 2.385 1.045 2.515 ;
 RECT 2.84 1.78 2.97 1.91 ;
 RECT 3.755 0.93 3.885 1.06 ;
 RECT 5.505 1.105 5.635 1.235 ;
 RECT 4.92 1.76 5.05 1.89 ;
 RECT 7.005 2.01 7.135 2.14 ;
 RECT 3.61 0.535 3.74 0.665 ;
 RECT 7.005 1.745 7.135 1.875 ;
 RECT 6.8 0.53 6.93 0.66 ;
 RECT 6.535 1.48 6.665 1.61 ;
 RECT 1.06 1.5 1.19 1.63 ;
 RECT 0.59 1.685 0.72 1.815 ;
 RECT 6.33 0.53 6.46 0.66 ;
 RECT 5.695 1.5 5.825 1.63 ;
 RECT 3.61 1.78 3.74 1.91 ;
 RECT 0.12 1.585 0.25 1.715 ;
 RECT 4.92 1.5 5.05 1.63 ;
 RECT 4.08 1.5 4.21 1.63 ;
 RECT 7.005 2.27 7.135 2.4 ;
 RECT 7.465 0.67 7.595 0.8 ;
 RECT 1.32 0.225 1.45 0.355 ;
 RECT 6.8 0.79 6.93 0.92 ;
 LAYER M1 ;
 RECT 5.385 0.45 5.525 0.82 ;
 RECT 5.69 1.54 5.83 1.945 ;
 RECT 5.825 0.96 5.965 1.075 ;
 RECT 5.825 1.215 5.965 1.4 ;
 RECT 5.385 0.82 5.965 0.96 ;
 RECT 5.69 1.4 5.965 1.54 ;
 RECT 5.825 1.075 6.115 1.215 ;
 RECT 4.445 0.44 4.585 1.1 ;
 RECT 4.445 1.24 4.585 1.68 ;
 RECT 4.445 1.1 5.685 1.24 ;
 RECT 1.425 0.53 1.565 0.865 ;
 RECT 2.51 1.625 2.65 1.775 ;
 RECT 1.425 0.865 2.87 1.005 ;
 RECT 2.73 1.005 2.87 1.485 ;
 RECT 2.365 0.53 2.505 0.865 ;
 RECT 2.32 1.775 2.65 1.915 ;
 RECT 2.51 1.485 2.87 1.625 ;
 RECT 3.01 0.67 3.15 0.925 ;
 RECT 3.01 1.065 3.15 1.775 ;
 RECT 2.77 0.53 3.15 0.67 ;
 RECT 2.79 1.775 3.15 1.915 ;
 RECT 3.01 0.925 3.935 1.065 ;
 RECT 3.29 1.205 4.215 1.345 ;
 RECT 4.075 0.365 4.215 1.205 ;
 RECT 4.075 1.345 4.215 1.68 ;
 RECT 3.3 2.205 3.44 2.375 ;
 RECT 1.055 2.065 3.44 2.205 ;
 RECT 1.055 0.36 1.195 2.065 ;
 RECT 1.055 0.22 1.5 0.36 ;
 RECT 3.3 2.375 4.775 2.515 ;
 RECT 0.115 0.72 0.255 1.155 ;
 RECT 0.115 1.295 0.255 1.785 ;
 RECT 0.68 1.12 0.91 1.155 ;
 RECT 0.68 1.295 0.91 1.33 ;
 RECT 0.115 1.155 0.91 1.295 ;
 RECT 2.545 2.485 2.685 2.58 ;
 RECT 0.865 2.485 1.095 2.555 ;
 RECT 0.865 2.345 2.69 2.485 ;
 END
END CGLNPRX2

MACRO CGLNPRX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.2 BY 2.88 ;
 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.165 1.99 0.44 2.36 ;
 END
 ANTENNAGATEAREA 0.063 ;
 END CLK

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.2 2.96 ;
 RECT 0.54 1.57 0.77 1.71 ;
 RECT 1.53 2.615 1.8 2.8 ;
 RECT 6.435 1.43 6.575 2.8 ;
 RECT 7.375 1.43 7.515 2.8 ;
 RECT 8.315 1.43 8.455 2.8 ;
 RECT 5.295 1.735 5.435 2.8 ;
 RECT 9.255 1.43 9.395 2.8 ;
 RECT 10.195 1.43 10.335 2.8 ;
 RECT 10.655 1.5 10.795 2.8 ;
 RECT 0.585 1.71 0.725 2.8 ;
 RECT 3.605 1.655 3.745 1.86 ;
 RECT 4.915 2 5.055 2.8 ;
 RECT 3.605 1.86 5.055 2 ;
 RECT 4.915 1.44 5.055 1.86 ;
 END
 END VDD

 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.96 1.145 2.36 1.4 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.2 0.08 ;
 RECT 3.605 0.08 3.745 0.74 ;
 RECT 1.85 0.585 2.08 0.725 ;
 RECT 5.495 0.08 5.635 0.83 ;
 RECT 7.375 0.08 7.515 0.975 ;
 RECT 9.255 0.08 9.395 0.975 ;
 RECT 8.315 0.08 8.455 0.975 ;
 RECT 10.195 0.08 10.335 0.975 ;
 RECT 4.915 0.08 5.055 0.955 ;
 RECT 0.585 0.08 0.725 0.99 ;
 RECT 6.435 0.08 6.575 0.975 ;
 RECT 10.655 0.08 10.795 0.85 ;
 RECT 1.895 0.08 2.035 0.585 ;
 END
 END VSS

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.905 1.12 9.865 1.26 ;
 RECT 9.725 2.055 9.865 2.45 ;
 RECT 9.725 1.76 10.055 2.055 ;
 RECT 7.845 1.26 7.985 2.45 ;
 RECT 7.845 0.475 7.985 1.12 ;
 RECT 6.905 1.26 7.045 2.45 ;
 RECT 6.905 0.475 7.045 1.12 ;
 RECT 8.785 1.26 8.925 2.45 ;
 RECT 8.785 0.475 8.925 1.12 ;
 RECT 9.725 1.26 9.865 1.76 ;
 RECT 9.725 0.475 9.865 1.12 ;
 END
 ANTENNADIFFAREA 2.488 ;
 END GCLK

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.455 1.395 1.795 1.74 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END SE

 OBS
 LAYER PO ;
 RECT 2.62 0.19 2.72 0.885 ;
 RECT 1.12 0.19 1.35 0.395 ;
 RECT 1.12 0.09 2.72 0.19 ;
 RECT 4.7 0.2 4.8 1.85 ;
 RECT 3.39 0.2 3.49 1.07 ;
 RECT 3.39 1.28 3.49 2.14 ;
 RECT 3.39 0.1 4.8 0.2 ;
 RECT 3.29 1.07 3.52 1.28 ;
 RECT 2.15 0.37 2.25 1.11 ;
 RECT 2.15 1.32 2.25 2.14 ;
 RECT 1.97 1.11 2.25 1.32 ;
 RECT 4.675 2.55 4.775 2.69 ;
 RECT 5.75 0.37 5.85 1.03 ;
 RECT 5.55 1.13 5.65 2.69 ;
 RECT 4.545 2.34 4.775 2.55 ;
 RECT 5.55 1.03 5.85 1.13 ;
 RECT 4.675 2.69 5.65 2.79 ;
 RECT 6.22 0.19 6.32 1.31 ;
 RECT 5.18 0.19 5.39 0.45 ;
 RECT 5.85 1.41 5.95 2.79 ;
 RECT 5.18 0.09 6.32 0.19 ;
 RECT 5.85 1.31 6.32 1.41 ;
 RECT 6.525 1.08 6.79 1.15 ;
 RECT 6.525 1.25 6.79 1.29 ;
 RECT 6.69 1.29 6.79 2.74 ;
 RECT 6.69 0.215 6.79 1.08 ;
 RECT 9.04 1.25 9.14 2.74 ;
 RECT 9.04 0.215 9.14 1.15 ;
 RECT 8.1 1.25 8.2 2.74 ;
 RECT 8.1 0.215 8.2 1.15 ;
 RECT 7.16 1.25 7.26 2.74 ;
 RECT 7.16 0.215 7.26 1.15 ;
 RECT 9.51 1.25 9.61 2.74 ;
 RECT 9.51 0.215 9.61 1.15 ;
 RECT 9.98 0.215 10.08 1.15 ;
 RECT 9.98 1.25 10.08 2.74 ;
 RECT 8.57 0.215 8.67 1.15 ;
 RECT 8.57 1.25 8.67 2.74 ;
 RECT 7.63 0.215 7.73 1.15 ;
 RECT 7.63 1.25 7.73 2.74 ;
 RECT 6.525 1.15 10.08 1.25 ;
 RECT 2.93 2.03 3.19 2.24 ;
 RECT 3.09 1.5 3.19 2.03 ;
 RECT 3.86 0.38 3.96 2.145 ;
 RECT 3.855 2.145 4.085 2.355 ;
 RECT 1.85 1.61 1.95 2.14 ;
 RECT 1.56 1.51 1.95 1.61 ;
 RECT 1.68 0.37 1.78 1.4 ;
 RECT 1.56 1.4 1.79 1.51 ;
 RECT 0.68 1.13 0.94 1.34 ;
 RECT 0.84 0.185 0.94 1.13 ;
 RECT 0.84 1.34 0.94 2.31 ;
 RECT 0.84 2.31 1.105 2.505 ;
 RECT 0.875 2.505 1.105 2.52 ;
 RECT 3.01 0.76 3.19 0.885 ;
 RECT 3.01 0.885 3.11 1.16 ;
 RECT 2.62 1.26 2.72 2.365 ;
 RECT 3.09 0.315 3.19 0.76 ;
 RECT 2.62 1.16 3.11 1.26 ;
 RECT 2.515 2.365 2.745 2.575 ;
 RECT 0.37 0.57 0.47 1.99 ;
 RECT 0.195 1.99 0.47 2.2 ;
 LAYER CO ;
 RECT 7.38 1.745 7.51 1.875 ;
 RECT 7.38 2.27 7.51 2.4 ;
 RECT 3.61 1.73 3.74 1.86 ;
 RECT 10.2 2.27 10.33 2.4 ;
 RECT 7.85 2.01 7.98 2.14 ;
 RECT 1.9 0.59 2.03 0.72 ;
 RECT 8.32 2.01 8.45 2.14 ;
 RECT 6.07 1.53 6.2 1.66 ;
 RECT 8.32 1.745 8.45 1.875 ;
 RECT 7.38 1.48 7.51 1.61 ;
 RECT 4.45 0.79 4.58 0.92 ;
 RECT 8.79 1.745 8.92 1.875 ;
 RECT 8.32 0.525 8.45 0.655 ;
 RECT 8.79 2.27 8.92 2.4 ;
 RECT 7.85 0.785 7.98 0.915 ;
 RECT 8.79 1.48 8.92 1.61 ;
 RECT 9.26 0.525 9.39 0.655 ;
 RECT 6.91 1.745 7.04 1.875 ;
 RECT 0.73 1.17 0.86 1.3 ;
 RECT 3.905 2.185 4.035 2.315 ;
 RECT 1.61 1.44 1.74 1.57 ;
 RECT 0.925 2.35 1.055 2.48 ;
 RECT 2.565 2.405 2.695 2.535 ;
 RECT 0.245 2.03 0.375 2.16 ;
 RECT 10.66 1.55 10.79 1.68 ;
 RECT 7.85 1.48 7.98 1.61 ;
 RECT 5.3 1.795 5.43 1.925 ;
 RECT 6.91 0.785 7.04 0.915 ;
 RECT 4.92 1.5 5.05 1.63 ;
 RECT 2.84 1.73 2.97 1.86 ;
 RECT 10.66 0.41 10.79 0.54 ;
 RECT 1.06 0.79 1.19 0.92 ;
 RECT 5.97 0.655 6.1 0.785 ;
 RECT 10.2 0.525 10.33 0.655 ;
 RECT 5.3 2.32 5.43 2.45 ;
 RECT 9.73 0.785 9.86 0.915 ;
 RECT 6.44 1.48 6.57 1.61 ;
 RECT 2.84 0.535 2.97 0.665 ;
 RECT 6.44 1.745 6.57 1.875 ;
 RECT 6.91 1.48 7.04 1.61 ;
 RECT 6.91 0.525 7.04 0.655 ;
 RECT 8.79 0.525 8.92 0.655 ;
 RECT 4.595 2.38 4.725 2.51 ;
 RECT 0.59 0.79 0.72 0.92 ;
 RECT 6.575 1.12 6.705 1.25 ;
 RECT 5.5 0.65 5.63 0.78 ;
 RECT 1.17 0.225 1.3 0.355 ;
 RECT 6.44 0.785 6.57 0.915 ;
 RECT 1.43 0.59 1.56 0.72 ;
 RECT 6.07 2.06 6.2 2.19 ;
 RECT 9.73 0.525 9.86 0.655 ;
 RECT 8.79 2.01 8.92 2.14 ;
 RECT 6.91 2.01 7.04 2.14 ;
 RECT 4.92 0.775 5.05 0.905 ;
 RECT 6.44 2.27 6.57 2.4 ;
 RECT 8.32 0.785 8.45 0.915 ;
 RECT 9.26 2.01 9.39 2.14 ;
 RECT 9.26 0.785 9.39 0.915 ;
 RECT 9.26 1.745 9.39 1.875 ;
 RECT 9.73 1.745 9.86 1.875 ;
 RECT 9.73 2.27 9.86 2.4 ;
 RECT 8.32 2.27 8.45 2.4 ;
 RECT 9.73 1.48 9.86 1.61 ;
 RECT 6.44 2.01 6.57 2.14 ;
 RECT 3.61 0.535 3.74 0.665 ;
 RECT 7.38 2.01 7.51 2.14 ;
 RECT 7.85 0.525 7.98 0.655 ;
 RECT 2.37 1.73 2.5 1.86 ;
 RECT 10.2 2.01 10.33 2.14 ;
 RECT 7.85 1.745 7.98 1.875 ;
 RECT 8.32 1.48 8.45 1.61 ;
 RECT 10.2 1.48 10.33 1.61 ;
 RECT 8.79 0.785 8.92 0.915 ;
 RECT 9.26 2.27 9.39 2.4 ;
 RECT 5.22 0.27 5.35 0.4 ;
 RECT 4.08 0.6 4.21 0.73 ;
 RECT 7.85 2.27 7.98 2.4 ;
 RECT 4.45 0.53 4.58 0.66 ;
 RECT 3.34 1.11 3.47 1.24 ;
 RECT 2.02 1.15 2.15 1.28 ;
 RECT 0.12 0.79 0.25 0.92 ;
 RECT 4.08 1.5 4.21 1.63 ;
 RECT 5.3 2.06 5.43 2.19 ;
 RECT 2.37 0.59 2.5 0.72 ;
 RECT 10.66 2.07 10.79 2.2 ;
 RECT 0.59 1.58 0.72 1.71 ;
 RECT 0.12 1.585 0.25 1.715 ;
 RECT 7.38 0.785 7.51 0.915 ;
 RECT 4.92 0.515 5.05 0.645 ;
 RECT 10.66 1.81 10.79 1.94 ;
 RECT 9.73 2.01 9.86 2.14 ;
 RECT 2.98 2.07 3.11 2.2 ;
 RECT 10.66 0.67 10.79 0.8 ;
 RECT 10.2 1.745 10.33 1.875 ;
 RECT 6.07 1.795 6.2 1.925 ;
 RECT 4.45 1.5 4.58 1.63 ;
 RECT 1.6 2.62 1.73 2.75 ;
 RECT 1.06 1.5 1.19 1.63 ;
 RECT 7.38 0.525 7.51 0.655 ;
 RECT 6.91 2.27 7.04 2.4 ;
 RECT 10.2 0.785 10.33 0.915 ;
 RECT 6.44 0.495 6.57 0.625 ;
 RECT 9.26 1.48 9.39 1.61 ;
 LAYER M1 ;
 RECT 4.075 0.365 4.215 1.105 ;
 RECT 3.29 1.105 4.215 1.245 ;
 RECT 4.075 1.245 4.215 1.68 ;
 RECT 5.965 0.595 6.105 1.12 ;
 RECT 6.065 1.26 6.205 2.275 ;
 RECT 5.965 1.12 6.755 1.255 ;
 RECT 5.965 1.255 6.71 1.26 ;
 RECT 6.525 1.115 6.755 1.12 ;
 RECT 6.57 1.26 6.71 1.27 ;
 RECT 1.425 0.53 1.565 0.865 ;
 RECT 2.365 0.53 2.505 0.865 ;
 RECT 2.32 1.725 2.65 1.865 ;
 RECT 2.51 1.005 2.65 1.725 ;
 RECT 1.425 0.865 2.65 1.005 ;
 RECT 1.055 0.36 1.195 2.025 ;
 RECT 1.055 0.22 1.35 0.36 ;
 RECT 1.055 2.03 3.16 2.165 ;
 RECT 1.055 2.025 3.13 2.03 ;
 RECT 3.02 2.205 3.16 2.51 ;
 RECT 2.93 2.165 3.16 2.205 ;
 RECT 3.02 2.51 4.775 2.515 ;
 RECT 3.02 2.515 4.77 2.65 ;
 RECT 4.545 2.375 4.775 2.51 ;
 RECT 4.445 0.44 4.585 1.1 ;
 RECT 4.445 1.24 4.585 1.68 ;
 RECT 4.445 1.1 5.355 1.24 ;
 RECT 5.215 0.22 5.355 1.1 ;
 RECT 0.115 0.72 0.255 1.165 ;
 RECT 0.115 1.305 0.255 1.79 ;
 RECT 0.68 1.13 0.91 1.165 ;
 RECT 0.68 1.305 0.91 1.34 ;
 RECT 0.115 1.165 0.91 1.305 ;
 RECT 2.79 1.725 3.45 1.865 ;
 RECT 3.31 1.865 3.45 2.23 ;
 RECT 2.835 0.455 2.975 1.725 ;
 RECT 3.855 2.145 4.085 2.23 ;
 RECT 3.31 2.23 4.085 2.37 ;
 RECT 0.875 2.475 1.105 2.525 ;
 RECT 0.875 2.31 1.105 2.335 ;
 RECT 0.875 2.335 2.745 2.475 ;
 RECT 2.48 2.475 2.745 2.605 ;
 END
END CGLNPRX8

MACRO CGLNPSX16
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 15.36 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.725 0.805 5.085 1.14 ;
 END
 ANTENNAGATEAREA 0.051 ;
 END SE

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 15.36 0.08 ;
 RECT 5.82 0.585 6.05 0.725 ;
 RECT 1.375 0.585 1.63 0.725 ;
 RECT 1.49 0.08 1.63 0.585 ;
 RECT 12.445 0.08 12.585 0.98 ;
 RECT 11.505 0.08 11.645 0.98 ;
 RECT 6.805 0.08 6.945 0.73 ;
 RECT 13.385 0.08 13.525 0.98 ;
 RECT 4.925 0.08 5.065 0.58 ;
 RECT 9.625 0.08 9.765 0.98 ;
 RECT 3.975 0.08 4.115 0.715 ;
 RECT 7.745 0.08 7.885 0.98 ;
 RECT 0.585 0.08 0.725 0.985 ;
 RECT 8.685 0.08 8.825 0.98 ;
 RECT 10.565 0.08 10.705 0.98 ;
 RECT 14.325 0.08 14.465 0.98 ;
 RECT 3.135 0.08 3.275 0.74 ;
 RECT 5.865 0.725 6.005 0.735 ;
 RECT 5.865 0.08 6.005 0.585 ;
 RECT 14.855 0.08 14.995 0.85 ;
 END
 END VSS

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.035 1.79 11.345 2.055 ;
 RECT 7.465 1.15 13.995 1.29 ;
 RECT 7.275 0.805 7.605 0.945 ;
 RECT 7.275 1.43 7.605 1.57 ;
 RECT 7.275 0.43 7.415 0.805 ;
 RECT 7.275 1.57 7.415 2.22 ;
 RECT 11.035 2.055 11.175 2.455 ;
 RECT 11.035 0.45 11.175 1.15 ;
 RECT 13.855 1.29 13.995 2.455 ;
 RECT 13.855 0.455 13.995 1.15 ;
 RECT 7.465 0.945 7.605 1.15 ;
 RECT 11.975 1.29 12.115 2.455 ;
 RECT 11.975 0.455 12.115 1.15 ;
 RECT 7.465 1.29 7.605 1.43 ;
 RECT 10.095 1.29 10.235 2.455 ;
 RECT 10.095 0.455 10.235 1.15 ;
 RECT 9.155 1.29 9.295 2.455 ;
 RECT 9.155 0.45 9.295 1.15 ;
 RECT 12.915 1.29 13.055 2.455 ;
 RECT 12.915 0.45 13.055 1.15 ;
 RECT 8.215 1.29 8.355 2.455 ;
 RECT 8.215 0.455 8.355 1.15 ;
 RECT 11.035 1.29 11.175 1.79 ;
 END
 ANTENNADIFFAREA 4.72 ;
 END GCLK

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 15.36 2.96 ;
 RECT 1.31 2.41 1.58 2.55 ;
 RECT 3.09 2.625 3.32 2.8 ;
 RECT 4.915 1.675 5.055 2.8 ;
 RECT 0.585 1.575 0.725 2.8 ;
 RECT 14.325 1.435 14.465 2.8 ;
 RECT 9.625 1.435 9.765 2.8 ;
 RECT 13.385 1.435 13.525 2.8 ;
 RECT 7.745 1.435 7.885 2.8 ;
 RECT 12.445 1.435 12.585 2.8 ;
 RECT 6.805 1.72 6.945 2.8 ;
 RECT 10.565 1.435 10.705 2.8 ;
 RECT 11.505 1.435 11.645 2.8 ;
 RECT 8.685 1.435 8.825 2.8 ;
 RECT 1.375 2.55 1.515 2.8 ;
 RECT 14.89 1.5 15.03 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.405 1.16 0.76 1.4 ;
 END
 ANTENNAGATEAREA 0.063 ;
 END CLK

 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 1.44 1.75 1.72 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 OBS
 LAYER PO ;
 RECT 4.7 1.065 4.8 1.85 ;
 RECT 4.7 0.28 4.8 0.855 ;
 RECT 4.7 0.855 4.955 1.065 ;
 RECT 2.92 0.315 3.02 1.17 ;
 RECT 2.92 1.38 3.02 2.14 ;
 RECT 2.82 1.17 3.05 1.38 ;
 RECT 4.23 1.1 4.33 1.28 ;
 RECT 4.4 1.38 4.5 1.85 ;
 RECT 4.23 0.28 4.33 0.89 ;
 RECT 4.05 0.89 4.33 1.1 ;
 RECT 4.23 1.28 4.5 1.38 ;
 RECT 5.49 1.235 6.215 1.335 ;
 RECT 6.115 1.13 6.215 1.235 ;
 RECT 6.115 1.335 6.215 2.79 ;
 RECT 5.49 1.15 5.75 1.235 ;
 RECT 5.49 1.335 5.74 1.36 ;
 RECT 5.64 1.36 5.74 2.79 ;
 RECT 6.115 1.055 6.22 1.13 ;
 RECT 6.12 0.37 6.22 1.055 ;
 RECT 5.65 0.37 5.75 1.15 ;
 RECT 1.68 0.37 1.78 1.44 ;
 RECT 1.68 1.65 1.78 2.14 ;
 RECT 1.52 1.44 1.78 1.65 ;
 RECT 2.15 0.19 2.25 0.885 ;
 RECT 1.12 0.09 2.25 0.19 ;
 RECT 1.12 0.19 1.35 0.4 ;
 RECT 6.59 0.19 6.69 2.79 ;
 RECT 5.17 0.96 5.27 2.69 ;
 RECT 5.18 0.19 5.28 0.865 ;
 RECT 5.17 0.865 5.28 0.96 ;
 RECT 4.55 2.425 4.785 2.655 ;
 RECT 4.685 2.655 4.785 2.69 ;
 RECT 5.18 0.09 6.69 0.19 ;
 RECT 4.685 2.69 5.27 2.79 ;
 RECT 3.39 1.1 3.49 2.14 ;
 RECT 3.39 0.38 3.49 0.89 ;
 RECT 3.235 0.89 3.49 1.1 ;
 RECT 7.06 0.28 7.16 1.09 ;
 RECT 7.06 1.3 7.16 2.745 ;
 RECT 9.41 0.28 9.51 1.175 ;
 RECT 9.41 1.275 9.51 2.745 ;
 RECT 12.7 0.28 12.8 1.175 ;
 RECT 12.7 1.275 12.8 2.745 ;
 RECT 10.82 0.28 10.92 1.175 ;
 RECT 10.82 1.275 10.92 2.745 ;
 RECT 13.64 0.28 13.74 1.175 ;
 RECT 13.64 1.275 13.74 2.745 ;
 RECT 8.94 0.28 9.04 1.175 ;
 RECT 8.94 1.275 9.04 2.745 ;
 RECT 11.76 0.28 11.86 1.175 ;
 RECT 11.76 1.275 11.86 2.745 ;
 RECT 13.17 0.28 13.27 1.175 ;
 RECT 13.17 1.275 13.27 2.745 ;
 RECT 11.29 0.28 11.39 1.175 ;
 RECT 11.29 1.275 11.39 2.745 ;
 RECT 9.88 0.28 9.98 1.175 ;
 RECT 9.88 1.275 9.98 2.745 ;
 RECT 7.53 0.28 7.63 1.175 ;
 RECT 7.53 1.275 7.63 2.745 ;
 RECT 14.11 0.28 14.21 1.175 ;
 RECT 14.11 1.275 14.21 2.745 ;
 RECT 12.23 0.28 12.33 1.175 ;
 RECT 12.23 1.275 12.33 2.745 ;
 RECT 10.35 0.28 10.45 1.175 ;
 RECT 10.35 1.275 10.45 2.745 ;
 RECT 8.47 0.28 8.57 1.175 ;
 RECT 8.47 1.275 8.57 2.745 ;
 RECT 8 0.28 8.1 1.175 ;
 RECT 8 1.275 8.1 2.745 ;
 RECT 7.06 1.09 7.29 1.175 ;
 RECT 7.06 1.275 7.29 1.3 ;
 RECT 7.06 1.175 14.21 1.275 ;
 RECT 2.62 1.56 2.72 2.095 ;
 RECT 2.455 2.095 2.72 2.305 ;
 RECT 2.15 1.26 2.25 2.645 ;
 RECT 0.84 0.28 0.94 2.305 ;
 RECT 2.62 0.315 2.72 0.89 ;
 RECT 0.84 2.405 0.94 2.645 ;
 RECT 0.115 2.305 0.94 2.405 ;
 RECT 0.115 2.24 0.345 2.305 ;
 RECT 0.115 2.405 0.345 2.45 ;
 RECT 2.54 0.89 2.72 0.99 ;
 RECT 2.54 0.99 2.64 1.16 ;
 RECT 2.15 1.16 2.64 1.26 ;
 RECT 0.84 2.645 2.25 2.745 ;
 RECT 0.37 1.16 0.635 1.37 ;
 RECT 0.37 1.37 0.47 2.06 ;
 RECT 0.37 0.57 0.47 1.16 ;
 LAYER CO ;
 RECT 0.455 1.2 0.585 1.33 ;
 RECT 6.335 1.775 6.465 1.905 ;
 RECT 8.22 1.75 8.35 1.88 ;
 RECT 7.75 0.505 7.88 0.635 ;
 RECT 8.22 0.765 8.35 0.895 ;
 RECT 4.93 0.4 5.06 0.53 ;
 RECT 7.28 0.5 7.41 0.63 ;
 RECT 8.22 1.485 8.35 1.615 ;
 RECT 13.86 2.275 13.99 2.405 ;
 RECT 12.45 1.75 12.58 1.88 ;
 RECT 12.45 2.015 12.58 2.145 ;
 RECT 14.33 2.015 14.46 2.145 ;
 RECT 0.12 0.79 0.25 0.92 ;
 RECT 11.98 0.765 12.11 0.895 ;
 RECT 7.28 1.485 7.41 1.615 ;
 RECT 2.37 0.535 2.5 0.665 ;
 RECT 1.38 2.415 1.51 2.545 ;
 RECT 5.865 1.77 5.995 1.9 ;
 RECT 7.75 1.485 7.88 1.615 ;
 RECT 9.63 1.75 9.76 1.88 ;
 RECT 11.51 2.015 11.64 2.145 ;
 RECT 8.22 2.015 8.35 2.145 ;
 RECT 12.92 2.275 13.05 2.405 ;
 RECT 14.33 1.75 14.46 1.88 ;
 RECT 11.98 2.015 12.11 2.145 ;
 RECT 10.1 0.505 10.23 0.635 ;
 RECT 11.04 2.275 11.17 2.405 ;
 RECT 12.92 2.015 13.05 2.145 ;
 RECT 10.1 2.015 10.23 2.145 ;
 RECT 4.15 1.5 4.28 1.63 ;
 RECT 3.61 0.6 3.74 0.73 ;
 RECT 14.86 0.67 14.99 0.8 ;
 RECT 10.1 1.485 10.23 1.615 ;
 RECT 6.81 2.035 6.94 2.165 ;
 RECT 7.28 1.75 7.41 1.88 ;
 RECT 9.63 0.505 9.76 0.635 ;
 RECT 9.16 0.765 9.29 0.895 ;
 RECT 8.69 2.275 8.82 2.405 ;
 RECT 8.69 1.75 8.82 1.88 ;
 RECT 13.86 1.485 13.99 1.615 ;
 RECT 13.39 0.505 13.52 0.635 ;
 RECT 11.51 0.765 11.64 0.895 ;
 RECT 14.33 0.765 14.46 0.895 ;
 RECT 1.9 0.59 2.03 0.72 ;
 RECT 12.92 0.765 13.05 0.895 ;
 RECT 10.57 2.275 10.7 2.405 ;
 RECT 1.17 0.23 1.3 0.36 ;
 RECT 1.06 0.79 1.19 0.92 ;
 RECT 9.63 2.015 9.76 2.145 ;
 RECT 14.86 0.41 14.99 0.54 ;
 RECT 12.92 1.485 13.05 1.615 ;
 RECT 6.81 0.55 6.94 0.68 ;
 RECT 5.39 2.035 5.52 2.165 ;
 RECT 10.57 0.505 10.7 0.635 ;
 RECT 13.39 0.765 13.52 0.895 ;
 RECT 7.75 2.015 7.88 2.145 ;
 RECT 10.57 2.015 10.7 2.145 ;
 RECT 8.69 0.765 8.82 0.895 ;
 RECT 13.39 1.75 13.52 1.88 ;
 RECT 10.57 1.75 10.7 1.88 ;
 RECT 14.33 0.505 14.46 0.635 ;
 RECT 13.86 0.765 13.99 0.895 ;
 RECT 9.16 0.5 9.29 0.63 ;
 RECT 0.12 1.585 0.25 1.715 ;
 RECT 1.43 0.59 1.56 0.72 ;
 RECT 5.87 0.59 6 0.72 ;
 RECT 5.4 0.405 5.53 0.535 ;
 RECT 11.51 1.485 11.64 1.615 ;
 RECT 11.04 2.015 11.17 2.145 ;
 RECT 13.39 1.485 13.52 1.615 ;
 RECT 1.9 1.78 2.03 1.91 ;
 RECT 9.63 0.765 9.76 0.895 ;
 RECT 10.57 1.485 10.7 1.615 ;
 RECT 11.98 1.485 12.11 1.615 ;
 RECT 11.98 0.505 12.11 0.635 ;
 RECT 7.11 1.13 7.24 1.26 ;
 RECT 12.92 1.75 13.05 1.88 ;
 RECT 4.45 0.53 4.58 0.66 ;
 RECT 8.69 2.015 8.82 2.145 ;
 RECT 10.1 0.765 10.23 0.895 ;
 RECT 6.81 2.295 6.94 2.425 ;
 RECT 1.57 1.48 1.7 1.61 ;
 RECT 8.22 2.275 8.35 2.405 ;
 RECT 14.895 1.81 15.025 1.94 ;
 RECT 13.86 2.015 13.99 2.145 ;
 RECT 14.895 1.55 15.025 1.68 ;
 RECT 4.6 2.47 4.73 2.6 ;
 RECT 5.865 2.03 5.995 2.16 ;
 RECT 12.45 0.505 12.58 0.635 ;
 RECT 9.16 2.275 9.29 2.405 ;
 RECT 7.75 0.765 7.88 0.895 ;
 RECT 13.39 2.275 13.52 2.405 ;
 RECT 5.39 1.775 5.52 1.905 ;
 RECT 13.39 2.015 13.52 2.145 ;
 RECT 4.775 0.895 4.905 1.025 ;
 RECT 3.61 1.78 3.74 1.91 ;
 RECT 3.98 0.53 4.11 0.66 ;
 RECT 8.69 1.485 8.82 1.615 ;
 RECT 7.75 2.275 7.88 2.405 ;
 RECT 12.45 1.485 12.58 1.615 ;
 RECT 6.34 0.59 6.47 0.72 ;
 RECT 10.57 0.765 10.7 0.895 ;
 RECT 14.33 1.485 14.46 1.615 ;
 RECT 9.16 1.75 9.29 1.88 ;
 RECT 12.45 2.275 12.58 2.405 ;
 RECT 4.92 1.775 5.05 1.905 ;
 RECT 11.04 0.765 11.17 0.895 ;
 RECT 6.81 1.77 6.94 1.9 ;
 RECT 9.16 1.485 9.29 1.615 ;
 RECT 14.33 2.275 14.46 2.405 ;
 RECT 8.22 0.505 8.35 0.635 ;
 RECT 5.865 1.51 5.995 1.64 ;
 RECT 0.59 0.79 0.72 0.92 ;
 RECT 3.14 0.535 3.27 0.665 ;
 RECT 2.37 1.78 2.5 1.91 ;
 RECT 10.1 2.275 10.23 2.405 ;
 RECT 2.87 1.21 3 1.34 ;
 RECT 11.98 1.75 12.11 1.88 ;
 RECT 11.04 0.5 11.17 0.63 ;
 RECT 11.51 2.275 11.64 2.405 ;
 RECT 13.86 1.75 13.99 1.88 ;
 RECT 7.28 2.015 7.41 2.145 ;
 RECT 5.54 1.19 5.67 1.32 ;
 RECT 4.1 0.93 4.23 1.06 ;
 RECT 3.285 0.93 3.415 1.06 ;
 RECT 3.14 2.63 3.27 2.76 ;
 RECT 2.505 2.135 2.635 2.265 ;
 RECT 0.165 2.28 0.295 2.41 ;
 RECT 7.75 1.75 7.88 1.88 ;
 RECT 9.63 2.275 9.76 2.405 ;
 RECT 11.04 1.75 11.17 1.88 ;
 RECT 0.59 1.625 0.72 1.755 ;
 RECT 12.45 0.765 12.58 0.895 ;
 RECT 11.98 2.275 12.11 2.405 ;
 RECT 13.86 0.505 13.99 0.635 ;
 RECT 8.69 0.505 8.82 0.635 ;
 RECT 6.335 2.295 6.465 2.425 ;
 RECT 12.92 0.5 13.05 0.63 ;
 RECT 11.51 0.505 11.64 0.635 ;
 RECT 10.1 1.75 10.23 1.88 ;
 RECT 11.51 1.75 11.64 1.88 ;
 RECT 5.39 2.295 5.52 2.425 ;
 RECT 6.335 2.035 6.465 2.165 ;
 RECT 9.16 2.015 9.29 2.145 ;
 RECT 4.92 2.295 5.05 2.425 ;
 RECT 7.28 0.765 7.41 0.895 ;
 RECT 4.92 2.035 5.05 2.165 ;
 RECT 11.04 1.485 11.17 1.615 ;
 RECT 1.06 1.5 1.19 1.63 ;
 RECT 14.895 2.07 15.025 2.2 ;
 RECT 9.63 1.485 9.76 1.615 ;
 LAYER M1 ;
 RECT 1.895 0.53 2.035 1.985 ;
 RECT 3.605 0.365 3.745 0.925 ;
 RECT 3.605 1.065 3.745 1.205 ;
 RECT 3.605 1.345 3.745 1.775 ;
 RECT 2.82 1.205 3.745 1.345 ;
 RECT 3.56 1.775 3.79 1.915 ;
 RECT 3.605 0.925 4.28 1.065 ;
 RECT 6.33 1.725 6.47 2.355 ;
 RECT 5.385 1.725 5.525 2.355 ;
 RECT 5.385 2.355 6.47 2.495 ;
 RECT 2.365 0.455 2.505 0.925 ;
 RECT 2.365 1.065 2.505 1.775 ;
 RECT 2.32 1.775 2.55 1.915 ;
 RECT 2.365 0.925 3.465 1.065 ;
 RECT 5.86 1.025 6 1.125 ;
 RECT 5.86 1.265 6 2.215 ;
 RECT 6.335 0.525 6.475 1.125 ;
 RECT 5.395 0.885 6 1.025 ;
 RECT 5.395 0.35 5.535 0.885 ;
 RECT 5.86 1.125 7.29 1.265 ;
 RECT 4.445 0.48 4.585 1.36 ;
 RECT 4.145 1.5 4.585 1.505 ;
 RECT 4.145 1.505 4.285 1.68 ;
 RECT 4.445 1.36 5.365 1.365 ;
 RECT 4.145 1.365 5.365 1.5 ;
 RECT 5.225 1.185 5.72 1.325 ;
 RECT 5.225 1.325 5.365 1.36 ;
 RECT 1.055 2.205 3.445 2.27 ;
 RECT 2.455 2.095 2.685 2.13 ;
 RECT 2.455 2.27 2.685 2.305 ;
 RECT 1.055 0.225 1.35 0.365 ;
 RECT 1.055 0.365 1.195 2.13 ;
 RECT 1.055 0.22 1.195 0.225 ;
 RECT 4.595 2.205 4.735 2.655 ;
 RECT 1.055 2.13 4.735 2.205 ;
 RECT 3.305 2.065 4.735 2.13 ;
 RECT 0.115 0.725 0.255 2.24 ;
 RECT 0.115 2.24 0.345 2.45 ;
 END
END CGLNPSX16

MACRO CGLNPSX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8 BY 2.88 ;
 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 1.16 1.925 1.4 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.43 0.565 7.48 0.705 ;
 RECT 7.24 0.705 7.48 0.765 ;
 RECT 7.24 0.525 7.48 0.565 ;
 RECT 6.7 0.705 6.84 2.47 ;
 END
 ANTENNADIFFAREA 0.57 ;
 END GCLK

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.195 2.11 0.615 2.36 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.925 0.84 5.24 1.09 ;
 END
 ANTENNAGATEAREA 0.051 ;
 END SE

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8 2.96 ;
 RECT 1.55 2.625 1.78 2.8 ;
 RECT 3.305 2.345 3.445 2.8 ;
 RECT 7.17 1.45 7.31 2.8 ;
 RECT 5.085 1.61 5.225 2.8 ;
 RECT 6.23 1.715 6.37 2.8 ;
 RECT 0.755 1.495 0.895 2.8 ;
 RECT 7.65 2.25 7.79 2.8 ;
 RECT 7.665 1.5 7.805 2.065 ;
 RECT 7.65 2.065 7.805 2.25 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8 0.08 ;
 RECT 1.545 0.585 1.8 0.725 ;
 RECT 6.965 0.08 7.105 0.355 ;
 RECT 6.025 0.08 6.165 0.68 ;
 RECT 3.305 0.08 3.445 0.74 ;
 RECT 0.755 0.08 0.895 0.99 ;
 RECT 5.085 0.08 5.225 0.68 ;
 RECT 4.145 0.08 4.285 0.715 ;
 RECT 1.66 0.08 1.8 0.585 ;
 RECT 7.63 0.08 7.77 0.85 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 2.32 1.26 2.42 2.35 ;
 RECT 2.79 0.315 2.89 0.89 ;
 RECT 2.71 0.89 2.89 0.99 ;
 RECT 2.71 0.99 2.81 1.16 ;
 RECT 2.32 1.16 2.81 1.26 ;
 RECT 2.21 2.35 2.42 2.58 ;
 RECT 4.22 0.89 4.5 1 ;
 RECT 4.4 0.28 4.5 0.89 ;
 RECT 4.22 1 4.67 1.1 ;
 RECT 4.57 1.1 4.67 1.85 ;
 RECT 2.79 1.56 2.89 2.03 ;
 RECT 2.61 2.03 2.89 2.24 ;
 RECT 2.32 0.19 2.42 0.885 ;
 RECT 1.29 0.09 2.42 0.19 ;
 RECT 1.29 0.19 1.52 0.4 ;
 RECT 1.85 0.37 1.95 1.19 ;
 RECT 1.85 1.4 1.95 2.14 ;
 RECT 1.69 1.19 1.95 1.4 ;
 RECT 3.09 0.315 3.19 1.17 ;
 RECT 3.09 1.38 3.19 2.14 ;
 RECT 2.99 1.17 3.22 1.38 ;
 RECT 5.34 0.28 5.44 2.4 ;
 RECT 4.72 2.27 4.95 2.4 ;
 RECT 4.72 2.4 5.44 2.5 ;
 RECT 3.405 0.89 3.66 1.1 ;
 RECT 3.56 0.38 3.66 0.89 ;
 RECT 3.56 1.1 3.66 2.14 ;
 RECT 6.055 1.04 6.38 1.15 ;
 RECT 6.055 1.15 7.055 1.25 ;
 RECT 6.485 1.25 6.585 2.76 ;
 RECT 6.75 0.28 6.85 1.15 ;
 RECT 6.28 0.28 6.38 1.04 ;
 RECT 6.955 1.25 7.055 2.76 ;
 RECT 5.81 0.28 5.91 0.75 ;
 RECT 5.645 0.85 5.745 1.08 ;
 RECT 5.645 1.29 5.745 2.5 ;
 RECT 5.645 0.75 5.91 0.85 ;
 RECT 5.625 1.08 5.855 1.29 ;
 RECT 1.01 1.355 1.11 2.31 ;
 RECT 1.01 2.31 1.3 2.52 ;
 RECT 1.01 0.57 1.11 1.145 ;
 RECT 0.825 1.145 1.11 1.355 ;
 RECT 0.54 0.57 0.64 2.13 ;
 RECT 0.35 2.13 0.64 2.34 ;
 RECT 4.87 0.87 5.155 1.08 ;
 RECT 4.87 0.28 4.97 0.87 ;
 RECT 4.87 1.08 4.97 1.85 ;
 LAYER CO ;
 RECT 6.235 1.765 6.365 1.895 ;
 RECT 6.705 2.29 6.835 2.42 ;
 RECT 4.62 0.53 4.75 0.66 ;
 RECT 6.235 2.03 6.365 2.16 ;
 RECT 2.54 0.535 2.67 0.665 ;
 RECT 0.29 0.79 0.42 0.92 ;
 RECT 6.105 1.08 6.235 1.21 ;
 RECT 7.67 2.07 7.8 2.2 ;
 RECT 5.865 1.51 5.995 1.64 ;
 RECT 7.67 1.81 7.8 1.94 ;
 RECT 6.705 1.765 6.835 1.895 ;
 RECT 5.56 0.5 5.69 0.63 ;
 RECT 0.29 1.565 0.42 1.695 ;
 RECT 1.6 2.63 1.73 2.76 ;
 RECT 2.07 1.78 2.2 1.91 ;
 RECT 1.12 2.35 1.25 2.48 ;
 RECT 1.74 1.23 1.87 1.36 ;
 RECT 3.78 1.78 3.91 1.91 ;
 RECT 7.67 1.55 7.8 1.68 ;
 RECT 5.865 1.77 5.995 1.9 ;
 RECT 2.07 0.59 2.2 0.72 ;
 RECT 6.235 2.29 6.365 2.42 ;
 RECT 5.09 0.5 5.22 0.63 ;
 RECT 4.32 1.5 4.45 1.63 ;
 RECT 3.455 0.93 3.585 1.06 ;
 RECT 5.675 1.12 5.805 1.25 ;
 RECT 7.175 2.03 7.305 2.16 ;
 RECT 3.31 0.535 3.44 0.665 ;
 RECT 7.175 1.765 7.305 1.895 ;
 RECT 6.97 0.155 7.1 0.285 ;
 RECT 5.09 1.7 5.22 1.83 ;
 RECT 6.705 1.5 6.835 1.63 ;
 RECT 1.23 1.685 1.36 1.815 ;
 RECT 0.76 1.565 0.89 1.695 ;
 RECT 6.5 0.57 6.63 0.7 ;
 RECT 0.875 1.185 1.005 1.315 ;
 RECT 0.4 2.17 0.53 2.3 ;
 RECT 4.975 0.91 5.105 1.04 ;
 RECT 7.175 2.29 7.305 2.42 ;
 RECT 7.635 0.67 7.765 0.8 ;
 RECT 2.25 2.4 2.38 2.53 ;
 RECT 7.175 1.5 7.305 1.63 ;
 RECT 2.54 1.78 2.67 1.91 ;
 RECT 3.31 2.395 3.44 2.525 ;
 RECT 5.09 1.96 5.22 2.09 ;
 RECT 5.865 2.03 5.995 2.16 ;
 RECT 4.27 0.93 4.4 1.06 ;
 RECT 4.15 0.53 4.28 0.66 ;
 RECT 2.66 2.07 2.79 2.2 ;
 RECT 1.34 0.23 1.47 0.36 ;
 RECT 7.635 0.41 7.765 0.54 ;
 RECT 6.03 0.5 6.16 0.63 ;
 RECT 1.6 0.59 1.73 0.72 ;
 RECT 0.76 0.79 0.89 0.92 ;
 RECT 3.04 1.21 3.17 1.34 ;
 RECT 6.705 2.03 6.835 2.16 ;
 RECT 1.23 0.79 1.36 0.92 ;
 RECT 3.78 0.6 3.91 0.73 ;
 RECT 4.77 2.315 4.9 2.445 ;
 LAYER M1 ;
 RECT 5.555 0.45 5.695 0.82 ;
 RECT 5.86 1.54 6 2.21 ;
 RECT 5.995 0.96 6.135 1.075 ;
 RECT 5.995 1.215 6.135 1.4 ;
 RECT 5.555 0.82 6.135 0.96 ;
 RECT 5.86 1.4 6.135 1.54 ;
 RECT 5.995 1.075 6.285 1.215 ;
 RECT 4.59 0.525 4.755 0.71 ;
 RECT 4.615 0.48 4.755 0.525 ;
 RECT 4.59 0.71 4.73 1.24 ;
 RECT 4.315 1.38 4.455 1.685 ;
 RECT 4.315 1.255 5.72 1.38 ;
 RECT 4.315 1.24 5.855 1.255 ;
 RECT 5.58 1.115 5.855 1.24 ;
 RECT 2.065 0.53 2.205 1.775 ;
 RECT 2.02 1.775 2.25 1.915 ;
 RECT 2.535 1.065 2.675 1.775 ;
 RECT 2.535 0.455 2.675 0.925 ;
 RECT 2.49 1.775 2.72 1.915 ;
 RECT 2.535 0.925 3.635 1.065 ;
 RECT 2.245 2.485 2.385 2.58 ;
 RECT 1.06 2.345 2.385 2.485 ;
 RECT 3.775 0.365 3.915 0.925 ;
 RECT 3.775 1.065 3.915 1.205 ;
 RECT 3.775 1.345 3.915 1.775 ;
 RECT 2.99 1.205 3.915 1.345 ;
 RECT 3.73 1.775 3.96 1.915 ;
 RECT 3.775 0.925 4.45 1.065 ;
 RECT 1.225 0.22 1.365 0.225 ;
 RECT 1.225 0.365 1.365 0.74 ;
 RECT 1.195 1.005 1.335 1.635 ;
 RECT 1.225 1.865 1.365 2.065 ;
 RECT 1.195 0.74 1.405 1.005 ;
 RECT 1.19 1.635 1.41 1.865 ;
 RECT 1.225 0.225 1.52 0.365 ;
 RECT 4.765 2.205 4.905 2.5 ;
 RECT 1.225 2.065 4.905 2.205 ;
 RECT 0.285 0.6 0.425 1.18 ;
 RECT 0.285 1.32 0.425 1.765 ;
 RECT 0.825 1.145 1.055 1.18 ;
 RECT 0.825 1.32 1.055 1.355 ;
 RECT 0.285 1.18 1.055 1.32 ;
 END
END CGLNPSX2

MACRO CGLNPSX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.96 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.96 2.96 ;
 RECT 0.71 1.765 0.94 1.905 ;
 RECT 1.55 2.625 1.78 2.8 ;
 RECT 7.17 1.435 7.31 2.8 ;
 RECT 8.51 2.085 8.65 2.8 ;
 RECT 5.085 1.715 5.225 2.8 ;
 RECT 6.23 1.715 6.37 2.8 ;
 RECT 8.11 1.96 8.25 2.8 ;
 RECT 3.305 2.345 3.445 2.8 ;
 RECT 0.755 1.905 0.895 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.96 0.08 ;
 RECT 1.53 0.585 1.915 0.725 ;
 RECT 0.755 0.08 0.895 0.985 ;
 RECT 4.145 0.08 4.285 0.715 ;
 RECT 6.965 0.08 7.105 0.98 ;
 RECT 6.025 0.08 6.165 0.68 ;
 RECT 3.305 0.08 3.445 0.74 ;
 RECT 5.085 0.08 5.225 0.68 ;
 RECT 7.905 0.08 8.045 0.98 ;
 RECT 1.775 0.08 1.915 0.585 ;
 RECT 8.475 0.08 8.615 0.85 ;
 END
 END VSS

 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 1.16 1.92 1.405 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.89 0.825 5.32 1.1 ;
 END
 ANTENNAGATEAREA 0.051 ;
 END SE

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.7 1.265 6.84 2.47 ;
 RECT 6.495 0.45 6.635 1.125 ;
 RECT 8.2 1.62 8.44 1.72 ;
 RECT 7.64 1.62 7.78 2.49 ;
 RECT 7.64 1.48 8.44 1.62 ;
 RECT 7.64 1.27 7.78 1.48 ;
 RECT 7.435 1.265 7.78 1.27 ;
 RECT 7.435 0.445 7.575 1.125 ;
 RECT 6.495 1.125 7.78 1.265 ;
 END
 ANTENNADIFFAREA 1.2 ;
 END GCLK

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 2.12 0.595 2.36 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 OBS
 LAYER PO ;
 RECT 1.85 0.37 1.95 1.19 ;
 RECT 1.85 1.4 1.95 2.14 ;
 RECT 1.69 1.19 1.95 1.4 ;
 RECT 3.09 0.315 3.19 1.17 ;
 RECT 3.09 1.38 3.19 2.14 ;
 RECT 2.99 1.17 3.22 1.38 ;
 RECT 5.81 0.28 5.91 0.75 ;
 RECT 5.645 0.85 5.745 1.08 ;
 RECT 5.645 1.29 5.745 2.52 ;
 RECT 5.645 0.75 5.91 0.85 ;
 RECT 5.625 1.08 5.855 1.29 ;
 RECT 5.34 0.28 5.44 2.425 ;
 RECT 4.72 2.295 4.95 2.425 ;
 RECT 4.72 2.425 5.44 2.525 ;
 RECT 4.87 1.065 4.97 1.85 ;
 RECT 4.87 0.28 4.97 0.855 ;
 RECT 4.87 0.855 5.125 1.065 ;
 RECT 4.22 0.89 4.5 1.1 ;
 RECT 4.4 0.28 4.5 0.89 ;
 RECT 4.4 1.1 4.5 1.28 ;
 RECT 4.57 1.38 4.67 1.85 ;
 RECT 4.4 1.28 4.67 1.38 ;
 RECT 3.405 0.89 3.66 1.1 ;
 RECT 3.56 0.38 3.66 0.89 ;
 RECT 3.56 1.1 3.66 2.14 ;
 RECT 2.79 1.56 2.89 2.03 ;
 RECT 2.61 2.03 2.89 2.24 ;
 RECT 1.375 0.09 2.42 0.19 ;
 RECT 2.32 0.19 2.42 0.885 ;
 RECT 1.375 0.19 1.605 0.405 ;
 RECT 2.32 1.26 2.42 2.35 ;
 RECT 2.79 0.315 2.89 0.89 ;
 RECT 2.71 0.89 2.89 0.99 ;
 RECT 2.71 0.99 2.81 1.16 ;
 RECT 2.32 1.16 2.81 1.26 ;
 RECT 2.21 2.35 2.42 2.58 ;
 RECT 6.055 1.04 6.38 1.15 ;
 RECT 6.055 1.15 7.995 1.25 ;
 RECT 6.28 0.255 6.38 1.04 ;
 RECT 7.69 0.255 7.79 1.15 ;
 RECT 7.425 1.25 7.525 2.76 ;
 RECT 7.22 0.255 7.32 1.15 ;
 RECT 6.955 1.25 7.055 2.76 ;
 RECT 6.75 0.255 6.85 1.15 ;
 RECT 6.485 1.25 6.585 2.76 ;
 RECT 7.895 1.25 7.995 2.76 ;
 RECT 0.82 1.2 1.11 1.41 ;
 RECT 1.01 1.41 1.11 2.31 ;
 RECT 1.01 2.31 1.265 2.52 ;
 RECT 1.01 0.56 1.11 1.2 ;
 RECT 0.54 0.57 0.64 2.12 ;
 RECT 0.355 2.12 0.64 2.33 ;
 LAYER CO ;
 RECT 4.32 1.5 4.45 1.63 ;
 RECT 6.105 1.08 6.235 1.21 ;
 RECT 4.77 2.34 4.9 2.47 ;
 RECT 4.27 0.93 4.4 1.06 ;
 RECT 5.56 0.5 5.69 0.63 ;
 RECT 4.945 0.895 5.075 1.025 ;
 RECT 8.48 0.67 8.61 0.8 ;
 RECT 3.455 0.93 3.585 1.06 ;
 RECT 8.515 2.395 8.645 2.525 ;
 RECT 8.48 0.41 8.61 0.54 ;
 RECT 8.515 2.135 8.645 2.265 ;
 RECT 2.25 2.4 2.38 2.53 ;
 RECT 1.23 0.79 1.36 0.92 ;
 RECT 5.09 1.765 5.22 1.895 ;
 RECT 6.705 1.765 6.835 1.895 ;
 RECT 3.78 1.78 3.91 1.91 ;
 RECT 0.29 1.77 0.42 1.9 ;
 RECT 3.78 0.6 3.91 0.73 ;
 RECT 6.705 2.03 6.835 2.16 ;
 RECT 1.23 1.77 1.36 1.9 ;
 RECT 6.705 2.29 6.835 2.42 ;
 RECT 3.04 1.21 3.17 1.34 ;
 RECT 2.07 0.59 2.2 0.72 ;
 RECT 7.175 2.03 7.305 2.16 ;
 RECT 5.865 1.77 5.995 1.9 ;
 RECT 6.705 1.5 6.835 1.63 ;
 RECT 3.31 2.395 3.44 2.525 ;
 RECT 3.31 0.535 3.44 0.665 ;
 RECT 6.97 0.765 7.1 0.895 ;
 RECT 1.6 0.59 1.73 0.72 ;
 RECT 0.76 0.79 0.89 0.92 ;
 RECT 0.87 1.24 1 1.37 ;
 RECT 0.405 2.16 0.535 2.29 ;
 RECT 6.03 0.5 6.16 0.63 ;
 RECT 6.97 0.505 7.1 0.635 ;
 RECT 5.675 1.12 5.805 1.25 ;
 RECT 5.09 2.025 5.22 2.155 ;
 RECT 2.54 1.78 2.67 1.91 ;
 RECT 6.235 2.03 6.365 2.16 ;
 RECT 6.235 1.765 6.365 1.895 ;
 RECT 2.07 1.78 2.2 1.91 ;
 RECT 4.15 0.53 4.28 0.66 ;
 RECT 1.6 2.63 1.73 2.76 ;
 RECT 7.175 1.765 7.305 1.895 ;
 RECT 1.74 1.23 1.87 1.36 ;
 RECT 0.29 0.79 0.42 0.92 ;
 RECT 1.085 2.35 1.215 2.48 ;
 RECT 5.865 1.51 5.995 1.64 ;
 RECT 0.76 1.77 0.89 1.9 ;
 RECT 5.09 0.5 5.22 0.63 ;
 RECT 7.91 0.765 8.04 0.895 ;
 RECT 7.91 0.505 8.04 0.635 ;
 RECT 7.44 0.765 7.57 0.895 ;
 RECT 7.44 0.505 7.57 0.635 ;
 RECT 8.115 2.29 8.245 2.42 ;
 RECT 8.115 2.03 8.245 2.16 ;
 RECT 7.645 2.03 7.775 2.16 ;
 RECT 7.645 1.5 7.775 1.63 ;
 RECT 7.645 1.765 7.775 1.895 ;
 RECT 7.645 2.29 7.775 2.42 ;
 RECT 2.66 2.07 2.79 2.2 ;
 RECT 7.175 1.5 7.305 1.63 ;
 RECT 5.865 2.03 5.995 2.16 ;
 RECT 4.62 0.53 4.75 0.66 ;
 RECT 6.5 0.5 6.63 0.63 ;
 RECT 7.175 2.29 7.305 2.42 ;
 RECT 6.5 0.765 6.63 0.895 ;
 RECT 2.54 0.535 2.67 0.665 ;
 RECT 1.425 0.235 1.555 0.365 ;
 RECT 6.235 2.29 6.365 2.42 ;
 LAYER M1 ;
 RECT 5.555 0.45 5.695 0.82 ;
 RECT 5.86 1.54 6 2.21 ;
 RECT 5.995 0.96 6.135 1.075 ;
 RECT 5.995 1.215 6.135 1.4 ;
 RECT 5.555 0.82 6.135 0.96 ;
 RECT 5.86 1.4 6.135 1.54 ;
 RECT 5.995 1.075 6.285 1.215 ;
 RECT 4.61 0.665 4.75 1.24 ;
 RECT 4.61 1.38 4.75 1.425 ;
 RECT 4.315 1.565 4.455 1.685 ;
 RECT 4.315 1.425 4.75 1.565 ;
 RECT 4.57 0.525 4.8 0.665 ;
 RECT 4.61 1.24 5.855 1.255 ;
 RECT 4.61 1.255 5.72 1.38 ;
 RECT 5.58 1.115 5.855 1.24 ;
 RECT 1.035 2.345 2.385 2.485 ;
 RECT 2.245 2.485 2.385 2.58 ;
 RECT 2.535 1.065 2.675 1.775 ;
 RECT 2.535 0.455 2.675 0.925 ;
 RECT 2.49 1.775 2.72 1.915 ;
 RECT 2.535 0.925 3.635 1.065 ;
 RECT 3.775 1.065 3.915 1.205 ;
 RECT 3.775 1.345 3.915 1.775 ;
 RECT 2.99 1.205 3.915 1.345 ;
 RECT 3.775 0.365 3.915 0.925 ;
 RECT 3.73 1.775 3.96 1.915 ;
 RECT 3.775 0.925 4.45 1.065 ;
 RECT 2.065 0.53 2.205 1.775 ;
 RECT 2.02 1.775 2.25 1.915 ;
 RECT 1.225 0.37 1.365 0.74 ;
 RECT 1.19 0.99 1.33 1.565 ;
 RECT 1.225 1.705 1.365 2.065 ;
 RECT 1.185 1.565 1.365 1.705 ;
 RECT 1.17 0.74 1.385 0.99 ;
 RECT 1.225 0.23 1.605 0.37 ;
 RECT 4.765 2.205 4.905 2.525 ;
 RECT 1.225 2.065 4.905 2.205 ;
 RECT 0.285 0.62 0.425 1.235 ;
 RECT 0.285 1.375 0.425 1.97 ;
 RECT 0.82 1.2 1.05 1.235 ;
 RECT 0.82 1.375 1.05 1.41 ;
 RECT 0.285 1.235 1.05 1.375 ;
 END
END CGLNPSX4

MACRO CGLNPSX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.88 BY 2.88 ;
 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.425 1.16 0.76 1.495 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.985 1.8 4.35 2.14 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END SE

 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 0.84 1.75 1.15 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.88 0.08 ;
 RECT 1.36 0.52 1.63 0.66 ;
 RECT 0.585 0.08 0.725 0.985 ;
 RECT 3.975 0.08 4.115 0.68 ;
 RECT 8.675 0.08 8.815 0.98 ;
 RECT 9.615 0.08 9.755 0.98 ;
 RECT 4.915 0.08 5.055 0.68 ;
 RECT 3.135 0.08 3.275 0.74 ;
 RECT 7.735 0.08 7.875 0.98 ;
 RECT 5.855 0.08 5.995 0.68 ;
 RECT 6.795 0.08 6.935 0.98 ;
 RECT 10.185 0.08 10.325 0.85 ;
 RECT 1.49 0.08 1.63 0.52 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.88 2.96 ;
 RECT 0.54 1.765 0.77 1.905 ;
 RECT 1.38 2.625 1.61 2.8 ;
 RECT 7 1.45 7.14 2.8 ;
 RECT 4.915 1.52 5.055 2.8 ;
 RECT 7.94 1.45 8.08 2.8 ;
 RECT 8.88 1.45 9.02 2.8 ;
 RECT 9.82 1.45 9.96 2.8 ;
 RECT 3.135 2.35 3.275 2.8 ;
 RECT 6.06 1.715 6.2 2.8 ;
 RECT 10.205 2.25 10.345 2.8 ;
 RECT 10.22 1.5 10.36 2.065 ;
 RECT 10.205 2.065 10.36 2.25 ;
 RECT 0.585 1.905 0.725 2.8 ;
 END
 END VDD

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.53 1.46 6.86 1.74 ;
 RECT 6.325 0.45 6.465 1.125 ;
 RECT 7.47 1.27 7.61 2.49 ;
 RECT 8.205 0.45 8.345 1.13 ;
 RECT 8.41 1.27 8.55 2.47 ;
 RECT 9.145 0.445 9.285 1.13 ;
 RECT 9.35 1.27 9.49 2.49 ;
 RECT 6.53 1.74 6.67 2.47 ;
 RECT 6.53 1.265 6.67 1.46 ;
 RECT 7.265 0.445 7.405 1.125 ;
 RECT 6.325 1.125 7.405 1.13 ;
 RECT 7.265 1.265 9.49 1.27 ;
 RECT 6.325 1.13 9.49 1.265 ;
 END
 ANTENNADIFFAREA 2.488 ;
 END GCLK

 OBS
 LAYER PO ;
 RECT 3.39 1.1 3.49 2.14 ;
 RECT 3.39 0.38 3.49 0.89 ;
 RECT 3.235 0.89 3.49 1.1 ;
 RECT 5.64 0.28 5.74 0.75 ;
 RECT 5.475 1.29 5.575 2.54 ;
 RECT 5.475 0.85 5.575 1.08 ;
 RECT 5.475 0.75 5.74 0.85 ;
 RECT 5.455 1.08 5.685 1.29 ;
 RECT 5.17 0.28 5.27 2.445 ;
 RECT 4.545 2.43 4.775 2.445 ;
 RECT 4.545 2.545 4.775 2.66 ;
 RECT 4.545 2.445 5.27 2.545 ;
 RECT 2.62 1.56 2.72 2.03 ;
 RECT 2.44 2.03 2.72 2.24 ;
 RECT 1.68 1.08 1.78 2.14 ;
 RECT 1.68 0.37 1.78 0.87 ;
 RECT 1.52 0.87 1.78 1.08 ;
 RECT 5.885 1.15 9.705 1.25 ;
 RECT 5.885 1.04 6.21 1.15 ;
 RECT 7.05 0.195 7.15 1.15 ;
 RECT 7.52 0.195 7.62 1.15 ;
 RECT 6.58 0.195 6.68 1.15 ;
 RECT 7.255 1.25 7.355 2.76 ;
 RECT 6.315 1.25 6.415 2.76 ;
 RECT 6.785 1.25 6.885 2.76 ;
 RECT 9.135 1.25 9.235 2.76 ;
 RECT 8.46 0.195 8.56 1.15 ;
 RECT 9.4 0.195 9.5 1.15 ;
 RECT 8.665 1.25 8.765 2.76 ;
 RECT 8.195 1.25 8.295 2.76 ;
 RECT 8.93 0.195 9.03 1.15 ;
 RECT 6.11 0.195 6.21 1.04 ;
 RECT 9.605 1.25 9.705 2.76 ;
 RECT 7.99 0.195 8.09 1.15 ;
 RECT 7.725 1.25 7.825 2.76 ;
 RECT 4.05 1.28 4.5 1.38 ;
 RECT 4.05 1.095 4.33 1.28 ;
 RECT 4.23 0.28 4.33 1.095 ;
 RECT 4.4 1.38 4.5 1.85 ;
 RECT 2.15 0.19 2.25 0.885 ;
 RECT 1.12 0.09 2.25 0.19 ;
 RECT 1.12 0.19 1.35 0.4 ;
 RECT 2.92 0.315 3.02 1.17 ;
 RECT 2.92 1.38 3.02 2.14 ;
 RECT 2.82 1.17 3.05 1.38 ;
 RECT 2.15 1.26 2.25 2.35 ;
 RECT 2.62 0.315 2.72 0.89 ;
 RECT 2.54 0.89 2.72 0.99 ;
 RECT 2.54 0.99 2.64 1.16 ;
 RECT 2.15 1.16 2.64 1.26 ;
 RECT 2.04 2.35 2.25 2.58 ;
 RECT 4.7 0.28 4.8 2.035 ;
 RECT 3.985 1.93 4.215 2.035 ;
 RECT 3.985 2.135 4.215 2.14 ;
 RECT 3.985 2.035 4.8 2.135 ;
 RECT 0.84 0.565 0.94 2.31 ;
 RECT 0.84 2.31 1.11 2.36 ;
 RECT 0.115 2.36 1.11 2.46 ;
 RECT 0.84 2.46 1.11 2.52 ;
 RECT 0.115 2.315 0.345 2.36 ;
 RECT 0.115 2.46 0.345 2.525 ;
 RECT 0.37 1.285 0.66 1.495 ;
 RECT 0.37 0.57 0.47 1.285 ;
 RECT 0.37 1.495 0.47 2.12 ;
 LAYER CO ;
 RECT 9.355 2.29 9.485 2.42 ;
 RECT 8.68 0.765 8.81 0.895 ;
 RECT 9.62 0.765 9.75 0.895 ;
 RECT 8.415 2.03 8.545 2.16 ;
 RECT 9.825 2.03 9.955 2.16 ;
 RECT 6.33 0.765 6.46 0.895 ;
 RECT 4.15 1.5 4.28 1.63 ;
 RECT 4.92 2.09 5.05 2.22 ;
 RECT 5.695 1.77 5.825 1.9 ;
 RECT 2.08 2.4 2.21 2.53 ;
 RECT 3.285 0.93 3.415 1.06 ;
 RECT 5.935 1.08 6.065 1.21 ;
 RECT 2.49 2.07 2.62 2.2 ;
 RECT 1.06 0.79 1.19 0.92 ;
 RECT 0.93 2.35 1.06 2.48 ;
 RECT 1.06 1.77 1.19 1.9 ;
 RECT 4.45 0.5 4.58 0.63 ;
 RECT 1.43 2.63 1.56 2.76 ;
 RECT 3.61 1.78 3.74 1.91 ;
 RECT 6.33 0.5 6.46 0.63 ;
 RECT 5.39 0.5 5.52 0.63 ;
 RECT 1.9 1.78 2.03 1.91 ;
 RECT 3.14 0.535 3.27 0.665 ;
 RECT 3.14 2.4 3.27 2.53 ;
 RECT 4.595 2.475 4.725 2.605 ;
 RECT 4.035 1.97 4.165 2.1 ;
 RECT 0.165 2.355 0.295 2.485 ;
 RECT 0.48 1.325 0.61 1.455 ;
 RECT 7.475 1.765 7.605 1.895 ;
 RECT 5.695 1.51 5.825 1.64 ;
 RECT 7.005 2.03 7.135 2.16 ;
 RECT 2.37 1.78 2.5 1.91 ;
 RECT 7.27 0.765 7.4 0.895 ;
 RECT 10.225 1.55 10.355 1.68 ;
 RECT 6.8 0.505 6.93 0.635 ;
 RECT 7.475 2.29 7.605 2.42 ;
 RECT 5.86 0.5 5.99 0.63 ;
 RECT 6.065 2.03 6.195 2.16 ;
 RECT 2.87 1.21 3 1.34 ;
 RECT 6.065 1.765 6.195 1.895 ;
 RECT 0.12 1.77 0.25 1.9 ;
 RECT 6.065 2.29 6.195 2.42 ;
 RECT 7.74 0.505 7.87 0.635 ;
 RECT 1.57 0.91 1.7 1.04 ;
 RECT 7.945 2.29 8.075 2.42 ;
 RECT 3.98 0.5 4.11 0.63 ;
 RECT 0.12 0.79 0.25 0.92 ;
 RECT 4.92 1.83 5.05 1.96 ;
 RECT 1.9 0.59 2.03 0.72 ;
 RECT 2.37 0.535 2.5 0.665 ;
 RECT 5.505 1.12 5.635 1.25 ;
 RECT 8.415 2.29 8.545 2.42 ;
 RECT 8.415 1.5 8.545 1.63 ;
 RECT 8.885 1.765 9.015 1.895 ;
 RECT 9.355 1.765 9.485 1.895 ;
 RECT 9.825 1.765 9.955 1.895 ;
 RECT 8.21 0.5 8.34 0.63 ;
 RECT 8.885 1.5 9.015 1.63 ;
 RECT 9.355 2.03 9.485 2.16 ;
 RECT 9.355 1.5 9.485 1.63 ;
 RECT 9.15 0.765 9.28 0.895 ;
 RECT 9.62 0.505 9.75 0.635 ;
 RECT 8.885 2.29 9.015 2.42 ;
 RECT 8.21 0.765 8.34 0.895 ;
 RECT 8.415 1.765 8.545 1.895 ;
 RECT 7.74 0.765 7.87 0.895 ;
 RECT 8.68 0.505 8.81 0.635 ;
 RECT 9.825 1.5 9.955 1.63 ;
 RECT 4.92 0.5 5.05 0.63 ;
 RECT 6.535 2.29 6.665 2.42 ;
 RECT 7.27 0.505 7.4 0.635 ;
 RECT 7.005 1.5 7.135 1.63 ;
 RECT 10.225 1.81 10.355 1.94 ;
 RECT 10.225 2.07 10.355 2.2 ;
 RECT 6.535 2.03 6.665 2.16 ;
 RECT 7.945 1.765 8.075 1.895 ;
 RECT 10.19 0.67 10.32 0.8 ;
 RECT 7.475 2.03 7.605 2.16 ;
 RECT 7.005 2.29 7.135 2.42 ;
 RECT 4.1 1.135 4.23 1.265 ;
 RECT 4.92 1.57 5.05 1.7 ;
 RECT 7.945 2.03 8.075 2.16 ;
 RECT 6.535 1.5 6.665 1.63 ;
 RECT 10.19 0.41 10.32 0.54 ;
 RECT 7.475 1.5 7.605 1.63 ;
 RECT 1.17 0.23 1.3 0.36 ;
 RECT 3.61 0.6 3.74 0.73 ;
 RECT 0.59 0.79 0.72 0.92 ;
 RECT 6.8 0.765 6.93 0.895 ;
 RECT 7.005 1.765 7.135 1.895 ;
 RECT 5.695 2.03 5.825 2.16 ;
 RECT 1.43 0.525 1.56 0.655 ;
 RECT 0.59 1.77 0.72 1.9 ;
 RECT 6.535 1.765 6.665 1.895 ;
 RECT 7.945 1.5 8.075 1.63 ;
 RECT 9.15 0.505 9.28 0.635 ;
 RECT 9.825 2.29 9.955 2.42 ;
 RECT 8.885 2.03 9.015 2.16 ;
 LAYER M1 ;
 RECT 1.895 0.53 2.035 1.775 ;
 RECT 1.85 1.775 2.08 1.915 ;
 RECT 2.075 2.485 2.215 2.58 ;
 RECT 0.88 2.345 2.215 2.485 ;
 RECT 5.385 0.45 5.525 0.82 ;
 RECT 5.69 1.54 5.83 2.21 ;
 RECT 5.825 0.96 5.965 1.075 ;
 RECT 5.825 1.215 5.965 1.4 ;
 RECT 5.385 0.82 5.965 0.96 ;
 RECT 5.69 1.4 5.965 1.54 ;
 RECT 5.825 1.075 6.115 1.215 ;
 RECT 2.365 0.455 2.505 0.925 ;
 RECT 2.365 1.065 2.505 1.775 ;
 RECT 2.32 1.775 2.55 1.915 ;
 RECT 2.365 0.925 3.465 1.065 ;
 RECT 3.605 1.345 3.745 1.775 ;
 RECT 2.82 1.27 3.745 1.345 ;
 RECT 3.605 0.365 3.745 1.13 ;
 RECT 3.56 1.775 3.79 1.915 ;
 RECT 2.82 1.205 4.285 1.27 ;
 RECT 3.605 1.13 4.285 1.205 ;
 RECT 4.445 0.45 4.585 1.24 ;
 RECT 4.445 1.38 4.585 1.495 ;
 RECT 4.08 1.495 4.585 1.635 ;
 RECT 5.41 1.115 5.685 1.24 ;
 RECT 4.445 1.24 5.685 1.255 ;
 RECT 4.445 1.255 5.55 1.38 ;
 RECT 1.055 0.365 1.195 2.065 ;
 RECT 1.055 0.225 1.35 0.365 ;
 RECT 1.055 2.065 3.555 2.205 ;
 RECT 3.415 2.205 3.555 2.52 ;
 RECT 3.415 2.52 4.73 2.66 ;
 RECT 4.59 2.425 4.73 2.52 ;
 RECT 0.115 0.71 0.255 2.315 ;
 RECT 0.115 2.315 0.345 2.525 ;
 END
END CGLNPSX8

MACRO CGLPPRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.36 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 1.43 1.95 1.735 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END SE

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.36 2.96 ;
 RECT 4.57 1.505 4.8 1.645 ;
 RECT 1.72 2.625 1.95 2.8 ;
 RECT 6.495 1.675 6.635 2.8 ;
 RECT 0.755 1.655 0.895 2.8 ;
 RECT 3.775 1.73 3.915 2.8 ;
 RECT 5.555 1.43 5.695 2.8 ;
 RECT 6.895 1.5 7.035 2.8 ;
 RECT 4.615 1.645 4.755 2.8 ;
 END
 END VDD

 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.1 1.145 2.37 1.425 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 2.12 0.615 2.36 ;
 END
 ANTENNAGATEAREA 0.063 ;
 END CLK

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.36 0.08 ;
 RECT 2.02 0.585 2.25 0.725 ;
 RECT 6.495 0.08 6.635 0.98 ;
 RECT 0.755 0.08 0.895 0.985 ;
 RECT 5.555 0.08 5.695 0.68 ;
 RECT 3.775 0.08 3.915 0.74 ;
 RECT 6.895 0.08 7.035 0.85 ;
 RECT 2.065 0.08 2.205 0.585 ;
 END
 END VSS

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.96 1.775 6.25 2.045 ;
 RECT 6.025 2.045 6.165 2.45 ;
 RECT 6.025 0.48 6.165 1.775 ;
 END
 ANTENNADIFFAREA 0.61 ;
 END GCLK

 OBS
 LAYER PO ;
 RECT 3.56 1.38 3.66 2.135 ;
 RECT 3.56 0.315 3.66 1.17 ;
 RECT 3.46 1.17 3.69 1.38 ;
 RECT 2.32 0.37 2.42 1.15 ;
 RECT 2.32 1.36 2.42 2.14 ;
 RECT 2.14 1.15 2.42 1.36 ;
 RECT 5.34 0.28 5.44 2.45 ;
 RECT 3.395 2.32 3.605 2.45 ;
 RECT 3.395 2.45 5.44 2.55 ;
 RECT 5.04 0.28 5.14 0.75 ;
 RECT 4.87 1.345 4.97 1.86 ;
 RECT 4.87 0.85 4.97 1.115 ;
 RECT 4.69 1.115 4.97 1.345 ;
 RECT 4.87 0.75 5.14 0.85 ;
 RECT 3.875 0.89 4.13 1.1 ;
 RECT 4.03 0.38 4.13 0.89 ;
 RECT 4.03 1.1 4.13 2.14 ;
 RECT 3.115 2.13 3.215 2.42 ;
 RECT 3.26 1.56 3.36 2.03 ;
 RECT 3.115 2.03 3.36 2.13 ;
 RECT 3.005 2.42 3.215 2.65 ;
 RECT 6.28 0.25 6.38 1.255 ;
 RECT 5.81 0.25 5.91 1.03 ;
 RECT 6.28 1.355 6.38 2.74 ;
 RECT 5.81 1.355 5.91 2.74 ;
 RECT 5.68 1.255 6.38 1.26 ;
 RECT 5.68 1.03 5.91 1.255 ;
 RECT 5.81 1.26 6.38 1.355 ;
 RECT 3.26 0.315 3.36 0.89 ;
 RECT 2.79 1.26 2.89 2.03 ;
 RECT 3.18 0.89 3.36 0.99 ;
 RECT 3.18 0.99 3.28 1.16 ;
 RECT 2.79 1.16 3.28 1.26 ;
 RECT 2.705 2.03 2.935 2.24 ;
 RECT 0.82 1.13 1.11 1.34 ;
 RECT 1.01 0.19 1.11 1.13 ;
 RECT 1.01 1.34 1.11 2.31 ;
 RECT 2.79 0.19 2.89 0.885 ;
 RECT 1.01 2.31 1.29 2.52 ;
 RECT 1.01 0.09 2.89 0.19 ;
 RECT 1.85 0.37 1.95 1.43 ;
 RECT 2.02 1.64 2.12 2.14 ;
 RECT 1.72 1.43 1.95 1.54 ;
 RECT 1.72 1.54 2.12 1.64 ;
 RECT 0.54 0.57 0.64 2.12 ;
 RECT 0.38 2.12 0.64 2.33 ;
 LAYER CO ;
 RECT 3.78 0.535 3.91 0.665 ;
 RECT 4.25 0.6 4.38 0.73 ;
 RECT 3.51 1.21 3.64 1.34 ;
 RECT 1.6 0.59 1.73 0.72 ;
 RECT 0.29 1.585 0.42 1.715 ;
 RECT 1.23 0.79 1.36 0.92 ;
 RECT 2.19 1.19 2.32 1.32 ;
 RECT 6.5 2.01 6.63 2.14 ;
 RECT 4.79 0.5 4.92 0.63 ;
 RECT 1.77 2.63 1.9 2.76 ;
 RECT 6.5 0.53 6.63 0.66 ;
 RECT 6.5 0.79 6.63 0.92 ;
 RECT 6.03 0.79 6.16 0.92 ;
 RECT 6.03 1.745 6.16 1.875 ;
 RECT 0.29 0.79 0.42 0.92 ;
 RECT 6.5 1.745 6.63 1.875 ;
 RECT 3.435 2.37 3.565 2.5 ;
 RECT 5.56 0.5 5.69 0.63 ;
 RECT 4.25 1.78 4.38 1.91 ;
 RECT 5.56 1.745 5.69 1.875 ;
 RECT 2.755 2.07 2.885 2.2 ;
 RECT 3.925 0.93 4.055 1.06 ;
 RECT 6.03 0.53 6.16 0.66 ;
 RECT 6.9 1.81 7.03 1.94 ;
 RECT 6.03 2.27 6.16 2.4 ;
 RECT 6.9 1.55 7.03 1.68 ;
 RECT 6.5 2.27 6.63 2.4 ;
 RECT 2.54 1.78 2.67 1.91 ;
 RECT 5.73 1.08 5.86 1.21 ;
 RECT 5.56 1.48 5.69 1.61 ;
 RECT 6.03 2.01 6.16 2.14 ;
 RECT 5.56 2.27 5.69 2.4 ;
 RECT 6.03 1.48 6.16 1.61 ;
 RECT 6.9 0.67 7.03 0.8 ;
 RECT 5.56 2.01 5.69 2.14 ;
 RECT 6.9 2.07 7.03 2.2 ;
 RECT 3.045 2.47 3.175 2.6 ;
 RECT 4.74 1.165 4.87 1.295 ;
 RECT 3.78 1.78 3.91 1.91 ;
 RECT 0.76 1.705 0.89 1.835 ;
 RECT 6.9 0.41 7.03 0.54 ;
 RECT 5.09 1.48 5.22 1.61 ;
 RECT 1.225 1.885 1.355 2.015 ;
 RECT 1.11 2.35 1.24 2.48 ;
 RECT 4.62 1.51 4.75 1.64 ;
 RECT 0.87 1.17 1 1.3 ;
 RECT 1.77 1.47 1.9 1.6 ;
 RECT 0.43 2.16 0.56 2.29 ;
 RECT 0.76 0.79 0.89 0.92 ;
 RECT 3.01 1.78 3.14 1.91 ;
 RECT 2.07 0.59 2.2 0.72 ;
 RECT 3.01 0.535 3.14 0.665 ;
 RECT 2.54 0.59 2.67 0.72 ;
 LAYER M1 ;
 RECT 5.085 0.975 5.225 1.08 ;
 RECT 5.085 1.22 5.225 1.66 ;
 RECT 4.785 0.45 4.925 0.835 ;
 RECT 4.785 0.835 5.225 0.975 ;
 RECT 5.725 1.03 5.865 1.08 ;
 RECT 5.725 1.22 5.865 1.26 ;
 RECT 5.085 1.08 5.865 1.22 ;
 RECT 1.595 0.53 1.735 0.865 ;
 RECT 2.535 1.005 2.675 1.775 ;
 RECT 2.535 0.53 2.675 0.865 ;
 RECT 1.595 0.865 2.675 1.005 ;
 RECT 2.49 1.775 2.72 1.915 ;
 RECT 4.245 0.365 4.385 1.205 ;
 RECT 4.245 1.345 4.385 1.96 ;
 RECT 4.735 1.115 4.875 1.205 ;
 RECT 3.46 1.205 4.875 1.345 ;
 RECT 3.005 0.455 3.145 0.925 ;
 RECT 3.005 1.065 3.145 1.775 ;
 RECT 2.96 1.775 3.19 1.915 ;
 RECT 3.005 0.925 4.105 1.065 ;
 RECT 3.04 2.485 3.18 2.65 ;
 RECT 1.06 2.345 3.18 2.485 ;
 RECT 1.19 1.13 1.33 1.88 ;
 RECT 1.19 0.99 1.365 1.13 ;
 RECT 1.225 0.715 1.365 0.99 ;
 RECT 1.09 1.88 1.43 2.065 ;
 RECT 1.09 2.065 3.57 2.205 ;
 RECT 3.43 2.205 3.57 2.55 ;
 RECT 0.285 0.57 0.425 1.165 ;
 RECT 0.285 1.305 0.425 1.79 ;
 RECT 0.82 1.13 1.05 1.165 ;
 RECT 0.82 1.305 1.05 1.34 ;
 RECT 0.285 1.165 1.05 1.305 ;
 END
END CGLPPRX2

MACRO CGLPPRX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.24 BY 2.88 ;
 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.085 1.145 2.395 1.435 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.24 2.96 ;
 RECT 1.72 2.62 1.95 2.8 ;
 RECT 7.435 1.425 7.575 2.8 ;
 RECT 8.375 1.425 8.515 2.8 ;
 RECT 5.555 1.425 5.695 2.8 ;
 RECT 0.755 1.58 0.895 2.8 ;
 RECT 4.515 2.34 4.655 2.8 ;
 RECT 3.725 2.34 3.865 2.8 ;
 RECT 9.315 1.425 9.455 2.8 ;
 RECT 6.495 1.425 6.635 2.8 ;
 RECT 9.715 1.495 9.855 2.8 ;
 END
 END VDD

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 1.42 1.945 1.72 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END SE

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 2.12 0.61 2.36 ;
 END
 ANTENNAGATEAREA 0.046 ;
 END CLK

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.24 0.08 ;
 RECT 2.02 0.585 2.25 0.725 ;
 RECT 5.555 0.08 5.695 0.685 ;
 RECT 7.435 0.08 7.575 0.97 ;
 RECT 8.375 0.08 8.515 0.97 ;
 RECT 9.315 0.08 9.455 0.97 ;
 RECT 0.755 0.08 0.895 0.97 ;
 RECT 3.775 0.08 3.915 0.735 ;
 RECT 6.495 0.08 6.635 0.97 ;
 RECT 9.715 0.08 9.855 0.845 ;
 RECT 2.065 0.08 2.205 0.585 ;
 END
 END VSS

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.775 1.76 9.105 2.06 ;
 RECT 8.845 2.06 8.985 2.545 ;
 RECT 6.025 1.115 8.985 1.255 ;
 RECT 8.845 1.255 8.985 1.76 ;
 RECT 8.845 0.47 8.985 1.115 ;
 RECT 6.025 1.255 6.165 2.53 ;
 RECT 6.025 0.47 6.165 1.115 ;
 RECT 6.965 1.255 7.105 2.525 ;
 RECT 6.965 0.47 7.105 1.115 ;
 RECT 7.905 1.255 8.045 2.55 ;
 RECT 7.905 0.47 8.045 1.115 ;
 END
 ANTENNADIFFAREA 2.4 ;
 END GCLK

 OBS
 LAYER PO ;
 RECT 3.875 0.885 4.13 1.095 ;
 RECT 4.03 0.375 4.13 0.885 ;
 RECT 4.03 1.095 4.13 2.135 ;
 RECT 3.26 0.31 3.36 0.885 ;
 RECT 2.79 1.255 2.89 2.025 ;
 RECT 3.18 0.885 3.36 0.985 ;
 RECT 3.18 0.985 3.28 1.155 ;
 RECT 2.79 1.155 3.28 1.255 ;
 RECT 2.705 2.025 2.935 2.235 ;
 RECT 3.56 1.375 3.66 2.135 ;
 RECT 3.56 0.31 3.66 1.165 ;
 RECT 3.46 1.165 3.69 1.375 ;
 RECT 5.34 0.09 5.44 2.425 ;
 RECT 5.18 2.425 5.44 2.59 ;
 RECT 5.18 2.59 5.41 2.635 ;
 RECT 3.26 1.555 3.36 2.345 ;
 RECT 3.15 2.345 3.36 2.575 ;
 RECT 2.32 0.37 2.42 1.14 ;
 RECT 2.32 1.35 2.42 2.135 ;
 RECT 2.135 1.14 2.42 1.35 ;
 RECT 5.645 1.075 5.91 1.145 ;
 RECT 5.81 0.27 5.91 1.075 ;
 RECT 9.1 0.27 9.2 1.145 ;
 RECT 9.1 1.245 9.2 2.775 ;
 RECT 6.28 0.27 6.38 1.145 ;
 RECT 6.28 1.245 6.38 2.775 ;
 RECT 6.75 0.27 6.85 1.145 ;
 RECT 6.75 1.245 6.85 2.775 ;
 RECT 8.63 0.27 8.73 1.145 ;
 RECT 8.63 1.245 8.73 2.775 ;
 RECT 8.16 0.27 8.26 1.145 ;
 RECT 8.16 1.245 8.26 2.775 ;
 RECT 7.69 0.27 7.79 1.145 ;
 RECT 7.69 1.245 7.79 2.775 ;
 RECT 5.645 1.245 5.91 1.285 ;
 RECT 5.81 1.285 5.91 2.775 ;
 RECT 7.22 0.27 7.32 1.145 ;
 RECT 7.22 1.245 7.32 2.775 ;
 RECT 5.645 1.145 9.2 1.245 ;
 RECT 5.04 0.09 5.14 1.11 ;
 RECT 4.87 1.34 4.97 2.54 ;
 RECT 4.74 1.21 4.97 1.34 ;
 RECT 4.74 1.11 5.14 1.21 ;
 RECT 1.01 0.19 1.11 1.16 ;
 RECT 1.01 1.37 1.11 2.305 ;
 RECT 2.79 0.19 2.89 0.88 ;
 RECT 1.01 2.305 1.265 2.515 ;
 RECT 0.82 1.16 1.11 1.37 ;
 RECT 1.01 0.09 2.89 0.19 ;
 RECT 1.7 1.425 1.95 1.535 ;
 RECT 1.85 0.37 1.95 1.425 ;
 RECT 2.02 1.635 2.12 2.135 ;
 RECT 1.7 1.535 2.12 1.635 ;
 RECT 0.54 0.555 0.64 2.12 ;
 RECT 0.38 2.12 0.64 2.33 ;
 LAYER CO ;
 RECT 7.91 2.305 8.04 2.435 ;
 RECT 8.38 1.515 8.51 1.645 ;
 RECT 8.85 2.305 8.98 2.435 ;
 RECT 7.91 1.78 8.04 1.91 ;
 RECT 8.85 0.78 8.98 0.91 ;
 RECT 9.32 2.045 9.45 2.175 ;
 RECT 9.32 2.305 9.45 2.435 ;
 RECT 7.44 2.045 7.57 2.175 ;
 RECT 6.97 1.515 7.1 1.645 ;
 RECT 7.91 2.045 8.04 2.175 ;
 RECT 8.85 1.78 8.98 1.91 ;
 RECT 6.97 0.52 7.1 0.65 ;
 RECT 9.32 1.78 9.45 1.91 ;
 RECT 7.44 2.305 7.57 2.435 ;
 RECT 6.5 2.305 6.63 2.435 ;
 RECT 9.72 1.805 9.85 1.935 ;
 RECT 1.085 2.345 1.215 2.475 ;
 RECT 9.72 1.545 9.85 1.675 ;
 RECT 1.6 0.59 1.73 0.72 ;
 RECT 3.01 1.775 3.14 1.905 ;
 RECT 2.54 1.775 2.67 1.905 ;
 RECT 3.51 1.205 3.64 1.335 ;
 RECT 2.185 1.18 2.315 1.31 ;
 RECT 0.29 0.775 0.42 0.905 ;
 RECT 1.77 2.625 1.9 2.755 ;
 RECT 7.91 0.52 8.04 0.65 ;
 RECT 4.25 1.775 4.38 1.905 ;
 RECT 7.91 1.515 8.04 1.645 ;
 RECT 0.29 1.63 0.42 1.76 ;
 RECT 2.07 0.59 2.2 0.72 ;
 RECT 3.925 0.925 4.055 1.055 ;
 RECT 4.79 0.52 4.92 0.65 ;
 RECT 1.23 2.015 1.36 2.145 ;
 RECT 4.52 2.43 4.65 2.56 ;
 RECT 0.76 0.775 0.89 0.905 ;
 RECT 0.87 1.2 1 1.33 ;
 RECT 1.75 1.465 1.88 1.595 ;
 RECT 0.43 2.16 0.56 2.29 ;
 RECT 1.23 0.775 1.36 0.905 ;
 RECT 5.56 2.045 5.69 2.175 ;
 RECT 5.56 1.775 5.69 1.905 ;
 RECT 4.79 0.78 4.92 0.91 ;
 RECT 8.38 2.045 8.51 2.175 ;
 RECT 6.97 1.78 7.1 1.91 ;
 RECT 7.44 1.515 7.57 1.645 ;
 RECT 9.72 0.665 9.85 0.795 ;
 RECT 3.78 0.53 3.91 0.66 ;
 RECT 9.72 0.405 9.85 0.535 ;
 RECT 0.76 1.66 0.89 1.79 ;
 RECT 5.09 1.515 5.22 1.645 ;
 RECT 4.25 0.595 4.38 0.725 ;
 RECT 3.19 2.395 3.32 2.525 ;
 RECT 3.01 0.53 3.14 0.66 ;
 RECT 9.72 2.065 9.85 2.195 ;
 RECT 6.5 0.78 6.63 0.91 ;
 RECT 8.38 1.78 8.51 1.91 ;
 RECT 9.32 0.52 9.45 0.65 ;
 RECT 6.03 0.78 6.16 0.91 ;
 RECT 6.97 2.045 7.1 2.175 ;
 RECT 6.03 0.52 6.16 0.65 ;
 RECT 2.755 2.065 2.885 2.195 ;
 RECT 4.79 1.16 4.92 1.29 ;
 RECT 5.23 2.465 5.36 2.595 ;
 RECT 5.56 0.49 5.69 0.62 ;
 RECT 6.03 1.78 6.16 1.91 ;
 RECT 6.5 0.52 6.63 0.65 ;
 RECT 6.03 2.045 6.16 2.175 ;
 RECT 6.5 1.515 6.63 1.645 ;
 RECT 7.91 0.78 8.04 0.91 ;
 RECT 8.85 0.52 8.98 0.65 ;
 RECT 6.03 1.515 6.16 1.645 ;
 RECT 5.56 1.515 5.69 1.645 ;
 RECT 8.38 0.78 8.51 0.91 ;
 RECT 8.38 2.305 8.51 2.435 ;
 RECT 3.73 2.39 3.86 2.52 ;
 RECT 2.54 0.59 2.67 0.72 ;
 RECT 9.32 1.515 9.45 1.645 ;
 RECT 8.38 0.52 8.51 0.65 ;
 RECT 6.97 0.78 7.1 0.91 ;
 RECT 6.03 2.305 6.16 2.435 ;
 RECT 6.5 2.045 6.63 2.175 ;
 RECT 7.44 1.78 7.57 1.91 ;
 RECT 7.44 0.78 7.57 0.91 ;
 RECT 6.5 1.78 6.63 1.91 ;
 RECT 5.695 1.115 5.825 1.245 ;
 RECT 9.32 0.78 9.45 0.91 ;
 RECT 6.97 2.305 7.1 2.435 ;
 RECT 8.85 1.515 8.98 1.645 ;
 RECT 7.44 0.52 7.57 0.65 ;
 RECT 8.85 2.045 8.98 2.175 ;
 LAYER M1 ;
 RECT 1.595 0.53 1.735 0.865 ;
 RECT 2.535 1.005 2.675 1.77 ;
 RECT 2.535 0.525 2.675 0.865 ;
 RECT 1.595 0.865 2.675 1.005 ;
 RECT 2.49 1.77 2.72 1.91 ;
 RECT 5.085 0.97 5.225 1.11 ;
 RECT 5.085 1.25 5.225 1.8 ;
 RECT 4.785 0.47 4.925 0.83 ;
 RECT 4.785 0.83 5.225 0.97 ;
 RECT 5.085 1.11 5.875 1.25 ;
 RECT 4.245 0.36 4.385 1.2 ;
 RECT 4.245 1.34 4.385 1.77 ;
 RECT 4.245 1.91 4.385 1.92 ;
 RECT 4.785 1.11 4.925 1.2 ;
 RECT 3.46 1.2 4.925 1.34 ;
 RECT 4.2 1.77 4.43 1.91 ;
 RECT 3.005 0.45 3.145 0.92 ;
 RECT 3.005 1.06 3.145 1.77 ;
 RECT 2.96 1.77 3.19 1.91 ;
 RECT 3.005 0.92 4.105 1.06 ;
 RECT 3.185 2.48 3.325 2.575 ;
 RECT 1.035 2.34 3.325 2.48 ;
 RECT 1.19 1.12 1.33 2.01 ;
 RECT 1.225 0.71 1.365 0.98 ;
 RECT 1.19 0.98 1.365 1.12 ;
 RECT 1.05 2.01 1.485 2.06 ;
 RECT 5.18 2.2 5.32 2.46 ;
 RECT 1.05 2.06 5.32 2.2 ;
 RECT 5.18 2.46 5.41 2.6 ;
 RECT 0.285 0.58 0.425 1.195 ;
 RECT 0.285 1.335 0.425 1.84 ;
 RECT 0.285 1.195 1.05 1.335 ;
 RECT 0.82 1.16 1.05 1.195 ;
 RECT 0.82 1.335 1.05 1.37 ;
 END
END CGLPPRX8

MACRO LSUPENCLX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.32 BY 5.76 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.32 2.96 ;
 RECT 1.685 3.395 1.945 3.535 ;
 RECT 1.325 2.085 1.6 2.225 ;
 RECT 2.46 2.96 2.88 3.645 ;
 RECT 2.285 2.02 2.425 2.8 ;
 RECT 3.255 2.1 3.395 2.8 ;
 RECT 4.22 2.1 4.36 2.8 ;
 RECT 5.185 2.1 5.325 2.8 ;
 RECT 6.2 2.1 6.34 2.8 ;
 RECT 6.975 2.1 7.115 2.8 ;
 RECT 6.975 2.96 7.115 3.475 ;
 RECT 1.75 3.535 1.89 3.58 ;
 RECT 1.75 2.96 1.89 3.395 ;
 RECT 1.425 2.225 1.565 2.8 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 3.72 1.96 3.745 ;
 RECT 2.05 3.11 2.32 3.25 ;
 RECT 1.555 3.885 1.96 4.04 ;
 RECT 1.555 3.745 2.255 3.885 ;
 RECT 2.115 3.25 2.255 3.745 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 8.32 5.2 ;
 RECT 2.07 4.26 2.49 4.665 ;
 RECT 2.215 4.665 2.355 5.04 ;
 RECT 1.745 4.3 1.885 5.04 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.6 1.475 2.905 1.81 ;
 RECT 2.765 0.935 2.905 1.475 ;
 RECT 7.445 2.4 7.93 2.62 ;
 RECT 2.765 1.82 7.595 1.96 ;
 RECT 2.765 1.96 2.905 2.29 ;
 RECT 2.765 1.81 2.905 1.82 ;
 RECT 3.745 1.96 3.885 2.29 ;
 RECT 3.745 0.935 3.885 1.82 ;
 RECT 4.715 1.96 4.855 2.29 ;
 RECT 4.715 0.935 4.855 1.82 ;
 RECT 5.71 1.96 5.85 2.29 ;
 RECT 5.71 0.935 5.85 1.82 ;
 RECT 7.445 1.96 7.585 2.4 ;
 END
 ANTENNADIFFAREA 2.218 ;
 END Q

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.8 4.17 7.3 4.755 ;
 END
 ANTENNAGATEAREA 0.16 ;
 END ENB

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.32 0.08 ;
 RECT 0.47 0.08 0.61 1.275 ;
 RECT 7.445 0.08 7.585 1.325 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 8.32 5.84 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 1.15 0.215 1.25 1.29 ;
 RECT 2.55 0.215 2.65 1.595 ;
 RECT 2.2 1.595 2.65 1.825 ;
 RECT 2.55 1.825 2.65 2.685 ;
 RECT 1.15 0.115 6.085 0.215 ;
 RECT 5.985 0.215 6.085 2.685 ;
 RECT 5.475 0.215 5.575 2.685 ;
 RECT 4.97 0.215 5.07 2.685 ;
 RECT 4.48 0.215 4.58 2.685 ;
 RECT 4 0.215 4.1 2.685 ;
 RECT 3.51 0.215 3.61 2.685 ;
 RECT 3.04 0.215 3.14 2.685 ;
 RECT 7.23 0.455 7.33 4.28 ;
 RECT 6.855 4.28 7.33 4.35 ;
 RECT 6.855 4.45 7.33 4.47 ;
 RECT 6.855 4.47 7.26 4.51 ;
 RECT 6.76 4.35 7.33 4.45 ;
 RECT 1.455 1.165 1.75 1.395 ;
 RECT 1.65 0.395 1.75 1.165 ;
 RECT 1 2.535 1.1 3.06 ;
 RECT 1.15 1.835 1.25 2.435 ;
 RECT 1 2.435 1.25 2.535 ;
 RECT 0.93 3.06 1.16 3.29 ;
 RECT 2.045 3.065 2.3 3.295 ;
 RECT 2.045 2.5 2.145 3.065 ;
 RECT 1.65 2.4 2.145 2.5 ;
 RECT 1.65 1.84 1.75 2.4 ;
 RECT 1.53 3.17 1.63 3.785 ;
 RECT 1.53 3.785 1.83 4.015 ;
 RECT 1.53 4.015 1.63 4.73 ;
 RECT 7.765 2.62 7.865 3.155 ;
 RECT 7.7 3.155 7.93 3.385 ;
 RECT 7.7 2.39 7.93 2.62 ;
 LAYER CO ;
 RECT 1.4 2.09 1.53 2.22 ;
 RECT 2.745 3.445 2.875 3.575 ;
 RECT 1.65 3.835 1.78 3.965 ;
 RECT 2.295 0.815 2.425 0.945 ;
 RECT 2.12 3.115 2.25 3.245 ;
 RECT 6.205 2.175 6.335 2.305 ;
 RECT 5.19 2.175 5.32 2.305 ;
 RECT 4.225 2.175 4.355 2.305 ;
 RECT 3.26 2.175 3.39 2.305 ;
 RECT 6.205 0.815 6.335 0.945 ;
 RECT 6.205 1.125 6.335 1.255 ;
 RECT 5.715 1.005 5.845 1.135 ;
 RECT 5.715 2.09 5.845 2.22 ;
 RECT 5.715 1.265 5.845 1.395 ;
 RECT 5.19 0.815 5.32 0.945 ;
 RECT 5.19 1.125 5.32 1.255 ;
 RECT 4.72 1.005 4.85 1.135 ;
 RECT 4.72 2.09 4.85 2.22 ;
 RECT 4.72 1.265 4.85 1.395 ;
 RECT 4.22 0.815 4.35 0.945 ;
 RECT 4.22 1.125 4.35 1.255 ;
 RECT 3.75 2.09 3.88 2.22 ;
 RECT 3.75 1.265 3.88 1.395 ;
 RECT 3.75 1.005 3.88 1.135 ;
 RECT 3.26 0.815 3.39 0.945 ;
 RECT 3.26 1.125 3.39 1.255 ;
 RECT 6.98 4.33 7.11 4.46 ;
 RECT 0.475 1.085 0.605 1.215 ;
 RECT 7.75 2.44 7.88 2.57 ;
 RECT 7.75 3.205 7.88 3.335 ;
 RECT 7.45 2.09 7.58 2.22 ;
 RECT 6.98 2.16 7.11 2.29 ;
 RECT 7.45 3.295 7.58 3.425 ;
 RECT 6.98 3.295 7.11 3.425 ;
 RECT 7.45 1.125 7.58 1.255 ;
 RECT 7.45 0.815 7.58 0.945 ;
 RECT 6.98 1.125 7.11 1.255 ;
 RECT 6.98 1.125 7.11 1.255 ;
 RECT 1.28 4.36 1.41 4.49 ;
 RECT 0.475 0.825 0.605 0.955 ;
 RECT 2.77 1.005 2.9 1.135 ;
 RECT 1.87 2.09 2 2.22 ;
 RECT 2.29 2.09 2.42 2.22 ;
 RECT 2.745 3.185 2.875 3.315 ;
 RECT 1.4 0.83 1.53 0.96 ;
 RECT 1.755 3.4 1.885 3.53 ;
 RECT 1.505 1.215 1.635 1.345 ;
 RECT 2.295 1.125 2.425 1.255 ;
 RECT 0.9 0.835 1.03 0.965 ;
 RECT 1.28 3.4 1.41 3.53 ;
 RECT 2.77 2.09 2.9 2.22 ;
 RECT 0.98 3.11 1.11 3.24 ;
 RECT 0.475 0.565 0.605 0.695 ;
 RECT 1.75 4.37 1.88 4.5 ;
 RECT 1.87 0.815 2 0.945 ;
 RECT 2.465 3.185 2.595 3.315 ;
 RECT 0.9 2.09 1.03 2.22 ;
 RECT 2.225 4.3 2.355 4.43 ;
 RECT 2.25 1.645 2.38 1.775 ;
 RECT 2.77 1.265 2.9 1.395 ;
 RECT 2.465 3.445 2.595 3.575 ;
 RECT 7.75 2.44 7.88 2.57 ;
 LAYER M1 ;
 RECT 5.185 0.38 5.325 1.385 ;
 RECT 4.215 0.38 4.355 1.385 ;
 RECT 3.255 0.38 3.395 1.385 ;
 RECT 1.395 0.38 1.535 1.02 ;
 RECT 2.29 0.38 2.43 1.385 ;
 RECT 6.975 0.38 7.115 1.325 ;
 RECT 6.2 0.38 6.34 1.385 ;
 RECT 1.395 0.24 7.115 0.38 ;
 RECT 0.895 0.76 1.035 1.45 ;
 RECT 0.895 1.59 1.035 2.29 ;
 RECT 1.5 1.165 1.64 1.45 ;
 RECT 0.895 1.45 1.64 1.59 ;
 RECT 1.275 3.245 1.415 4.56 ;
 RECT 0.93 3.105 1.415 3.245 ;
 RECT 7.39 3.1 7.985 3.51 ;
 RECT 1.865 0.745 2.005 1.64 ;
 RECT 1.865 1.78 2.005 2.29 ;
 RECT 1.865 1.64 2.46 1.78 ;
 RECT 2.2 1.6 2.46 1.64 ;
 RECT 2.2 1.78 2.46 1.83 ;
 END
END LSUPENCLX4

MACRO CGLPPSX16
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 16.32 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.04 1.765 4.41 2.04 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END SE

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 16.32 2.96 ;
 RECT 4.51 1.525 4.74 1.665 ;
 RECT 1.53 2.355 1.67 2.8 ;
 RECT 8.625 1.43 8.765 2.8 ;
 RECT 11.445 1.43 11.585 2.8 ;
 RECT 12.385 1.43 12.525 2.8 ;
 RECT 0.695 1.66 0.835 2.8 ;
 RECT 3.245 1.73 3.385 2.8 ;
 RECT 5.42 1.95 5.56 2.8 ;
 RECT 5.71 2.325 5.85 2.8 ;
 RECT 13.325 1.43 13.465 2.8 ;
 RECT 14.265 1.43 14.405 2.8 ;
 RECT 15.205 1.43 15.345 2.8 ;
 RECT 7.685 1.43 7.825 2.8 ;
 RECT 9.565 1.43 9.705 2.8 ;
 RECT 6.745 1.44 6.885 2.8 ;
 RECT 10.505 1.43 10.645 2.8 ;
 RECT 15.725 1.5 15.865 2.8 ;
 RECT 4.55 1.665 4.69 2.8 ;
 END
 END VDD

 PIN EN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.56 1.115 1.865 1.405 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END EN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 16.32 0.08 ;
 RECT 1.485 0.585 1.74 0.725 ;
 RECT 4.51 0.585 4.74 0.725 ;
 RECT 14.265 0.08 14.405 0.975 ;
 RECT 7.685 0.08 7.825 0.94 ;
 RECT 10.505 0.08 10.645 0.975 ;
 RECT 3.245 0.08 3.385 0.74 ;
 RECT 1.6 0.08 1.74 0.585 ;
 RECT 13.325 0.08 13.465 0.975 ;
 RECT 12.385 0.08 12.525 0.975 ;
 RECT 15.205 0.08 15.345 0.975 ;
 RECT 0.695 0.08 0.835 0.985 ;
 RECT 9.565 0.08 9.705 0.975 ;
 RECT 11.445 0.08 11.585 0.975 ;
 RECT 5.805 0.08 5.945 0.785 ;
 RECT 8.625 0.08 8.765 0.975 ;
 RECT 15.725 0.08 15.865 0.85 ;
 RECT 4.555 0.08 4.695 0.585 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 2.105 0.555 2.36 ;
 END
 ANTENNAGATEAREA 0.063 ;
 END CLK

 PIN GCLK
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.6 1.48 14.875 1.72 ;
 RECT 14.735 1.72 14.875 2.45 ;
 RECT 12.855 1.26 12.995 2.45 ;
 RECT 12.855 0.475 12.995 1.12 ;
 RECT 13.795 1.26 13.935 2.45 ;
 RECT 13.795 0.475 13.935 1.12 ;
 RECT 11.915 1.26 12.055 2.45 ;
 RECT 11.915 0.475 12.055 1.12 ;
 RECT 10.975 1.26 11.115 2.45 ;
 RECT 10.975 0.475 11.115 1.12 ;
 RECT 10.035 1.26 10.175 2.45 ;
 RECT 10.035 0.475 10.175 1.12 ;
 RECT 8.155 1.26 8.295 2.45 ;
 RECT 8.155 0.475 8.295 1.12 ;
 RECT 9.095 1.26 9.235 2.45 ;
 RECT 9.095 0.475 9.235 1.12 ;
 RECT 8.155 1.12 14.875 1.26 ;
 RECT 14.735 1.26 14.875 1.48 ;
 RECT 14.735 0.475 14.875 1.12 ;
 END
 ANTENNADIFFAREA 4.976 ;
 END GCLK

 OBS
 LAYER PO ;
 RECT 4.81 0.19 4.91 1.88 ;
 RECT 3.5 0.19 3.6 0.89 ;
 RECT 3.5 1.1 3.6 2.14 ;
 RECT 3.345 0.89 3.6 1.1 ;
 RECT 3.5 0.09 4.91 0.19 ;
 RECT 5.11 1.2 5.345 1.23 ;
 RECT 5.11 0.37 5.21 1.2 ;
 RECT 5.115 1.33 5.38 1.41 ;
 RECT 5.28 1.41 5.38 1.88 ;
 RECT 5.11 1.23 5.38 1.33 ;
 RECT 3.03 0.315 3.13 1.17 ;
 RECT 3.03 1.38 3.13 2.14 ;
 RECT 2.93 1.17 3.16 1.38 ;
 RECT 7.47 0.09 7.57 2.625 ;
 RECT 6.06 0.09 6.16 2.625 ;
 RECT 2.885 2.625 7.57 2.725 ;
 RECT 2.885 2.43 3.095 2.625 ;
 RECT 2.73 0.315 2.83 0.89 ;
 RECT 2.26 1.26 2.36 2.03 ;
 RECT 2.65 0.89 2.83 0.99 ;
 RECT 2.65 0.99 2.75 1.16 ;
 RECT 2.26 1.16 2.75 1.26 ;
 RECT 2.185 2.03 2.415 2.24 ;
 RECT 7 0.09 7.1 2.22 ;
 RECT 6.53 0.09 6.63 2.215 ;
 RECT 6.4 2.215 6.63 2.22 ;
 RECT 6.4 2.32 6.63 2.445 ;
 RECT 6.4 2.22 7.1 2.32 ;
 RECT 7.775 1.08 8.04 1.15 ;
 RECT 7.775 1.25 8.04 1.29 ;
 RECT 7.94 1.29 8.04 2.74 ;
 RECT 9.82 0.22 9.92 1.15 ;
 RECT 9.82 1.25 9.92 2.74 ;
 RECT 7.94 0.22 8.04 1.08 ;
 RECT 7.775 1.15 15.09 1.25 ;
 RECT 14.99 1.25 15.09 2.74 ;
 RECT 14.99 0.22 15.09 1.15 ;
 RECT 12.64 1.25 12.74 2.74 ;
 RECT 12.64 0.22 12.74 1.15 ;
 RECT 13.11 0.22 13.21 1.15 ;
 RECT 13.11 1.25 13.21 2.74 ;
 RECT 14.52 0.22 14.62 1.15 ;
 RECT 14.52 1.25 14.62 2.74 ;
 RECT 13.58 1.25 13.68 2.74 ;
 RECT 13.58 0.22 13.68 1.15 ;
 RECT 14.05 1.25 14.15 2.74 ;
 RECT 14.05 0.22 14.15 1.15 ;
 RECT 12.17 0.22 12.27 1.15 ;
 RECT 12.17 1.25 12.27 2.74 ;
 RECT 11.7 1.25 11.8 2.74 ;
 RECT 11.7 0.22 11.8 1.15 ;
 RECT 8.41 0.22 8.51 1.15 ;
 RECT 8.41 1.25 8.51 2.74 ;
 RECT 9.35 1.25 9.45 2.74 ;
 RECT 9.35 0.22 9.45 1.15 ;
 RECT 10.76 1.25 10.86 2.74 ;
 RECT 10.76 0.22 10.86 1.15 ;
 RECT 8.88 0.22 8.98 1.15 ;
 RECT 8.88 1.25 8.98 2.74 ;
 RECT 10.29 1.25 10.39 2.74 ;
 RECT 10.29 0.22 10.39 1.15 ;
 RECT 11.23 1.25 11.33 2.74 ;
 RECT 11.23 0.22 11.33 1.15 ;
 RECT 1.79 1.4 1.89 2.14 ;
 RECT 1.79 0.37 1.89 1.19 ;
 RECT 1.615 1.19 1.89 1.4 ;
 RECT 0.95 1.34 1.05 2.655 ;
 RECT 0.95 0.19 1.05 1.13 ;
 RECT 2.73 1.56 2.83 2.035 ;
 RECT 2.6 2.135 2.7 2.655 ;
 RECT 2.6 2.035 2.83 2.135 ;
 RECT 0.95 2.655 2.7 2.755 ;
 RECT 2.26 0.19 2.36 0.885 ;
 RECT 0.78 1.13 1.05 1.34 ;
 RECT 0.95 0.09 2.36 0.19 ;
 RECT 4.34 0.37 4.44 1.78 ;
 RECT 4.175 1.78 4.44 1.99 ;
 RECT 0.48 0.57 0.58 2.12 ;
 RECT 0.325 2.12 0.58 2.33 ;
 LAYER CO ;
 RECT 13.33 1.48 13.46 1.61 ;
 RECT 14.27 2.01 14.4 2.14 ;
 RECT 13.8 1.48 13.93 1.61 ;
 RECT 14.74 2.01 14.87 2.14 ;
 RECT 0.83 1.17 0.96 1.3 ;
 RECT 4.225 1.82 4.355 1.95 ;
 RECT 0.375 2.16 0.505 2.29 ;
 RECT 13.33 2.01 13.46 2.14 ;
 RECT 11.92 2.27 12.05 2.4 ;
 RECT 15.21 2.27 15.34 2.4 ;
 RECT 14.27 1.745 14.4 1.875 ;
 RECT 13.8 1.745 13.93 1.875 ;
 RECT 15.21 2.01 15.34 2.14 ;
 RECT 11.92 2.01 12.05 2.14 ;
 RECT 15.73 0.41 15.86 0.54 ;
 RECT 3.395 0.93 3.525 1.06 ;
 RECT 2.235 2.07 2.365 2.2 ;
 RECT 8.63 0.525 8.76 0.655 ;
 RECT 10.04 0.525 10.17 0.655 ;
 RECT 7.69 1.74 7.82 1.87 ;
 RECT 11.45 0.525 11.58 0.655 ;
 RECT 8.63 1.745 8.76 1.875 ;
 RECT 8.16 0.785 8.29 0.915 ;
 RECT 10.04 2.27 10.17 2.4 ;
 RECT 10.98 2.27 11.11 2.4 ;
 RECT 8.16 2.01 8.29 2.14 ;
 RECT 10.51 0.525 10.64 0.655 ;
 RECT 8.16 0.525 8.29 0.655 ;
 RECT 10.51 1.48 10.64 1.61 ;
 RECT 7.69 0.495 7.82 0.625 ;
 RECT 11.45 1.745 11.58 1.875 ;
 RECT 9.1 1.48 9.23 1.61 ;
 RECT 8.63 2.01 8.76 2.14 ;
 RECT 9.1 0.785 9.23 0.915 ;
 RECT 9.1 0.525 9.23 0.655 ;
 RECT 9.1 2.27 9.23 2.4 ;
 RECT 11.92 1.745 12.05 1.875 ;
 RECT 11.92 0.785 12.05 0.915 ;
 RECT 11.92 0.525 12.05 0.655 ;
 RECT 14.74 1.48 14.87 1.61 ;
 RECT 15.21 1.745 15.34 1.875 ;
 RECT 13.33 2.27 13.46 2.4 ;
 RECT 8.16 2.27 8.29 2.4 ;
 RECT 10.04 1.745 10.17 1.875 ;
 RECT 0.23 1.585 0.36 1.715 ;
 RECT 4.09 0.59 4.22 0.72 ;
 RECT 10.98 1.745 11.11 1.875 ;
 RECT 5.33 0.59 5.46 0.72 ;
 RECT 11.45 2.27 11.58 2.4 ;
 RECT 10.51 2.27 10.64 2.4 ;
 RECT 9.57 2.01 9.7 2.14 ;
 RECT 9.57 1.745 9.7 1.875 ;
 RECT 7.69 2.01 7.82 2.14 ;
 RECT 0.23 0.79 0.36 0.92 ;
 RECT 15.73 1.81 15.86 1.94 ;
 RECT 4.56 1.53 4.69 1.66 ;
 RECT 8.63 1.48 8.76 1.61 ;
 RECT 9.57 0.785 9.7 0.915 ;
 RECT 3.25 0.535 3.38 0.665 ;
 RECT 6.75 1.49 6.88 1.62 ;
 RECT 10.98 0.525 11.11 0.655 ;
 RECT 15.73 0.67 15.86 0.8 ;
 RECT 9.57 2.27 9.7 2.4 ;
 RECT 4.09 1.49 4.22 1.62 ;
 RECT 3.25 1.78 3.38 1.91 ;
 RECT 8.16 1.48 8.29 1.61 ;
 RECT 11.45 0.785 11.58 0.915 ;
 RECT 8.16 1.745 8.29 1.875 ;
 RECT 15.73 2.07 15.86 2.2 ;
 RECT 2.925 2.48 3.055 2.61 ;
 RECT 7.22 0.31 7.35 0.44 ;
 RECT 7.22 0.57 7.35 0.7 ;
 RECT 6.75 0.785 6.88 0.915 ;
 RECT 6.28 0.31 6.41 0.44 ;
 RECT 6.28 0.57 6.41 0.7 ;
 RECT 5.81 0.57 5.94 0.7 ;
 RECT 7.22 1.75 7.35 1.88 ;
 RECT 7.22 1.49 7.35 1.62 ;
 RECT 12.86 1.48 12.99 1.61 ;
 RECT 15.21 1.48 15.34 1.61 ;
 RECT 10.51 0.785 10.64 0.915 ;
 RECT 2.01 1.78 2.14 1.91 ;
 RECT 7.69 1.48 7.82 1.61 ;
 RECT 10.51 2.01 10.64 2.14 ;
 RECT 1.17 1.5 1.3 1.63 ;
 RECT 2.98 1.21 3.11 1.34 ;
 RECT 7.825 1.12 7.955 1.25 ;
 RECT 9.1 2.01 9.23 2.14 ;
 RECT 13.8 0.785 13.93 0.915 ;
 RECT 14.74 1.745 14.87 1.875 ;
 RECT 6.75 1.75 6.88 1.88 ;
 RECT 10.04 2.01 10.17 2.14 ;
 RECT 3.72 0.6 3.85 0.73 ;
 RECT 10.04 0.785 10.17 0.915 ;
 RECT 0.7 0.79 0.83 0.92 ;
 RECT 5.165 1.24 5.295 1.37 ;
 RECT 10.98 0.785 11.11 0.915 ;
 RECT 9.57 1.48 9.7 1.61 ;
 RECT 10.98 2.01 11.11 2.14 ;
 RECT 9.1 1.745 9.23 1.875 ;
 RECT 7.69 0.76 7.82 0.89 ;
 RECT 1.535 2.405 1.665 2.535 ;
 RECT 15.21 0.525 15.34 0.655 ;
 RECT 13.33 1.745 13.46 1.875 ;
 RECT 14.74 0.525 14.87 0.655 ;
 RECT 12.39 0.525 12.52 0.655 ;
 RECT 15.21 0.785 15.34 0.915 ;
 RECT 12.39 1.745 12.52 1.875 ;
 RECT 14.27 0.525 14.4 0.655 ;
 RECT 2.48 1.78 2.61 1.91 ;
 RECT 8.63 0.785 8.76 0.915 ;
 RECT 10.51 1.745 10.64 1.875 ;
 RECT 11.45 2.01 11.58 2.14 ;
 RECT 2.01 0.59 2.14 0.72 ;
 RECT 5.81 0.31 5.94 0.44 ;
 RECT 5.425 2 5.555 2.13 ;
 RECT 12.39 2.27 12.52 2.4 ;
 RECT 12.86 1.745 12.99 1.875 ;
 RECT 13.8 0.525 13.93 0.655 ;
 RECT 14.27 1.48 14.4 1.61 ;
 RECT 12.39 2.01 12.52 2.14 ;
 RECT 14.27 0.785 14.4 0.915 ;
 RECT 13.8 2.27 13.93 2.4 ;
 RECT 12.86 0.785 12.99 0.915 ;
 RECT 12.39 1.48 12.52 1.61 ;
 RECT 14.74 2.27 14.87 2.4 ;
 RECT 12.86 0.525 12.99 0.655 ;
 RECT 13.33 0.785 13.46 0.915 ;
 RECT 12.86 2.01 12.99 2.14 ;
 RECT 13.33 0.525 13.46 0.655 ;
 RECT 12.86 2.27 12.99 2.4 ;
 RECT 13.8 2.01 13.93 2.14 ;
 RECT 14.74 0.785 14.87 0.915 ;
 RECT 11.92 1.48 12.05 1.61 ;
 RECT 4.56 0.59 4.69 0.72 ;
 RECT 5.715 2.375 5.845 2.505 ;
 RECT 1.665 1.23 1.795 1.36 ;
 RECT 10.98 1.48 11.11 1.61 ;
 RECT 2.48 0.535 2.61 0.665 ;
 RECT 7.69 2.27 7.82 2.4 ;
 RECT 9.57 0.525 9.7 0.655 ;
 RECT 15.73 1.55 15.86 1.68 ;
 RECT 11.45 1.48 11.58 1.61 ;
 RECT 6.28 1.75 6.41 1.88 ;
 RECT 0.7 1.71 0.83 1.84 ;
 RECT 3.72 1.78 3.85 1.91 ;
 RECT 1.54 0.59 1.67 0.72 ;
 RECT 5.03 1.53 5.16 1.66 ;
 RECT 8.63 2.27 8.76 2.4 ;
 RECT 10.04 1.48 10.17 1.61 ;
 RECT 6.28 1.49 6.41 1.62 ;
 RECT 1.17 0.79 1.3 0.92 ;
 RECT 6.45 2.26 6.58 2.39 ;
 RECT 14.27 2.27 14.4 2.4 ;
 RECT 12.39 0.785 12.52 0.915 ;
 LAYER M1 ;
 RECT 7.215 0.4 7.355 0.76 ;
 RECT 6.275 0.26 7.355 0.4 ;
 RECT 6.275 0.4 6.415 0.75 ;
 RECT 2.475 0.455 2.615 0.925 ;
 RECT 2.475 1.065 2.615 1.775 ;
 RECT 2.43 1.775 2.66 1.915 ;
 RECT 2.475 0.925 3.575 1.065 ;
 RECT 2.005 0.53 2.145 1.775 ;
 RECT 1.96 1.775 2.19 1.915 ;
 RECT 6.275 1.105 7.355 1.11 ;
 RECT 7.215 1.25 7.355 1.93 ;
 RECT 6.745 0.73 6.885 1.105 ;
 RECT 6.275 1.245 6.415 1.93 ;
 RECT 7.215 1.245 8.005 1.25 ;
 RECT 6.275 1.115 8.005 1.245 ;
 RECT 6.275 1.11 7.96 1.115 ;
 RECT 7.775 1.25 8.005 1.255 ;
 RECT 2.93 1.205 3.855 1.345 ;
 RECT 3.715 0.365 3.855 1.205 ;
 RECT 3.715 1.345 3.855 2 ;
 RECT 5.525 0.725 5.665 1.525 ;
 RECT 5.28 0.585 5.665 0.725 ;
 RECT 4.98 1.525 6.13 1.665 ;
 RECT 5.99 1.665 6.13 2.07 ;
 RECT 6.445 2.21 6.585 2.445 ;
 RECT 5.99 2.07 6.585 2.21 ;
 RECT 1.165 0.715 1.305 1.545 ;
 RECT 1.675 2.065 3.06 2.205 ;
 RECT 2.92 2.205 3.06 2.66 ;
 RECT 1.165 1.545 1.815 1.685 ;
 RECT 1.675 1.685 1.815 2.065 ;
 RECT 4.04 1.385 4.305 1.625 ;
 RECT 4.085 0.505 4.225 1.245 ;
 RECT 4.04 1.245 5.345 1.375 ;
 RECT 5.115 1.235 5.345 1.245 ;
 RECT 4.04 1.375 5.295 1.385 ;
 RECT 0.225 0.52 0.365 1.165 ;
 RECT 0.225 1.305 0.365 1.81 ;
 RECT 0.225 1.165 1.01 1.305 ;
 RECT 0.78 1.13 1.01 1.165 ;
 RECT 0.78 1.305 1.01 1.34 ;
 END
END CGLPPSX16

MACRO LSUPENCLX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 15.36 BY 5.76 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 15.36 2.96 ;
 RECT 1.685 3.395 1.945 3.535 ;
 RECT 1.325 2.085 1.6 2.225 ;
 RECT 2.46 2.96 2.88 3.645 ;
 RECT 14.775 2.1 14.915 2.8 ;
 RECT 2.285 2.02 2.425 2.8 ;
 RECT 3.255 2.1 3.395 2.8 ;
 RECT 4.22 2.1 4.36 2.8 ;
 RECT 5.185 2.1 5.325 2.8 ;
 RECT 6.2 2.1 6.34 2.8 ;
 RECT 7.195 2.1 7.335 2.8 ;
 RECT 8.18 2.1 8.32 2.8 ;
 RECT 9.165 2.1 9.305 2.8 ;
 RECT 10.155 2.1 10.295 2.8 ;
 RECT 12.875 2.1 13.015 2.8 ;
 RECT 13.815 2.1 13.955 2.8 ;
 RECT 1.75 3.535 1.89 3.58 ;
 RECT 1.75 2.96 1.89 3.395 ;
 RECT 1.425 2.225 1.565 2.8 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 3.885 1.96 4.04 ;
 RECT 1.555 3.72 1.96 3.745 ;
 RECT 2.05 3.11 2.32 3.25 ;
 RECT 1.555 3.745 2.255 3.885 ;
 RECT 2.115 3.25 2.255 3.745 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 15.36 5.2 ;
 RECT 2.07 4.26 2.49 4.665 ;
 RECT 2.215 4.665 2.355 5.04 ;
 RECT 1.745 4.3 1.885 5.04 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.6 1.475 2.905 1.81 ;
 RECT 2.765 0.935 2.905 1.475 ;
 RECT 2.765 1.82 14.43 1.96 ;
 RECT 2.765 1.96 2.905 2.29 ;
 RECT 2.765 1.81 2.905 1.82 ;
 RECT 14.29 1.96 14.43 2.295 ;
 RECT 3.745 1.96 3.885 2.29 ;
 RECT 3.745 0.935 3.885 1.82 ;
 RECT 4.715 1.96 4.855 2.29 ;
 RECT 4.715 0.935 4.855 1.82 ;
 RECT 5.71 1.96 5.85 2.29 ;
 RECT 5.71 0.935 5.85 1.82 ;
 RECT 6.705 1.96 6.845 2.29 ;
 RECT 6.705 0.935 6.845 1.82 ;
 RECT 7.69 1.96 7.83 2.29 ;
 RECT 7.69 0.935 7.83 1.82 ;
 RECT 8.675 1.96 8.815 2.29 ;
 RECT 8.675 0.935 8.815 1.82 ;
 RECT 9.665 1.96 9.805 2.29 ;
 RECT 9.665 0.935 9.805 1.82 ;
 RECT 10.645 0.935 10.785 1.82 ;
 RECT 11.615 0.935 11.755 1.82 ;
 RECT 13.345 1.96 13.485 2.295 ;
 END
 ANTENNADIFFAREA 6.91 ;
 END Q

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.7 4.17 13.2 4.755 ;
 END
 ANTENNAGATEAREA 0.6 ;
 END ENB

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 15.36 0.08 ;
 RECT 0.47 0.08 0.61 1.275 ;
 RECT 13.345 0.08 13.485 1.325 ;
 RECT 14.295 0.08 14.435 1.325 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 15.36 5.84 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 12.755 4.28 13.23 4.35 ;
 RECT 13.13 1.845 13.23 4.28 ;
 RECT 12.755 4.47 13.16 4.51 ;
 RECT 12.755 4.45 13.23 4.47 ;
 RECT 13.6 0.32 13.7 1.745 ;
 RECT 13.13 0.32 13.23 1.745 ;
 RECT 13.6 1.845 13.7 2.76 ;
 RECT 14.55 0.32 14.65 1.745 ;
 RECT 14.55 1.845 14.65 2.77 ;
 RECT 14.07 0.32 14.17 1.745 ;
 RECT 14.07 1.845 14.17 2.775 ;
 RECT 13.13 1.745 14.65 1.845 ;
 RECT 12.66 4.35 13.23 4.45 ;
 RECT 1.455 1.165 1.75 1.395 ;
 RECT 1.65 0.395 1.75 1.165 ;
 RECT 0.93 3.06 1.25 3.225 ;
 RECT 1.15 1.765 1.25 3.06 ;
 RECT 0.93 3.225 1.16 3.29 ;
 RECT 2.045 3.065 2.3 3.295 ;
 RECT 2.045 2.5 2.145 3.065 ;
 RECT 1.65 2.4 2.145 2.5 ;
 RECT 1.65 1.84 1.75 2.4 ;
 RECT 1.53 3.17 1.63 3.785 ;
 RECT 1.53 3.785 1.83 4.015 ;
 RECT 1.53 4.015 1.63 4.73 ;
 RECT 2.55 0.215 2.65 1.595 ;
 RECT 2.2 1.595 2.65 1.825 ;
 RECT 2.55 1.825 2.65 2.905 ;
 RECT 1.15 0.215 1.25 1.29 ;
 RECT 5.985 0.215 6.085 2.935 ;
 RECT 5.475 0.215 5.575 2.935 ;
 RECT 4.97 0.215 5.07 2.935 ;
 RECT 4.48 0.215 4.58 2.935 ;
 RECT 4 0.215 4.1 2.935 ;
 RECT 3.51 0.215 3.61 2.935 ;
 RECT 3.04 0.215 3.14 2.935 ;
 RECT 11.9 0.215 12 1.635 ;
 RECT 11.4 0.215 11.5 1.635 ;
 RECT 10.915 0.215 11.015 1.635 ;
 RECT 8.44 0.215 8.54 2.935 ;
 RECT 8.95 0.215 9.05 2.935 ;
 RECT 7.455 0.215 7.555 2.935 ;
 RECT 7.965 0.215 8.065 2.935 ;
 RECT 6.47 0.215 6.57 2.935 ;
 RECT 6.98 0.215 7.08 2.935 ;
 RECT 10.41 0.215 10.51 1.635 ;
 RECT 9.43 0.215 9.53 2.935 ;
 RECT 9.94 0.215 10.04 2.935 ;
 RECT 1.15 0.115 12 0.215 ;
 LAYER CO ;
 RECT 11.14 0.815 11.27 0.945 ;
 RECT 10.65 1.005 10.78 1.135 ;
 RECT 10.65 1.265 10.78 1.395 ;
 RECT 10.16 0.815 10.29 0.945 ;
 RECT 9.67 1.265 9.8 1.395 ;
 RECT 10.16 1.125 10.29 1.255 ;
 RECT 9.67 1.005 9.8 1.135 ;
 RECT 8.68 2.09 8.81 2.22 ;
 RECT 9.17 2.175 9.3 2.305 ;
 RECT 9.17 0.815 9.3 0.945 ;
 RECT 8.68 1.265 8.81 1.395 ;
 RECT 9.17 1.125 9.3 1.255 ;
 RECT 8.68 1.005 8.81 1.135 ;
 RECT 7.695 2.09 7.825 2.22 ;
 RECT 8.185 2.175 8.315 2.305 ;
 RECT 8.185 0.815 8.315 0.945 ;
 RECT 7.695 1.265 7.825 1.395 ;
 RECT 8.185 1.125 8.315 1.255 ;
 RECT 7.695 1.005 7.825 1.135 ;
 RECT 1.505 1.215 1.635 1.345 ;
 RECT 2.295 1.125 2.425 1.255 ;
 RECT 0.9 0.835 1.03 0.965 ;
 RECT 1.28 3.4 1.41 3.53 ;
 RECT 2.77 2.09 2.9 2.22 ;
 RECT 0.98 3.11 1.11 3.24 ;
 RECT 0.475 0.565 0.605 0.695 ;
 RECT 1.75 4.37 1.88 4.5 ;
 RECT 1.87 0.815 2 0.945 ;
 RECT 2.465 3.185 2.595 3.315 ;
 RECT 0.9 2.09 1.03 2.22 ;
 RECT 2.225 4.3 2.355 4.43 ;
 RECT 2.25 1.645 2.38 1.775 ;
 RECT 2.77 1.265 2.9 1.395 ;
 RECT 2.465 3.445 2.595 3.575 ;
 RECT 1.4 2.09 1.53 2.22 ;
 RECT 2.745 3.445 2.875 3.575 ;
 RECT 1.65 3.835 1.78 3.965 ;
 RECT 2.295 0.815 2.425 0.945 ;
 RECT 2.12 3.115 2.25 3.245 ;
 RECT 6.71 2.09 6.84 2.22 ;
 RECT 7.2 2.175 7.33 2.305 ;
 RECT 7.2 0.815 7.33 0.945 ;
 RECT 6.71 1.265 6.84 1.395 ;
 RECT 7.2 1.125 7.33 1.255 ;
 RECT 6.71 1.005 6.84 1.135 ;
 RECT 6.205 2.175 6.335 2.305 ;
 RECT 5.19 2.175 5.32 2.305 ;
 RECT 4.225 2.175 4.355 2.305 ;
 RECT 9.67 2.09 9.8 2.22 ;
 RECT 10.16 2.175 10.29 2.305 ;
 RECT 3.26 2.175 3.39 2.305 ;
 RECT 6.205 0.815 6.335 0.945 ;
 RECT 6.205 1.125 6.335 1.255 ;
 RECT 5.715 1.005 5.845 1.135 ;
 RECT 5.715 2.09 5.845 2.22 ;
 RECT 5.715 1.265 5.845 1.395 ;
 RECT 5.19 0.815 5.32 0.945 ;
 RECT 5.19 1.125 5.32 1.255 ;
 RECT 4.72 1.005 4.85 1.135 ;
 RECT 4.72 2.09 4.85 2.22 ;
 RECT 4.72 1.265 4.85 1.395 ;
 RECT 4.22 0.815 4.35 0.945 ;
 RECT 4.22 1.125 4.35 1.255 ;
 RECT 3.75 2.09 3.88 2.22 ;
 RECT 3.75 1.265 3.88 1.395 ;
 RECT 3.75 1.005 3.88 1.135 ;
 RECT 3.26 0.815 3.39 0.945 ;
 RECT 3.26 1.125 3.39 1.255 ;
 RECT 12.88 4.33 13.01 4.46 ;
 RECT 0.475 1.085 0.605 1.215 ;
 RECT 13.35 2.09 13.48 2.22 ;
 RECT 12.88 2.16 13.01 2.29 ;
 RECT 13.35 1.125 13.48 1.255 ;
 RECT 13.35 0.815 13.48 0.945 ;
 RECT 12.88 1.125 13.01 1.255 ;
 RECT 12.88 1.125 13.01 1.255 ;
 RECT 1.28 4.36 1.41 4.49 ;
 RECT 0.475 0.825 0.605 0.955 ;
 RECT 2.77 1.005 2.9 1.135 ;
 RECT 1.87 2.09 2 2.22 ;
 RECT 2.29 2.09 2.42 2.22 ;
 RECT 2.745 3.185 2.875 3.315 ;
 RECT 1.4 0.83 1.53 0.96 ;
 RECT 1.755 3.4 1.885 3.53 ;
 RECT 14.78 2.16 14.91 2.29 ;
 RECT 14.295 2.09 14.425 2.22 ;
 RECT 13.82 2.16 13.95 2.29 ;
 RECT 14.77 1.125 14.9 1.255 ;
 RECT 14.77 1.125 14.9 1.255 ;
 RECT 14.3 0.815 14.43 0.945 ;
 RECT 14.3 1.125 14.43 1.255 ;
 RECT 13.82 1.125 13.95 1.255 ;
 RECT 13.82 1.125 13.95 1.255 ;
 RECT 12.12 1.125 12.25 1.255 ;
 RECT 12.12 0.815 12.25 0.945 ;
 RECT 11.62 1.005 11.75 1.135 ;
 RECT 11.62 1.265 11.75 1.395 ;
 RECT 11.14 1.125 11.27 1.255 ;
 LAYER M1 ;
 RECT 0.895 0.76 1.035 1.45 ;
 RECT 0.895 1.59 1.035 2.29 ;
 RECT 1.5 1.165 1.64 1.45 ;
 RECT 0.895 1.45 1.64 1.59 ;
 RECT 13.815 0.585 13.955 1.54 ;
 RECT 11.135 0.38 11.275 1.385 ;
 RECT 10.155 0.38 10.295 1.385 ;
 RECT 9.165 0.38 9.305 1.385 ;
 RECT 8.18 0.38 8.32 1.385 ;
 RECT 7.195 0.38 7.335 1.385 ;
 RECT 6.2 0.38 6.34 1.385 ;
 RECT 5.185 0.38 5.325 1.385 ;
 RECT 4.215 0.38 4.355 1.385 ;
 RECT 3.255 0.38 3.395 1.385 ;
 RECT 1.395 0.38 1.535 1.02 ;
 RECT 2.29 0.38 2.43 1.385 ;
 RECT 12.875 0.38 13.015 1.54 ;
 RECT 1.395 0.24 13.015 0.38 ;
 RECT 12.115 0.38 12.255 1.385 ;
 RECT 14.765 0.575 14.905 1.54 ;
 RECT 12.875 1.54 14.905 1.68 ;
 RECT 1.275 3.245 1.415 4.56 ;
 RECT 0.93 3.105 1.415 3.245 ;
 RECT 1.865 0.745 2.005 1.64 ;
 RECT 1.865 1.78 2.005 2.29 ;
 RECT 1.865 1.64 2.46 1.78 ;
 RECT 2.2 1.6 2.46 1.64 ;
 RECT 2.2 1.78 2.46 1.83 ;
 END
END LSUPENCLX8

MACRO LSUPENX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 5.76 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 1.685 3.395 1.945 3.535 ;
 RECT 2.46 2.96 2.88 3.645 ;
 RECT 3.63 2.1 3.77 2.8 ;
 RECT 3.63 2.96 3.77 3.475 ;
 RECT 4.55 2.11 4.69 2.8 ;
 RECT 1.75 3.535 1.89 3.58 ;
 RECT 1.75 2.96 1.89 3.395 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 3.72 1.96 3.745 ;
 RECT 2.05 3.11 2.32 3.25 ;
 RECT 1.555 3.885 1.96 4.04 ;
 RECT 1.555 3.745 2.255 3.885 ;
 RECT 2.115 3.25 2.255 3.745 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 5.44 5.2 ;
 RECT 2.07 4.26 2.49 4.665 ;
 RECT 2.215 4.665 2.355 5.04 ;
 RECT 1.745 4.3 1.885 5.04 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.6 1.475 3.745 1.615 ;
 RECT 2.765 0.89 2.905 1.475 ;
 RECT 2.765 1.81 2.905 2.29 ;
 RECT 2.6 1.615 2.92 1.81 ;
 RECT 3.605 0.955 3.745 1.475 ;
 END
 ANTENNADIFFAREA 0.522 ;
 END Q

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.795 1.14 5.27 1.42 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END ENB

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 2.29 0.08 2.43 1.385 ;
 RECT 0.47 0.08 0.61 1.275 ;
 RECT 1.395 0.08 1.535 1.02 ;
 RECT 3.135 0.08 3.275 1.325 ;
 RECT 4.075 0.08 4.215 1.325 ;
 RECT 4.985 0.08 5.125 0.87 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 5.44 5.84 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 1 2.535 1.1 3.06 ;
 RECT 1.15 1.865 1.25 2.435 ;
 RECT 1 2.435 1.25 2.535 ;
 RECT 0.93 3.06 1.16 3.29 ;
 RECT 1.53 3.17 1.63 3.785 ;
 RECT 1.53 3.785 1.83 4.015 ;
 RECT 1.53 4.015 1.63 4.73 ;
 RECT 1.15 0.23 1.25 1.29 ;
 RECT 2.55 0.23 2.65 1.595 ;
 RECT 2.2 1.595 2.65 1.825 ;
 RECT 2.55 1.825 2.65 2.7 ;
 RECT 1.15 0.13 2.65 0.23 ;
 RECT 1.65 2.4 2.145 2.5 ;
 RECT 2.045 2.5 2.145 3.065 ;
 RECT 2.045 3.065 2.3 3.295 ;
 RECT 1.65 1.84 1.75 2.4 ;
 RECT 1.455 1.165 1.75 1.395 ;
 RECT 1.65 0.47 1.75 1.165 ;
 RECT 4.805 1.4 4.905 2.52 ;
 RECT 4.77 0.445 4.87 1.175 ;
 RECT 4.77 1.175 5.235 1.4 ;
 RECT 3.86 1.485 3.985 1.615 ;
 RECT 3.885 1.615 3.985 3.73 ;
 RECT 3.86 0.505 3.96 1.485 ;
 RECT 3.39 1.49 3.515 1.615 ;
 RECT 3.415 1.615 3.515 3.73 ;
 RECT 3.39 0.505 3.49 1.49 ;
 RECT 4.36 0.29 4.59 0.405 ;
 RECT 3.39 0.405 4.59 0.505 ;
 RECT 4.23 2.665 4.33 2.865 ;
 RECT 4.42 2.965 4.52 3.155 ;
 RECT 4.165 2.43 4.395 2.665 ;
 RECT 4.355 3.155 4.585 3.385 ;
 RECT 4.23 2.865 4.52 2.965 ;
 LAYER CO ;
 RECT 1.28 3.4 1.41 3.53 ;
 RECT 2.77 1.995 2.9 2.125 ;
 RECT 0.98 3.11 1.11 3.24 ;
 RECT 0.475 0.565 0.605 0.695 ;
 RECT 1.75 4.37 1.88 4.5 ;
 RECT 1.87 0.815 2 0.945 ;
 RECT 2.465 3.185 2.595 3.315 ;
 RECT 0.9 2.09 1.03 2.22 ;
 RECT 2.225 4.3 2.355 4.43 ;
 RECT 2.25 1.645 2.38 1.775 ;
 RECT 2.77 1.125 2.9 1.255 ;
 RECT 2.465 3.445 2.595 3.575 ;
 RECT 1.4 2.09 1.53 2.22 ;
 RECT 2.745 3.445 2.875 3.575 ;
 RECT 1.65 3.835 1.78 3.965 ;
 RECT 2.12 3.115 2.25 3.245 ;
 RECT 5.025 2.16 5.155 2.29 ;
 RECT 4.555 2.16 4.685 2.29 ;
 RECT 4.99 0.685 5.12 0.815 ;
 RECT 4.52 0.685 4.65 0.815 ;
 RECT 0.475 1.085 0.605 1.215 ;
 RECT 4.405 3.205 4.535 3.335 ;
 RECT 4.105 2.09 4.235 2.22 ;
 RECT 3.165 2.09 3.295 2.22 ;
 RECT 3.635 2.16 3.765 2.29 ;
 RECT 3.165 3.295 3.295 3.425 ;
 RECT 4.105 3.295 4.235 3.425 ;
 RECT 3.635 3.295 3.765 3.425 ;
 RECT 4.08 1.125 4.21 1.255 ;
 RECT 4.08 0.815 4.21 0.945 ;
 RECT 3.61 1.125 3.74 1.255 ;
 RECT 3.14 0.815 3.27 0.945 ;
 RECT 3.14 1.125 3.27 1.255 ;
 RECT 3.61 1.125 3.74 1.255 ;
 RECT 1.28 4.36 1.41 4.49 ;
 RECT 0.475 0.825 0.605 0.955 ;
 RECT 1.87 2.09 2 2.22 ;
 RECT 2.29 1.99 2.42 2.12 ;
 RECT 2.745 3.185 2.875 3.315 ;
 RECT 1.4 0.83 1.53 0.96 ;
 RECT 1.755 3.4 1.885 3.53 ;
 RECT 1.505 1.215 1.635 1.345 ;
 RECT 2.295 1.125 2.425 1.255 ;
 RECT 0.9 0.835 1.03 0.965 ;
 RECT 5.055 1.215 5.185 1.345 ;
 RECT 4.41 0.33 4.54 0.46 ;
 RECT 4.215 2.47 4.345 2.6 ;
 LAYER M1 ;
 RECT 3.16 3.225 3.3 3.615 ;
 RECT 4.1 3.15 4.575 3.41 ;
 RECT 4.1 3.41 4.24 3.615 ;
 RECT 3.16 3.615 4.24 3.755 ;
 RECT 0.895 0.76 1.035 1.45 ;
 RECT 0.895 1.59 1.035 2.29 ;
 RECT 1.5 1.165 1.64 1.45 ;
 RECT 0.895 1.45 1.64 1.59 ;
 RECT 1.275 3.245 1.415 4.56 ;
 RECT 0.93 3.105 1.415 3.245 ;
 RECT 1.865 0.745 2.005 1.64 ;
 RECT 1.865 1.78 2.005 2.29 ;
 RECT 1.865 1.64 2.46 1.78 ;
 RECT 2.2 1.6 2.46 1.64 ;
 RECT 2.2 1.78 2.46 1.83 ;
 RECT 4.515 0.51 4.655 1.825 ;
 RECT 4.36 0.29 4.655 0.51 ;
 RECT 5.02 1.965 5.16 2.36 ;
 RECT 4.515 1.825 5.16 1.965 ;
 RECT 1.425 2.225 1.565 2.51 ;
 RECT 2.285 2.125 2.425 2.51 ;
 RECT 1.325 2.085 1.6 2.225 ;
 RECT 2.22 1.985 2.49 2.125 ;
 RECT 3.16 1.96 3.3 2.51 ;
 RECT 1.425 2.51 3.3 2.65 ;
 RECT 3.16 1.82 4.24 1.96 ;
 RECT 4.1 1.96 4.24 2.41 ;
 RECT 4.1 2.41 4.395 2.66 ;
 END
END LSUPENX1

MACRO LSUPENX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.72 BY 5.76 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.955 1.57 6 1.71 ;
 RECT 4.97 1.71 5.11 1.755 ;
 RECT 4.97 1.525 5.11 1.57 ;
 RECT 5.57 1.81 5.71 2.175 ;
 RECT 5.57 1.71 6 1.81 ;
 RECT 5.57 1.03 5.71 1.395 ;
 RECT 5.57 1.395 6 1.57 ;
 END
 ANTENNADIFFAREA 0.656 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.855 3.11 5.125 3.25 ;
 RECT 4.36 3.86 4.855 4.04 ;
 RECT 4.92 3.25 5.06 3.72 ;
 RECT 4.36 3.72 5.06 3.86 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.72 2.96 ;
 RECT 4.49 3.395 4.75 3.535 ;
 RECT 2.085 2.275 2.225 2.8 ;
 RECT 5.265 2.96 5.685 3.645 ;
 RECT 3.03 2.2 3.17 2.8 ;
 RECT 1.145 1.94 1.285 2.8 ;
 RECT 0.305 2.18 0.445 2.8 ;
 RECT 4.555 3.535 4.695 3.58 ;
 RECT 4.555 2.96 4.695 3.395 ;
 END
 END VSS

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.035 6.72 5.195 ;
 RECT 4.875 4.26 5.295 4.665 ;
 RECT 5.02 4.665 5.16 5.035 ;
 RECT 4.55 4.3 4.69 5.035 ;
 END
 END VDDL

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.455 1.14 1.735 1.42 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END ENB

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.83 0.08 ;
 RECT 6.14 0.08 6.28 1.315 ;
 RECT 4.17 0.08 4.31 1.02 ;
 RECT 0.75 0.08 0.89 1.025 ;
 RECT 5.095 0.08 5.235 1.385 ;
 RECT 3.03 0.08 3.17 1.13 ;
 RECT 2.08 0.08 2.22 1.315 ;
 RECT 1.71 0.08 1.85 0.98 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 6.72 5.84 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 4.43 0.49 4.53 1.175 ;
 RECT 4.33 1.175 4.56 1.405 ;
 RECT 3.8 2.475 4.055 2.575 ;
 RECT 3.8 2.575 3.9 3.105 ;
 RECT 3.955 1.87 4.055 2.475 ;
 RECT 3.735 3.105 3.965 3.335 ;
 RECT 4.85 2.545 4.95 3.065 ;
 RECT 4.455 1.87 4.555 2.445 ;
 RECT 4.85 3.065 5.105 3.295 ;
 RECT 4.455 2.445 4.95 2.545 ;
 RECT 4.335 3.175 4.435 3.785 ;
 RECT 4.335 3.785 4.635 4.015 ;
 RECT 4.335 4.015 4.435 4.73 ;
 RECT 4.925 1.525 5.155 1.585 ;
 RECT 4.925 1.685 5.155 1.755 ;
 RECT 3.355 1.22 3.77 1.585 ;
 RECT 3.355 1.585 5.155 1.685 ;
 RECT 2.34 0.23 2.44 1.51 ;
 RECT 2.34 0.13 2.915 0.23 ;
 RECT 2.815 0.23 2.915 2.725 ;
 RECT 2.34 1.74 2.44 2.63 ;
 RECT 1.4 1.78 1.5 2.63 ;
 RECT 1.87 1.775 1.97 2.63 ;
 RECT 1.4 2.63 2.44 2.73 ;
 RECT 2.15 1.51 2.44 1.74 ;
 RECT 5.355 0.225 5.455 0.79 ;
 RECT 5.355 0.89 5.455 2.7 ;
 RECT 5.355 0.79 5.935 0.89 ;
 RECT 5.835 0.89 5.935 2.7 ;
 RECT 3.955 0.225 4.055 1.29 ;
 RECT 3.955 0.13 5.455 0.225 ;
 RECT 3.955 0.125 5.45 0.13 ;
 RECT 4.72 0.225 4.95 0.43 ;
 RECT 0.56 1.36 0.66 2.58 ;
 RECT 0.56 1.26 1.7 1.36 ;
 RECT 1.47 1.175 1.7 1.26 ;
 RECT 1.47 1.36 1.7 1.385 ;
 RECT 1.495 0.555 1.595 1.175 ;
 LAYER CO ;
 RECT 3.035 0.91 3.165 1.04 ;
 RECT 2.085 0.815 2.215 0.945 ;
 RECT 2.56 1.125 2.69 1.255 ;
 RECT 2.085 1.125 2.215 1.255 ;
 RECT 3.035 0.545 3.165 0.675 ;
 RECT 2.56 0.815 2.69 0.945 ;
 RECT 0.31 2.23 0.44 2.36 ;
 RECT 0.78 2.23 0.91 2.36 ;
 RECT 1.245 0.795 1.375 0.925 ;
 RECT 1.715 0.795 1.845 0.925 ;
 RECT 2.225 1.56 2.355 1.69 ;
 RECT 1.15 2.01 1.28 2.14 ;
 RECT 1.15 2.27 1.28 2.4 ;
 RECT 4.38 1.225 4.51 1.355 ;
 RECT 4.56 3.4 4.69 3.53 ;
 RECT 4.085 4.36 4.215 4.49 ;
 RECT 5.55 3.445 5.68 3.575 ;
 RECT 4.65 0.815 4.78 0.945 ;
 RECT 4.975 1.575 5.105 1.705 ;
 RECT 0.755 0.825 0.885 0.955 ;
 RECT 4.175 0.83 4.305 0.96 ;
 RECT 5.575 1.985 5.705 2.115 ;
 RECT 3.705 0.835 3.835 0.965 ;
 RECT 0.755 0.565 0.885 0.695 ;
 RECT 5.095 1.985 5.225 2.115 ;
 RECT 3.785 3.15 3.915 3.28 ;
 RECT 4.205 2.09 4.335 2.22 ;
 RECT 4.925 3.115 5.055 3.245 ;
 RECT 4.085 3.4 4.215 3.53 ;
 RECT 4.455 3.835 4.585 3.965 ;
 RECT 5.55 3.185 5.68 3.315 ;
 RECT 4.555 4.37 4.685 4.5 ;
 RECT 5.575 1.125 5.705 1.255 ;
 RECT 5.03 4.3 5.16 4.43 ;
 RECT 5.27 3.185 5.4 3.315 ;
 RECT 5.1 1.125 5.23 1.255 ;
 RECT 3.705 2.09 3.835 2.22 ;
 RECT 4.675 2.09 4.805 2.22 ;
 RECT 5.27 3.445 5.4 3.575 ;
 RECT 6.145 1.985 6.275 2.115 ;
 RECT 6.145 1.125 6.275 1.255 ;
 RECT 3.42 1.275 3.55 1.405 ;
 RECT 2.09 2.35 2.22 2.48 ;
 RECT 1.62 2.085 1.75 2.215 ;
 RECT 1.62 2.35 1.75 2.48 ;
 RECT 2.56 2.35 2.69 2.48 ;
 RECT 3.035 2.27 3.165 2.4 ;
 RECT 2.56 2.085 2.69 2.215 ;
 RECT 4.77 0.26 4.9 0.39 ;
 RECT 1.52 1.215 1.65 1.345 ;
 LAYER M1 ;
 RECT 1.175 0.93 1.315 1.57 ;
 RECT 1.165 0.79 1.445 0.93 ;
 RECT 0.775 1.71 0.915 2.43 ;
 RECT 0.775 1.57 2.415 1.71 ;
 RECT 2.115 1.48 2.415 1.57 ;
 RECT 2.115 1.71 2.415 1.78 ;
 RECT 4.08 3.285 4.22 4.56 ;
 RECT 3.78 3.1 3.92 3.145 ;
 RECT 3.78 3.285 3.92 3.335 ;
 RECT 3.735 3.145 4.22 3.285 ;
 RECT 2.555 0.745 2.695 1.27 ;
 RECT 3.415 1.225 3.555 1.27 ;
 RECT 3.415 1.41 3.555 1.545 ;
 RECT 2.555 1.27 3.555 1.41 ;
 RECT 3.7 0.76 3.84 1.225 ;
 RECT 3.7 1.365 3.84 2.29 ;
 RECT 4.375 1.175 4.515 1.225 ;
 RECT 3.7 1.225 4.515 1.365 ;
 RECT 4.375 1.365 4.515 1.415 ;
 RECT 2.555 2.06 2.695 2.55 ;
 RECT 1.615 1.915 1.755 1.92 ;
 RECT 1.615 2.06 1.755 2.55 ;
 RECT 4.2 2.225 4.34 2.515 ;
 RECT 1.615 1.92 3.56 2.06 ;
 RECT 3.42 2.06 3.56 2.515 ;
 RECT 5.09 1.92 5.23 2.515 ;
 RECT 4.2 2.065 4.34 2.085 ;
 RECT 4.13 2.085 4.405 2.225 ;
 RECT 3.42 2.515 6.28 2.645 ;
 RECT 6.14 1.88 6.28 2.515 ;
 RECT 3.425 2.645 6.28 2.655 ;
 RECT 4.645 0.22 4.95 0.43 ;
 RECT 4.645 0.43 4.785 0.905 ;
 RECT 4.645 0.905 4.81 1.015 ;
 RECT 4.67 1.015 4.81 2.29 ;
 END
END LSUPENX2

MACRO LSUPENX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.68 BY 5.76 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.545 3.565 2.025 3.915 ;
 END
 ANTENNAGATEAREA 0.143 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 7.68 5.2 ;
 RECT 2.125 4.14 2.545 4.545 ;
 RECT 1.735 4.065 1.875 5.04 ;
 RECT 2.27 4.545 2.41 5.04 ;
 END
 END VDDL

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.02 1.49 7.325 1.795 ;
 END
 ANTENNAGATEAREA 0.092 ;
 END ENB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.68 2.96 ;
 RECT 3.5 2.96 3.92 3.645 ;
 RECT 7.21 1.995 7.35 2.8 ;
 RECT 1.74 2.96 1.88 3.35 ;
 RECT 5.425 2.135 5.565 2.8 ;
 RECT 4.485 2.135 4.625 2.8 ;
 RECT 6.37 2.135 6.51 2.8 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.7 1.795 2.84 2.285 ;
 RECT 2.7 0.74 2.84 1.46 ;
 RECT 3.64 1.6 3.78 2.305 ;
 RECT 3.64 0.74 3.78 1.46 ;
 RECT 4.955 0.74 5.095 1.46 ;
 RECT 2.7 1.6 3.13 1.795 ;
 RECT 2.7 1.46 5.1 1.6 ;
 END
 ANTENNADIFFAREA 1.708 ;
 END Q

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.68 0.08 ;
 RECT 7.215 0.08 7.355 1.31 ;
 RECT 2.225 0.08 2.365 1.3 ;
 RECT 1.3 0.08 1.44 1.11 ;
 RECT 3.17 0.08 3.31 1.3 ;
 RECT 0.405 0.08 0.545 1.27 ;
 RECT 4.11 0.08 4.25 1.3 ;
 RECT 4.485 0.08 4.625 1.32 ;
 RECT 5.425 0.08 5.565 1.32 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 7.68 5.84 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 1.52 2.895 1.62 3.585 ;
 RECT 1.52 3.585 1.82 3.815 ;
 RECT 1.52 3.815 1.62 4.575 ;
 RECT 1.585 1.885 1.685 2.78 ;
 RECT 1.52 2.78 1.685 2.895 ;
 RECT 1.085 0.11 3.995 0.21 ;
 RECT 1.085 0.21 1.185 1.49 ;
 RECT 2.485 0.21 2.585 1.46 ;
 RECT 1.85 1.46 2.585 1.695 ;
 RECT 2.485 1.695 2.585 2.74 ;
 RECT 3.895 0.21 3.995 2.74 ;
 RECT 3.425 0.21 3.525 2.745 ;
 RECT 2.955 0.21 3.055 2.74 ;
 RECT 6.995 0.75 7.095 1.545 ;
 RECT 6.995 1.545 7.25 1.755 ;
 RECT 6.995 1.755 7.095 2.605 ;
 RECT 0.8 2.805 0.9 3.1 ;
 RECT 1.085 1.875 1.185 2.705 ;
 RECT 0.8 2.705 1.185 2.805 ;
 RECT 0.74 3.1 0.97 3.31 ;
 RECT 1.395 1.495 1.655 1.705 ;
 RECT 1.555 0.495 1.655 1.495 ;
 RECT 5.685 1.64 5.785 2.655 ;
 RECT 5.21 0.125 5.31 1.54 ;
 RECT 5.21 1.64 5.31 2.655 ;
 RECT 4.74 0.125 4.84 1.54 ;
 RECT 4.74 1.64 4.84 2.66 ;
 RECT 4.74 1.54 6.31 1.64 ;
 RECT 6.08 1.5 6.31 1.54 ;
 RECT 6.08 1.64 6.31 1.71 ;
 RECT 6.155 1.71 6.255 2.655 ;
 LAYER CO ;
 RECT 3.785 3.445 3.915 3.575 ;
 RECT 1.745 3.14 1.875 3.27 ;
 RECT 1.805 2.245 1.935 2.375 ;
 RECT 4.96 2.04 5.09 2.17 ;
 RECT 3.505 3.445 3.635 3.575 ;
 RECT 3.175 0.81 3.305 0.94 ;
 RECT 4.96 1.12 5.09 1.25 ;
 RECT 1.305 0.91 1.435 1.04 ;
 RECT 3.645 2.085 3.775 2.215 ;
 RECT 4.125 2.085 4.255 2.215 ;
 RECT 4.115 1.12 4.245 1.25 ;
 RECT 3.645 1.12 3.775 1.25 ;
 RECT 4.115 0.81 4.245 0.94 ;
 RECT 3.645 0.81 3.775 0.94 ;
 RECT 4.49 1.12 4.62 1.25 ;
 RECT 4.49 0.81 4.62 0.94 ;
 RECT 5.43 2.235 5.56 2.365 ;
 RECT 3.785 3.185 3.915 3.315 ;
 RECT 3.505 3.185 3.635 3.315 ;
 RECT 5.43 0.81 5.56 0.94 ;
 RECT 0.41 1.08 0.54 1.21 ;
 RECT 2.705 2.085 2.835 2.215 ;
 RECT 2.705 0.81 2.835 0.94 ;
 RECT 3.175 2.085 3.305 2.215 ;
 RECT 0.835 1.1 0.965 1.23 ;
 RECT 4.96 0.81 5.09 0.94 ;
 RECT 2.23 0.81 2.36 0.94 ;
 RECT 4.49 2.215 4.62 2.345 ;
 RECT 4.96 1.12 5.09 1.25 ;
 RECT 0.41 0.82 0.54 0.95 ;
 RECT 0.41 0.56 0.54 0.69 ;
 RECT 2.28 4.25 2.41 4.38 ;
 RECT 2.705 1.12 2.835 1.25 ;
 RECT 1.335 2.235 1.465 2.365 ;
 RECT 1.775 1.1 1.905 1.23 ;
 RECT 1.64 3.635 1.77 3.765 ;
 RECT 4.96 0.81 5.09 0.94 ;
 RECT 0.835 2.235 0.965 2.365 ;
 RECT 3.175 1.12 3.305 1.25 ;
 RECT 6.745 2.035 6.875 2.165 ;
 RECT 7.215 2.1 7.345 2.23 ;
 RECT 6.745 1.165 6.875 1.295 ;
 RECT 7.22 1.11 7.35 1.24 ;
 RECT 6.375 2.235 6.505 2.365 ;
 RECT 5.905 2.14 6.035 2.27 ;
 RECT 1.27 3.195 1.4 3.325 ;
 RECT 1.27 4.005 1.4 4.135 ;
 RECT 2.225 2.085 2.355 2.215 ;
 RECT 5.43 1.12 5.56 1.25 ;
 RECT 2.23 1.12 2.36 1.25 ;
 RECT 1.74 4.14 1.87 4.27 ;
 RECT 1.9 1.525 2.03 1.655 ;
 RECT 7.07 1.585 7.2 1.715 ;
 RECT 0.79 3.14 0.92 3.27 ;
 RECT 1.445 1.535 1.575 1.665 ;
 RECT 6.13 1.54 6.26 1.67 ;
 LAYER M1 ;
 RECT 4.955 1.99 5.095 2.41 ;
 RECT 3.17 2.015 3.31 2.52 ;
 RECT 1.36 2.37 1.5 2.52 ;
 RECT 2.22 2.015 2.36 2.52 ;
 RECT 1.26 2.23 1.535 2.37 ;
 RECT 4.12 1.99 4.26 2.52 ;
 RECT 1.36 2.52 4.26 2.66 ;
 RECT 5.9 1.99 6.04 2.41 ;
 RECT 4.12 1.85 6.04 1.99 ;
 RECT 1.77 1.695 1.91 2.24 ;
 RECT 1.77 1.03 1.91 1.485 ;
 RECT 1.77 1.485 2.08 1.695 ;
 RECT 1.735 2.24 2.005 2.38 ;
 RECT 1.265 3.26 1.405 4.215 ;
 RECT 0.74 3.12 1.405 3.26 ;
 RECT 0.74 3.1 0.97 3.12 ;
 RECT 0.74 3.26 0.97 3.31 ;
 RECT 0.83 0.875 0.97 1.565 ;
 RECT 0.83 1.705 0.97 2.435 ;
 RECT 1.395 1.495 1.625 1.565 ;
 RECT 0.83 1.565 1.625 1.705 ;
 RECT 6.74 1.095 6.88 1.465 ;
 RECT 6.74 1.71 6.88 2.295 ;
 RECT 6.08 1.465 6.88 1.71 ;
 END
END LSUPENX4

MACRO LSUPENX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.92 BY 5.76 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.545 3.575 2.04 3.93 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 9.92 5.2 ;
 RECT 2.06 4.075 2.48 4.48 ;
 RECT 1.735 4.08 1.875 5.04 ;
 RECT 2.205 4.48 2.345 5.04 ;
 END
 END VDDL

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.92 2.96 ;
 RECT 3.915 2.96 4.335 3.655 ;
 RECT 1.74 2.96 1.88 3.4 ;
 RECT 9.375 1.96 9.515 2.8 ;
 RECT 7.365 2 7.505 2.8 ;
 RECT 6.425 2.005 6.565 2.8 ;
 RECT 8.305 1.995 8.445 2.8 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.75 1.785 2.89 2.215 ;
 RECT 2.745 1.58 3.18 1.785 ;
 RECT 2.75 0.72 2.89 1.44 ;
 RECT 4.63 1.58 4.77 2.285 ;
 RECT 3.69 1.58 3.83 2.215 ;
 RECT 5.57 1.58 5.71 2.285 ;
 RECT 2.745 1.56 7.03 1.58 ;
 RECT 2.745 1.45 7.035 1.56 ;
 RECT 4.63 0.72 4.77 1.44 ;
 RECT 3.69 0.72 3.83 1.44 ;
 RECT 5.57 0.72 5.71 1.44 ;
 RECT 6.895 0.715 7.035 1.44 ;
 RECT 2.75 1.44 7.035 1.45 ;
 END
 ANTENNADIFFAREA 2.984 ;
 END Q

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.92 0.08 ;
 RECT 0.455 0.08 0.595 1.26 ;
 RECT 3.22 0.08 3.36 1.3 ;
 RECT 2.275 0.08 2.415 1.3 ;
 RECT 5.1 0.08 5.24 1.3 ;
 RECT 1.38 0.08 1.52 0.915 ;
 RECT 6.04 0.08 6.18 1.3 ;
 RECT 9.38 0.08 9.52 1.235 ;
 RECT 4.16 0.08 4.3 1.3 ;
 RECT 7.365 0.08 7.505 1.295 ;
 RECT 6.425 0.08 6.565 1.295 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 9.92 5.84 ;
 END
 END VDDH

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.185 1.455 9.68 1.81 ;
 END
 ANTENNAGATEAREA 0.092 ;
 END ENB

 OBS
 LAYER PO ;
 RECT 9.16 0.575 9.26 1.495 ;
 RECT 9.16 1.495 9.46 1.725 ;
 RECT 9.16 1.725 9.26 2.7 ;
 RECT 1.52 2.83 1.62 3.615 ;
 RECT 1.52 3.615 1.82 3.845 ;
 RECT 1.52 3.845 1.62 4.865 ;
 RECT 1.635 1.71 1.735 2.71 ;
 RECT 1.52 2.71 1.735 2.83 ;
 RECT 1.135 0.09 5.925 0.19 ;
 RECT 2.535 1.585 2.635 2.735 ;
 RECT 1.135 0.19 1.235 1.265 ;
 RECT 2.535 0.19 2.635 1.485 ;
 RECT 1.935 1.49 2.635 1.585 ;
 RECT 1.935 1.585 2.165 1.7 ;
 RECT 2.07 1.485 2.635 1.49 ;
 RECT 5.825 0.19 5.925 2.745 ;
 RECT 5.355 0.19 5.455 2.745 ;
 RECT 4.885 0.19 4.985 2.745 ;
 RECT 4.415 0.19 4.515 2.745 ;
 RECT 3.945 0.19 4.045 2.745 ;
 RECT 3.475 0.19 3.575 2.745 ;
 RECT 3.005 0.19 3.105 2.73 ;
 RECT 1.48 1.31 1.735 1.435 ;
 RECT 1.48 1.435 1.71 1.52 ;
 RECT 1.635 0.385 1.735 1.31 ;
 RECT 8.09 1.475 8.42 1.515 ;
 RECT 8.09 1.615 8.42 1.685 ;
 RECT 6.68 1.515 8.42 1.615 ;
 RECT 6.68 0.1 6.78 1.515 ;
 RECT 6.68 1.615 6.78 2.71 ;
 RECT 7.62 0.1 7.72 1.515 ;
 RECT 7.62 1.615 7.72 2.71 ;
 RECT 7.15 0.1 7.25 1.515 ;
 RECT 7.15 1.615 7.25 2.71 ;
 RECT 8.09 0.1 8.19 1.475 ;
 RECT 8.09 1.685 8.19 2.71 ;
 RECT 0.725 2.795 0.825 3.13 ;
 RECT 1.135 1.71 1.235 2.695 ;
 RECT 0.725 2.695 1.235 2.795 ;
 RECT 0.665 3.13 0.895 3.34 ;
 LAYER CO ;
 RECT 2.28 1.1 2.41 1.23 ;
 RECT 3.225 0.79 3.355 0.92 ;
 RECT 4.165 0.79 4.295 0.92 ;
 RECT 9.28 1.54 9.41 1.67 ;
 RECT 8.91 2.025 9.04 2.155 ;
 RECT 8.91 1.035 9.04 1.165 ;
 RECT 9.385 1.035 9.515 1.165 ;
 RECT 9.38 2.145 9.51 2.275 ;
 RECT 8.31 2.075 8.44 2.205 ;
 RECT 7.84 2.075 7.97 2.205 ;
 RECT 5.575 1.1 5.705 1.23 ;
 RECT 6.045 1.1 6.175 1.23 ;
 RECT 5.575 2.015 5.705 2.145 ;
 RECT 6.045 2.015 6.175 2.145 ;
 RECT 6.045 0.79 6.175 0.92 ;
 RECT 5.575 0.79 5.705 0.92 ;
 RECT 1.74 4.265 1.87 4.395 ;
 RECT 3.92 3.195 4.05 3.325 ;
 RECT 7.37 2.075 7.5 2.205 ;
 RECT 3.695 0.79 3.825 0.92 ;
 RECT 4.165 1.1 4.295 1.23 ;
 RECT 6.9 0.785 7.03 0.915 ;
 RECT 2.755 0.79 2.885 0.92 ;
 RECT 2.28 0.79 2.41 0.92 ;
 RECT 1.385 2.065 1.515 2.195 ;
 RECT 2.215 4.165 2.345 4.295 ;
 RECT 6.9 2.07 7.03 2.2 ;
 RECT 6.9 0.785 7.03 0.915 ;
 RECT 1.385 0.715 1.515 0.845 ;
 RECT 1.27 3.2 1.4 3.33 ;
 RECT 3.92 3.455 4.05 3.585 ;
 RECT 0.46 1.06 0.59 1.19 ;
 RECT 2.755 2.015 2.885 2.145 ;
 RECT 7.37 0.785 7.5 0.915 ;
 RECT 6.9 1.095 7.03 1.225 ;
 RECT 4.2 3.195 4.33 3.325 ;
 RECT 1.745 3.2 1.875 3.33 ;
 RECT 6.43 2.075 6.56 2.205 ;
 RECT 2.755 1.1 2.885 1.23 ;
 RECT 0.46 0.54 0.59 0.67 ;
 RECT 6.43 0.785 6.56 0.915 ;
 RECT 4.2 3.455 4.33 3.585 ;
 RECT 4.165 2.015 4.295 2.145 ;
 RECT 3.225 2.015 3.355 2.145 ;
 RECT 0.885 2.065 1.015 2.195 ;
 RECT 1.64 3.66 1.77 3.79 ;
 RECT 1.27 4.145 1.4 4.275 ;
 RECT 0.46 0.8 0.59 0.93 ;
 RECT 5.105 1.1 5.235 1.23 ;
 RECT 2.275 2.015 2.405 2.145 ;
 RECT 1.855 2.065 1.985 2.195 ;
 RECT 1.855 0.905 1.985 1.035 ;
 RECT 5.105 0.79 5.235 0.92 ;
 RECT 4.635 1.1 4.765 1.23 ;
 RECT 3.225 1.1 3.355 1.23 ;
 RECT 4.635 2.015 4.765 2.145 ;
 RECT 6.43 1.095 6.56 1.225 ;
 RECT 7.37 1.095 7.5 1.225 ;
 RECT 1.985 1.53 2.115 1.66 ;
 RECT 1.53 1.35 1.66 1.48 ;
 RECT 8.24 1.515 8.37 1.645 ;
 RECT 0.715 3.17 0.845 3.3 ;
 RECT 6.9 2.07 7.03 2.2 ;
 RECT 3.695 1.1 3.825 1.23 ;
 RECT 3.695 2.015 3.825 2.145 ;
 RECT 5.105 2.015 5.235 2.145 ;
 RECT 0.885 0.905 1.015 1.035 ;
 RECT 6.9 1.095 7.03 1.225 ;
 RECT 4.635 0.79 4.765 0.92 ;
 LAYER M1 ;
 RECT 5.1 1.945 5.24 2.505 ;
 RECT 4.16 1.945 4.3 2.505 ;
 RECT 3.22 1.945 3.36 2.505 ;
 RECT 1.41 2.2 1.55 2.505 ;
 RECT 2.27 1.945 2.41 2.505 ;
 RECT 1.31 2.06 1.585 2.2 ;
 RECT 6.895 1.86 7.035 2.33 ;
 RECT 6.04 1.86 6.18 2.505 ;
 RECT 1.41 2.505 6.18 2.645 ;
 RECT 7.835 1.86 7.975 2.33 ;
 RECT 6.04 1.72 7.975 1.86 ;
 RECT 1.85 0.835 1.99 1.49 ;
 RECT 1.85 1.49 2.165 1.7 ;
 RECT 1.85 1.7 1.99 2.265 ;
 RECT 0.88 0.835 1.02 1.425 ;
 RECT 0.88 1.565 1.02 2.265 ;
 RECT 0.88 1.425 1.71 1.565 ;
 RECT 1.48 1.31 1.71 1.425 ;
 RECT 8.905 0.93 9.045 1.465 ;
 RECT 8.905 1.695 9.045 2.23 ;
 RECT 8.12 1.465 9.045 1.695 ;
 RECT 1.265 3.125 1.405 3.13 ;
 RECT 1.265 3.27 1.405 4.345 ;
 RECT 0.665 3.27 0.895 3.34 ;
 RECT 0.665 3.13 1.405 3.27 ;
 END
END LSUPENX8

MACRO LSUPX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 5.76 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 3.86 2.05 4.04 ;
 RECT 2.05 3.11 2.32 3.25 ;
 RECT 1.555 3.72 2.255 3.86 ;
 RECT 2.115 3.25 2.255 3.72 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 3.84 5.2 ;
 RECT 2.07 4.26 2.49 4.665 ;
 RECT 2.215 4.665 2.355 5.04 ;
 RECT 1.745 4.3 1.885 5.04 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.765 1.395 3.195 1.81 ;
 RECT 2.765 0.745 2.905 1.395 ;
 RECT 2.765 1.81 2.905 2.29 ;
 END
 ANTENNADIFFAREA 0.49 ;
 END Q

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 1.395 0.08 1.535 1.02 ;
 RECT 0.47 0.08 0.61 1.025 ;
 RECT 2.29 0.08 2.43 1.385 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 3.84 5.84 ;
 END
 END VDDH

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 RECT 1.685 3.42 1.945 3.56 ;
 RECT 1.325 2.085 1.6 2.225 ;
 RECT 2.46 2.96 2.88 3.645 ;
 RECT 2.285 2.02 2.425 2.8 ;
 RECT 1.75 2.96 1.89 3.42 ;
 RECT 1.425 2.225 1.565 2.8 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 1.15 1.865 1.25 3.06 ;
 RECT 1.12 3.06 1.35 3.29 ;
 RECT 1.455 1.165 1.75 1.395 ;
 RECT 1.65 0.47 1.75 1.165 ;
 RECT 1.53 3.2 1.63 3.785 ;
 RECT 1.53 3.785 1.83 4.015 ;
 RECT 1.53 4.015 1.63 4.73 ;
 RECT 2.045 3.065 2.3 3.295 ;
 RECT 2.045 2.5 2.145 3.065 ;
 RECT 1.65 2.4 2.145 2.5 ;
 RECT 1.65 1.84 1.75 2.4 ;
 RECT 2.55 0.23 2.65 1.595 ;
 RECT 2.55 1.825 2.65 2.7 ;
 RECT 2.36 1.595 2.65 1.825 ;
 RECT 1.15 0.23 1.25 1.29 ;
 RECT 1.15 0.13 2.65 0.23 ;
 LAYER CO ;
 RECT 2.745 3.185 2.875 3.315 ;
 RECT 2.745 3.445 2.875 3.575 ;
 RECT 2.12 3.115 2.25 3.245 ;
 RECT 1.17 3.11 1.3 3.24 ;
 RECT 1.87 0.815 2 0.945 ;
 RECT 2.29 2.09 2.42 2.22 ;
 RECT 1.4 0.83 1.53 0.96 ;
 RECT 0.475 0.565 0.605 0.695 ;
 RECT 2.295 0.815 2.425 0.945 ;
 RECT 1.87 2.09 2 2.22 ;
 RECT 0.475 0.825 0.605 0.955 ;
 RECT 1.4 2.09 1.53 2.22 ;
 RECT 0.9 2.09 1.03 2.22 ;
 RECT 0.9 0.835 1.03 0.965 ;
 RECT 2.77 2.09 2.9 2.22 ;
 RECT 2.41 1.645 2.54 1.775 ;
 RECT 1.505 1.215 1.635 1.345 ;
 RECT 2.77 1.125 2.9 1.255 ;
 RECT 2.77 0.815 2.9 0.945 ;
 RECT 2.295 1.125 2.425 1.255 ;
 RECT 2.225 4.3 2.355 4.43 ;
 RECT 1.755 3.425 1.885 3.555 ;
 RECT 1.75 4.37 1.88 4.5 ;
 RECT 1.65 3.835 1.78 3.965 ;
 RECT 1.28 4.36 1.41 4.49 ;
 RECT 1.28 3.425 1.41 3.555 ;
 RECT 2.465 3.185 2.595 3.315 ;
 RECT 2.465 3.445 2.595 3.575 ;
 LAYER M1 ;
 RECT 1.865 0.745 2.005 1.64 ;
 RECT 1.865 1.78 2.005 2.29 ;
 RECT 1.865 1.64 2.59 1.78 ;
 RECT 0.895 0.76 1.035 1.45 ;
 RECT 0.895 1.59 1.035 2.29 ;
 RECT 1.5 1.165 1.64 1.45 ;
 RECT 0.895 1.45 1.64 1.59 ;
 RECT 1.275 3.245 1.415 4.56 ;
 RECT 1.1 3.105 1.415 3.245 ;
 END
END LSUPX1

MACRO LSUPX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 5.76 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 RECT 1.685 3.44 1.945 3.58 ;
 RECT 1.325 2.085 1.6 2.225 ;
 RECT 2.46 2.96 2.88 3.645 ;
 RECT 2.285 2.02 2.425 2.8 ;
 RECT 3.245 2.02 3.385 2.8 ;
 RECT 1.75 2.96 1.89 3.44 ;
 RECT 1.425 2.225 1.565 2.8 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 3.86 2.05 4.04 ;
 RECT 2.05 3.11 2.32 3.25 ;
 RECT 1.555 3.72 2.255 3.86 ;
 RECT 2.115 3.25 2.255 3.72 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 3.84 5.2 ;
 RECT 2.07 4.26 2.49 4.665 ;
 RECT 2.215 4.665 2.355 5.04 ;
 RECT 1.745 4.3 1.885 5.04 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.765 1.395 3.195 1.81 ;
 RECT 2.765 0.745 2.905 1.395 ;
 RECT 2.765 1.81 2.905 2.29 ;
 END
 ANTENNADIFFAREA 0.618 ;
 END Q

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 1.395 0.08 1.535 1.02 ;
 RECT 0.47 0.08 0.61 1.025 ;
 RECT 2.29 0.08 2.43 1.385 ;
 RECT 3.24 0.08 3.38 1.205 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 3.84 5.84 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 1.15 1.865 1.25 3.06 ;
 RECT 1.085 3.06 1.315 3.29 ;
 RECT 1.15 0.23 1.25 1.29 ;
 RECT 2.55 0.23 2.65 1.595 ;
 RECT 3.02 0.23 3.12 2.7 ;
 RECT 2.36 1.595 2.65 1.825 ;
 RECT 2.55 1.825 2.65 2.7 ;
 RECT 1.15 0.13 3.12 0.23 ;
 RECT 1.455 1.165 1.75 1.395 ;
 RECT 1.65 0.47 1.75 1.165 ;
 RECT 1.53 3.225 1.63 3.785 ;
 RECT 1.53 3.785 1.83 4.015 ;
 RECT 1.53 4.015 1.63 4.73 ;
 RECT 2.045 3.065 2.3 3.295 ;
 RECT 2.045 2.5 2.145 3.065 ;
 RECT 1.65 2.4 2.145 2.5 ;
 RECT 1.65 1.84 1.75 2.4 ;
 LAYER CO ;
 RECT 3.25 2.09 3.38 2.22 ;
 RECT 3.245 0.91 3.375 1.04 ;
 RECT 3.245 0.545 3.375 0.675 ;
 RECT 2.745 3.185 2.875 3.315 ;
 RECT 2.745 3.445 2.875 3.575 ;
 RECT 2.12 3.115 2.25 3.245 ;
 RECT 1.135 3.11 1.265 3.24 ;
 RECT 1.87 0.815 2 0.945 ;
 RECT 2.29 2.09 2.42 2.22 ;
 RECT 1.4 0.83 1.53 0.96 ;
 RECT 0.475 0.565 0.605 0.695 ;
 RECT 2.295 0.815 2.425 0.945 ;
 RECT 1.87 2.09 2 2.22 ;
 RECT 0.475 0.825 0.605 0.955 ;
 RECT 1.4 2.09 1.53 2.22 ;
 RECT 0.9 2.09 1.03 2.22 ;
 RECT 0.9 0.835 1.03 0.965 ;
 RECT 2.77 2.09 2.9 2.22 ;
 RECT 2.41 1.645 2.54 1.775 ;
 RECT 1.505 1.215 1.635 1.345 ;
 RECT 2.77 1.125 2.9 1.255 ;
 RECT 2.77 0.815 2.9 0.945 ;
 RECT 2.295 1.125 2.425 1.255 ;
 RECT 2.225 4.3 2.355 4.43 ;
 RECT 1.755 3.445 1.885 3.575 ;
 RECT 1.75 4.37 1.88 4.5 ;
 RECT 1.65 3.835 1.78 3.965 ;
 RECT 1.28 4.36 1.41 4.49 ;
 RECT 1.28 3.445 1.41 3.575 ;
 RECT 2.465 3.185 2.595 3.315 ;
 RECT 2.465 3.445 2.595 3.575 ;
 LAYER M1 ;
 RECT 1.865 0.745 2.005 1.64 ;
 RECT 1.865 1.78 2.005 2.29 ;
 RECT 1.865 1.64 2.59 1.78 ;
 RECT 0.895 0.76 1.035 1.45 ;
 RECT 0.895 1.59 1.035 2.29 ;
 RECT 1.5 1.165 1.64 1.45 ;
 RECT 0.895 1.45 1.64 1.59 ;
 RECT 1.275 3.245 1.415 4.56 ;
 RECT 1.065 3.105 1.415 3.245 ;
 END
END LSUPX2

MACRO LSUPX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 5.76 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 1.685 3.44 1.945 3.58 ;
 RECT 1.325 2.085 1.6 2.225 ;
 RECT 2.46 2.96 2.88 3.645 ;
 RECT 2.285 2.02 2.425 2.8 ;
 RECT 3.245 2.02 3.385 2.8 ;
 RECT 4.195 2.02 4.335 2.8 ;
 RECT 1.75 2.96 1.89 3.44 ;
 RECT 1.425 2.225 1.565 2.8 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 3.86 2.05 4.04 ;
 RECT 2.05 3.11 2.32 3.25 ;
 RECT 1.555 3.72 2.255 3.86 ;
 RECT 2.115 3.25 2.255 3.72 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 4.48 5.2 ;
 RECT 2.07 4.26 2.49 4.665 ;
 RECT 2.215 4.665 2.355 5.04 ;
 RECT 1.745 4.3 1.885 5.04 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.765 1.81 2.905 2.29 ;
 RECT 2.765 0.745 2.905 1.395 ;
 RECT 2.765 1.64 3.855 1.78 ;
 RECT 2.765 1.78 3.195 1.81 ;
 RECT 2.765 1.395 3.195 1.64 ;
 RECT 3.715 1.78 3.855 2.29 ;
 RECT 3.715 0.745 3.855 1.64 ;
 END
 ANTENNADIFFAREA 1.236 ;
 END Q

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 1.395 0.08 1.535 1.02 ;
 RECT 0.47 0.08 0.61 1.025 ;
 RECT 2.29 0.08 2.43 1.385 ;
 RECT 3.24 0.08 3.38 1.205 ;
 RECT 4.19 0.08 4.33 1.205 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 4.48 5.84 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 1.15 1.865 1.25 3.06 ;
 RECT 1.115 3.06 1.345 3.29 ;
 RECT 3.02 0.23 3.12 1.62 ;
 RECT 3.02 1.62 4.07 1.72 ;
 RECT 3.02 1.72 3.12 2.7 ;
 RECT 3.97 0.13 4.07 1.62 ;
 RECT 3.97 1.72 4.07 2.7 ;
 RECT 3.5 0.13 3.6 1.62 ;
 RECT 3.5 1.72 3.6 2.7 ;
 RECT 1.15 0.23 1.25 1.29 ;
 RECT 2.55 0.23 2.65 1.595 ;
 RECT 2.36 1.595 2.65 1.825 ;
 RECT 2.55 1.825 2.65 2.7 ;
 RECT 1.15 0.13 3.12 0.23 ;
 RECT 1.455 1.165 1.75 1.395 ;
 RECT 1.65 0.47 1.75 1.165 ;
 RECT 1.53 3.22 1.63 3.785 ;
 RECT 1.53 3.785 1.83 4.015 ;
 RECT 1.53 4.015 1.63 4.73 ;
 RECT 2.045 3.065 2.3 3.295 ;
 RECT 2.045 2.5 2.145 3.065 ;
 RECT 1.65 2.4 2.145 2.5 ;
 RECT 1.65 1.84 1.75 2.4 ;
 LAYER CO ;
 RECT 3.72 0.815 3.85 0.945 ;
 RECT 4.195 0.545 4.325 0.675 ;
 RECT 3.72 2.09 3.85 2.22 ;
 RECT 4.2 2.09 4.33 2.22 ;
 RECT 3.72 1.125 3.85 1.255 ;
 RECT 3.25 2.09 3.38 2.22 ;
 RECT 3.245 0.91 3.375 1.04 ;
 RECT 3.245 0.545 3.375 0.675 ;
 RECT 2.745 3.185 2.875 3.315 ;
 RECT 2.745 3.445 2.875 3.575 ;
 RECT 2.12 3.115 2.25 3.245 ;
 RECT 1.165 3.11 1.295 3.24 ;
 RECT 1.87 0.815 2 0.945 ;
 RECT 2.29 2.09 2.42 2.22 ;
 RECT 1.4 0.83 1.53 0.96 ;
 RECT 0.475 0.565 0.605 0.695 ;
 RECT 2.295 0.815 2.425 0.945 ;
 RECT 1.87 2.09 2 2.22 ;
 RECT 0.475 0.825 0.605 0.955 ;
 RECT 1.4 2.09 1.53 2.22 ;
 RECT 0.9 2.09 1.03 2.22 ;
 RECT 0.9 0.835 1.03 0.965 ;
 RECT 2.77 2.09 2.9 2.22 ;
 RECT 2.41 1.645 2.54 1.775 ;
 RECT 1.505 1.215 1.635 1.345 ;
 RECT 2.77 1.125 2.9 1.255 ;
 RECT 2.77 0.815 2.9 0.945 ;
 RECT 2.295 1.125 2.425 1.255 ;
 RECT 2.225 4.3 2.355 4.43 ;
 RECT 1.755 3.445 1.885 3.575 ;
 RECT 1.75 4.37 1.88 4.5 ;
 RECT 1.65 3.835 1.78 3.965 ;
 RECT 1.28 4.36 1.41 4.49 ;
 RECT 1.28 3.445 1.41 3.575 ;
 RECT 2.465 3.185 2.595 3.315 ;
 RECT 2.465 3.445 2.595 3.575 ;
 RECT 4.195 0.91 4.325 1.04 ;
 LAYER M1 ;
 RECT 1.865 0.745 2.005 1.64 ;
 RECT 1.865 1.78 2.005 2.29 ;
 RECT 1.865 1.64 2.59 1.78 ;
 RECT 0.895 0.76 1.035 1.45 ;
 RECT 0.895 1.59 1.035 2.29 ;
 RECT 1.5 1.165 1.64 1.45 ;
 RECT 0.895 1.45 1.64 1.59 ;
 RECT 1.275 3.245 1.415 4.56 ;
 RECT 1.095 3.105 1.415 3.245 ;
 END
END LSUPX4

MACRO LSUPX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.4 BY 5.76 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.4 2.96 ;
 RECT 1.685 3.415 1.945 3.555 ;
 RECT 1.325 2.085 1.6 2.225 ;
 RECT 2.46 2.96 2.88 3.645 ;
 RECT 2.285 2.02 2.425 2.8 ;
 RECT 3.245 2.02 3.385 2.8 ;
 RECT 5.14 2.02 5.28 2.8 ;
 RECT 6.09 2.02 6.23 2.8 ;
 RECT 4.19 2.02 4.33 2.8 ;
 RECT 1.75 2.96 1.89 3.415 ;
 RECT 1.425 2.225 1.565 2.8 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.05 3.11 2.32 3.25 ;
 RECT 1.555 3.835 2.05 4.04 ;
 RECT 2.115 3.25 2.255 3.695 ;
 RECT 1.555 3.695 2.255 3.835 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 6.4 5.2 ;
 RECT 2.07 4.26 2.49 4.665 ;
 RECT 2.215 4.665 2.355 5.04 ;
 RECT 1.745 4.3 1.885 5.04 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.765 1.81 2.905 2.29 ;
 RECT 2.765 0.745 2.905 1.395 ;
 RECT 2.765 1.78 3.195 1.81 ;
 RECT 2.765 1.395 3.195 1.64 ;
 RECT 3.715 1.78 3.855 2.29 ;
 RECT 3.715 0.745 3.855 1.64 ;
 RECT 4.66 1.78 4.8 2.29 ;
 RECT 4.66 0.745 4.8 1.64 ;
 RECT 5.61 1.78 5.75 2.29 ;
 RECT 5.61 0.745 5.75 1.64 ;
 RECT 2.765 1.64 5.75 1.78 ;
 END
 ANTENNADIFFAREA 2.472 ;
 END Q

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.4 0.08 ;
 RECT 1.395 0.08 1.535 1.02 ;
 RECT 0.47 0.08 0.61 1.025 ;
 RECT 2.29 0.08 2.43 1.385 ;
 RECT 3.24 0.08 3.38 1.205 ;
 RECT 4.19 0.08 4.33 1.205 ;
 RECT 5.135 0.08 5.275 1.205 ;
 RECT 6.085 0.08 6.225 1.205 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 6.4 5.84 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 1.15 1.865 1.25 3.055 ;
 RECT 1.115 3.055 1.345 3.285 ;
 RECT 1.455 1.165 1.75 1.395 ;
 RECT 1.65 0.47 1.75 1.165 ;
 RECT 1.53 3.195 1.63 3.785 ;
 RECT 1.53 3.785 1.83 4.015 ;
 RECT 1.53 4.015 1.63 4.73 ;
 RECT 2.045 3.065 2.3 3.295 ;
 RECT 2.045 2.5 2.145 3.065 ;
 RECT 1.65 2.4 2.145 2.5 ;
 RECT 1.65 1.84 1.75 2.4 ;
 RECT 3.02 1.62 5.965 1.72 ;
 RECT 2.55 0.23 2.65 1.595 ;
 RECT 2.36 1.595 2.65 1.825 ;
 RECT 2.55 1.825 2.65 2.7 ;
 RECT 1.15 0.23 1.25 1.29 ;
 RECT 3.02 0.23 3.12 1.62 ;
 RECT 3.5 0.13 3.6 1.62 ;
 RECT 3.5 1.72 3.6 2.7 ;
 RECT 3.02 1.72 3.12 2.7 ;
 RECT 3.97 0.13 4.07 1.62 ;
 RECT 3.97 1.72 4.07 2.7 ;
 RECT 5.865 0.13 5.965 1.62 ;
 RECT 5.865 1.72 5.965 2.7 ;
 RECT 5.395 0.13 5.495 1.62 ;
 RECT 5.395 1.72 5.495 2.7 ;
 RECT 4.915 0.13 5.015 1.62 ;
 RECT 4.915 1.72 5.015 2.7 ;
 RECT 4.445 0.13 4.545 1.62 ;
 RECT 4.445 1.72 4.545 2.7 ;
 RECT 1.15 0.13 3.12 0.23 ;
 LAYER CO ;
 RECT 3.72 2.09 3.85 2.22 ;
 RECT 3.72 1.125 3.85 1.255 ;
 RECT 3.25 2.09 3.38 2.22 ;
 RECT 3.245 0.91 3.375 1.04 ;
 RECT 3.245 0.545 3.375 0.675 ;
 RECT 2.745 3.185 2.875 3.315 ;
 RECT 2.745 3.445 2.875 3.575 ;
 RECT 2.12 3.115 2.25 3.245 ;
 RECT 1.165 3.105 1.295 3.235 ;
 RECT 1.87 0.815 2 0.945 ;
 RECT 2.29 2.09 2.42 2.22 ;
 RECT 1.4 0.83 1.53 0.96 ;
 RECT 0.475 0.565 0.605 0.695 ;
 RECT 2.295 0.815 2.425 0.945 ;
 RECT 1.87 2.09 2 2.22 ;
 RECT 0.475 0.825 0.605 0.955 ;
 RECT 1.4 2.09 1.53 2.22 ;
 RECT 0.9 2.09 1.03 2.22 ;
 RECT 0.9 0.835 1.03 0.965 ;
 RECT 2.77 2.09 2.9 2.22 ;
 RECT 2.41 1.645 2.54 1.775 ;
 RECT 1.505 1.215 1.635 1.345 ;
 RECT 2.77 1.125 2.9 1.255 ;
 RECT 2.77 0.815 2.9 0.945 ;
 RECT 2.295 1.125 2.425 1.255 ;
 RECT 2.225 4.3 2.355 4.43 ;
 RECT 1.755 3.42 1.885 3.55 ;
 RECT 1.75 4.37 1.88 4.5 ;
 RECT 1.65 3.835 1.78 3.965 ;
 RECT 1.28 4.36 1.41 4.49 ;
 RECT 1.28 3.425 1.41 3.555 ;
 RECT 2.465 3.185 2.595 3.315 ;
 RECT 2.465 3.445 2.595 3.575 ;
 RECT 5.14 0.91 5.27 1.04 ;
 RECT 4.665 0.815 4.795 0.945 ;
 RECT 5.14 0.545 5.27 0.675 ;
 RECT 4.195 2.09 4.325 2.22 ;
 RECT 5.615 2.09 5.745 2.22 ;
 RECT 6.09 0.91 6.22 1.04 ;
 RECT 6.095 2.09 6.225 2.22 ;
 RECT 5.615 0.815 5.745 0.945 ;
 RECT 5.615 1.125 5.745 1.255 ;
 RECT 6.09 0.545 6.22 0.675 ;
 RECT 4.195 0.955 4.325 1.085 ;
 RECT 4.665 2.09 4.795 2.22 ;
 RECT 5.145 2.09 5.275 2.22 ;
 RECT 4.665 1.125 4.795 1.255 ;
 RECT 3.72 0.815 3.85 0.945 ;
 RECT 4.195 0.545 4.325 0.675 ;
 LAYER M1 ;
 RECT 1.865 0.745 2.005 1.64 ;
 RECT 1.865 1.78 2.005 2.29 ;
 RECT 1.865 1.64 2.59 1.78 ;
 RECT 0.895 0.76 1.035 1.45 ;
 RECT 0.895 1.59 1.035 2.29 ;
 RECT 1.5 1.165 1.64 1.45 ;
 RECT 0.895 1.45 1.64 1.59 ;
 RECT 1.095 3.105 1.415 3.24 ;
 RECT 1.275 3.24 1.415 4.56 ;
 RECT 1.095 3.1 1.405 3.105 ;
 END
END LSUPX8

MACRO RDFFNSRARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 26.88 BY 2.88 ;
 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.01 0.735 5.13 0.875 ;
 RECT 7.145 0.85 8.005 0.99 ;
 RECT 9.875 1.09 12.245 1.23 ;
 RECT 4.01 0.485 4.25 0.735 ;
 RECT 4.99 0.36 5.13 0.735 ;
 RECT 12.105 0.81 12.245 1.09 ;
 RECT 12.105 0.6 12.395 0.81 ;
 RECT 7.145 0.36 7.285 0.85 ;
 RECT 4.99 0.22 7.285 0.36 ;
 RECT 7.865 0.385 8.005 0.85 ;
 RECT 9.875 0.385 10.015 1.09 ;
 RECT 7.865 0.245 10.01 0.255 ;
 RECT 7.865 0.255 10.015 0.385 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 26.88 0.08 ;
 RECT 23.7 0.08 23.94 0.26 ;
 RECT 15.105 0.335 15.37 0.495 ;
 RECT 7.425 0.57 7.695 0.71 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 4.615 0.08 4.85 0.595 ;
 RECT 21.35 0.08 21.49 0.36 ;
 RECT 11.35 0.08 11.49 0.945 ;
 RECT 12.855 0.08 12.995 0.525 ;
 RECT 22.565 0.08 22.705 0.35 ;
 RECT 2.015 0.08 2.155 0.39 ;
 RECT 17.625 0.08 17.765 0.82 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 15.16 0.08 15.3 0.335 ;
 RECT 7.49 0.08 7.63 0.57 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 26.88 2.96 ;
 RECT 1.945 2.34 2.195 2.8 ;
 RECT 15.075 2.57 15.215 2.8 ;
 RECT 17.54 2.57 17.68 2.8 ;
 RECT 11.95 2.57 12.09 2.8 ;
 RECT 12.85 2.57 12.99 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.27 1.98 1.41 2.8 ;
 RECT 7.3 2.375 7.44 2.8 ;
 RECT 5.2 2.07 5.34 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.475 1.65 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.765 0.22 1.13 0.615 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.465 1.205 14.82 1.445 ;
 RECT 14.67 0.915 14.81 1.205 ;
 RECT 14.67 1.7 15.815 1.84 ;
 RECT 14.67 1.84 14.81 1.885 ;
 RECT 14.67 1.445 14.81 1.7 ;
 RECT 15.675 1.84 15.815 1.885 ;
 RECT 15.675 0.915 15.815 1.7 ;
 END
 ANTENNADIFFAREA 0.774 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 16.945 1.095 17.205 1.335 ;
 RECT 17.065 0.51 17.205 1.095 ;
 RECT 18.125 1.905 18.265 1.91 ;
 RECT 17.065 1.765 18.265 1.905 ;
 RECT 18.125 0.56 18.265 1.765 ;
 RECT 17.065 1.905 17.205 1.915 ;
 RECT 17.065 1.335 17.205 1.765 ;
 END
 ANTENNADIFFAREA 0.632 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.88 1.135 7.27 1.49 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 25.26 1.435 25.6 1.8 ;
 RECT 23.58 1.99 25.445 2.13 ;
 RECT 21.35 2.22 23.72 2.36 ;
 RECT 23.58 1.435 23.72 1.99 ;
 RECT 25.305 1.8 25.445 1.99 ;
 RECT 21.35 1.39 21.49 2.22 ;
 RECT 22.735 1.37 22.875 2.22 ;
 RECT 23.58 2.13 23.72 2.22 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.03 0.59 20.4 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 OBS
 LAYER PO ;
 RECT 21.915 1.205 22.015 2 ;
 RECT 21.135 0.855 21.235 2.2 ;
 RECT 24 1.125 24.1 2.2 ;
 RECT 20.17 0.755 21.705 0.84 ;
 RECT 20.17 0.84 21.7 0.855 ;
 RECT 21.605 0.215 21.705 0.755 ;
 RECT 21.135 0.21 21.235 0.755 ;
 RECT 20.17 0.595 20.4 0.755 ;
 RECT 21.135 2.2 24.1 2.3 ;
 RECT 6.855 1.45 6.955 1.655 ;
 RECT 6.855 1.755 6.955 2.57 ;
 RECT 6.855 1.655 7.815 1.755 ;
 RECT 7.715 1.755 7.815 2.355 ;
 RECT 6.855 0.655 6.955 1.13 ;
 RECT 6.855 1.23 6.955 1.24 ;
 RECT 5.94 0.66 6.04 1.13 ;
 RECT 6.855 1.24 7.11 1.45 ;
 RECT 5.94 1.13 6.955 1.23 ;
 RECT 10.155 0.795 10.32 0.925 ;
 RECT 9.475 0.885 9.705 0.925 ;
 RECT 9.475 1.025 9.705 1.095 ;
 RECT 9.475 0.925 10.32 1.025 ;
 RECT 10.155 0.585 10.385 0.795 ;
 RECT 13.105 1.635 13.205 1.66 ;
 RECT 13.105 1.66 13.36 1.87 ;
 RECT 13.105 1.87 13.205 2.565 ;
 RECT 13.685 0.295 15.035 0.39 ;
 RECT 13.685 0.29 14.985 0.295 ;
 RECT 14.935 0.39 15.035 1.4 ;
 RECT 14.935 1.5 15.035 2.37 ;
 RECT 15.425 0.51 15.525 1.4 ;
 RECT 15.425 1.5 15.525 2.37 ;
 RECT 13.685 0.225 13.915 0.29 ;
 RECT 13.685 0.39 13.915 0.435 ;
 RECT 14.935 1.4 15.525 1.5 ;
 RECT 13.38 1.25 13.64 1.3 ;
 RECT 13.54 0.61 13.64 1.25 ;
 RECT 13.38 1.4 13.64 1.46 ;
 RECT 13.54 1.46 13.64 2.56 ;
 RECT 14.07 0.84 14.17 1.3 ;
 RECT 13.38 1.3 14.17 1.4 ;
 RECT 14.055 0.63 14.285 0.84 ;
 RECT 12.205 0.81 12.305 2.21 ;
 RECT 12.165 0.6 12.395 0.81 ;
 RECT 11.735 0.535 11.9 0.625 ;
 RECT 10.88 0.455 11.9 0.535 ;
 RECT 10.96 0.435 11.9 0.455 ;
 RECT 10.88 0.535 11.11 0.665 ;
 RECT 11.735 0.835 11.835 2.21 ;
 RECT 11.735 0.625 11.965 0.835 ;
 RECT 25.01 0.195 25.11 2.665 ;
 RECT 24 0.095 25.11 0.195 ;
 RECT 20.375 1.245 20.475 2.665 ;
 RECT 20.375 1.2 20.66 1.245 ;
 RECT 24 0.195 24.1 0.945 ;
 RECT 20.43 1.035 20.66 1.1 ;
 RECT 20.375 2.665 25.11 2.765 ;
 RECT 20.375 1.1 20.705 1.2 ;
 RECT 8.145 2.69 10.055 2.695 ;
 RECT 9.955 2.54 10.055 2.69 ;
 RECT 8.935 2.695 10.055 2.79 ;
 RECT 8.145 0.655 8.245 2.595 ;
 RECT 8.145 2.595 9.035 2.69 ;
 RECT 9.955 2.33 10.185 2.54 ;
 RECT 21.61 1.245 21.71 2.02 ;
 RECT 21.48 1.035 21.71 1.245 ;
 RECT 24.31 2.27 24.595 2.48 ;
 RECT 24.31 1.2 24.41 2.27 ;
 RECT 24.31 0.375 24.41 0.99 ;
 RECT 24.31 0.99 24.56 1.2 ;
 RECT 22.825 0.38 22.925 0.96 ;
 RECT 22.825 1.06 22.925 1.14 ;
 RECT 23.19 0.22 23.42 0.28 ;
 RECT 22.825 0.28 23.42 0.38 ;
 RECT 23.19 0.38 23.42 0.43 ;
 RECT 22.825 1.14 23.095 1.24 ;
 RECT 22.995 1.24 23.095 1.84 ;
 RECT 22.405 0.935 22.635 0.96 ;
 RECT 22.405 1.06 22.635 1.145 ;
 RECT 22.405 0.96 22.925 1.06 ;
 RECT 2.305 1.62 2.405 2.675 ;
 RECT 2.37 0.185 9.28 0.195 ;
 RECT 9.18 0.195 9.28 1.29 ;
 RECT 2.37 0.195 4.525 0.285 ;
 RECT 2.37 0.285 2.47 1.52 ;
 RECT 10.075 1.39 10.27 1.405 ;
 RECT 3.19 1.565 3.29 2.675 ;
 RECT 1.87 1.44 2.115 1.52 ;
 RECT 1.87 1.62 2.115 1.69 ;
 RECT 1.87 1.52 2.47 1.62 ;
 RECT 4.425 0.285 4.525 1.24 ;
 RECT 4.425 0.095 9.28 0.185 ;
 RECT 9.18 1.29 10.27 1.39 ;
 RECT 2.305 2.675 3.29 2.775 ;
 RECT 10.075 1.405 10.305 1.615 ;
 RECT 5.475 0.475 5.66 0.5 ;
 RECT 13.11 0.205 13.21 1.18 ;
 RECT 10.57 0.105 13.21 0.205 ;
 RECT 10.57 0.205 10.67 1.91 ;
 RECT 9.75 1.71 9.85 1.91 ;
 RECT 8.665 0.475 8.765 1.61 ;
 RECT 9.215 1.71 9.315 2.445 ;
 RECT 9.75 1.91 10.67 2.01 ;
 RECT 8.665 1.61 9.85 1.71 ;
 RECT 5.475 0.375 8.765 0.475 ;
 RECT 5.43 0.5 5.66 0.71 ;
 RECT 5.93 1.575 6.03 2.485 ;
 RECT 6.44 1.41 6.67 1.475 ;
 RECT 6.44 1.575 6.67 1.62 ;
 RECT 5.93 1.475 6.67 1.575 ;
 RECT 5.29 1.61 5.555 1.82 ;
 RECT 5.455 1.82 5.555 2.49 ;
 RECT 5.085 0.66 5.185 1.51 ;
 RECT 5.085 1.51 5.555 1.61 ;
 RECT 7.75 0.655 7.85 1.24 ;
 RECT 7.62 1.24 7.85 1.475 ;
 RECT 1.53 0.655 1.63 1.495 ;
 RECT 1.335 1.495 1.63 1.745 ;
 RECT 1.53 1.745 1.63 2.37 ;
 RECT 4.985 1.79 5.085 2.465 ;
 RECT 4.77 2.465 5.085 2.71 ;
 RECT 0.815 0.27 1.155 0.52 ;
 RECT 1.055 0.52 1.155 2.465 ;
 RECT 3.685 1.33 3.825 1.475 ;
 RECT 3.685 1.71 3.785 2.475 ;
 RECT 3.725 0.65 3.825 1.33 ;
 RECT 3.685 1.475 3.915 1.71 ;
 RECT 3.235 0.705 3.335 1.165 ;
 RECT 2.795 1.27 2.895 1.445 ;
 RECT 3.235 0.47 3.52 0.705 ;
 RECT 2.795 1.17 3.335 1.265 ;
 RECT 3.025 1.165 3.335 1.17 ;
 RECT 2.795 1.265 3.17 1.27 ;
 RECT 2.65 1.445 2.895 1.69 ;
 RECT 4.125 0.715 4.225 1.61 ;
 RECT 4.16 1.71 4.26 2.48 ;
 RECT 4.125 1.61 4.26 1.71 ;
 RECT 4.005 0.485 4.245 0.715 ;
 RECT 17.905 0.195 18.005 1.33 ;
 RECT 19.59 0.195 19.69 0.22 ;
 RECT 17.905 0.095 19.69 0.195 ;
 RECT 17.31 1.2 17.52 1.33 ;
 RECT 17.31 1.43 17.52 1.435 ;
 RECT 17.31 1.33 18.005 1.43 ;
 RECT 17.325 0.385 17.425 1.2 ;
 RECT 17.325 1.435 17.425 2.575 ;
 RECT 17.905 1.43 18.005 2.575 ;
 RECT 19.59 0.22 19.82 0.43 ;
 RECT 21.915 0.215 22.015 0.995 ;
 RECT 21.915 0.995 22.155 1.205 ;
 LAYER CO ;
 RECT 12.86 0.33 12.99 0.46 ;
 RECT 13.76 1.78 13.89 1.91 ;
 RECT 12.855 2.64 12.985 2.77 ;
 RECT 12.46 0.96 12.59 1.09 ;
 RECT 12.425 1.705 12.555 1.835 ;
 RECT 11.955 2.64 12.085 2.77 ;
 RECT 11.485 1.7 11.615 1.83 ;
 RECT 7.305 2.445 7.435 2.575 ;
 RECT 25.31 1.475 25.44 1.605 ;
 RECT 23.75 0.12 23.88 0.25 ;
 RECT 23.585 1.49 23.715 1.62 ;
 RECT 24.53 1.465 24.66 1.595 ;
 RECT 24.53 0.595 24.66 0.725 ;
 RECT 22.57 0.12 22.7 0.25 ;
 RECT 22.74 1.445 22.87 1.575 ;
 RECT 23.215 1.405 23.345 1.535 ;
 RECT 23.075 0.595 23.205 0.725 ;
 RECT 22.135 1.485 22.265 1.615 ;
 RECT 22.135 0.435 22.265 0.565 ;
 RECT 21.355 1.475 21.485 1.605 ;
 RECT 20.885 1.425 21.015 1.555 ;
 RECT 20.635 0.505 20.765 0.635 ;
 RECT 4.06 0.53 4.19 0.66 ;
 RECT 3.435 2.07 3.565 2.2 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 4.665 0.455 4.795 0.585 ;
 RECT 2.705 1.49 2.835 1.62 ;
 RECT 4.81 2.515 4.94 2.645 ;
 RECT 3.455 0.88 3.585 1.01 ;
 RECT 0.875 0.325 1.005 0.455 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 5.205 2.135 5.335 2.265 ;
 RECT 2.015 2.345 2.145 2.475 ;
 RECT 6.16 2.07 6.29 2.2 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.805 2.115 0.935 2.245 ;
 RECT 3.905 2.125 4.035 2.255 ;
 RECT 2.59 0.905 2.72 1.035 ;
 RECT 2.94 2.105 3.07 2.235 ;
 RECT 1.88 0.875 2.01 1.005 ;
 RECT 1.275 2.05 1.405 2.18 ;
 RECT 4.385 1.825 4.515 1.955 ;
 RECT 1.395 1.55 1.525 1.68 ;
 RECT 2.02 0.21 2.15 0.34 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 4.735 2.125 4.865 2.255 ;
 RECT 1.75 1.995 1.88 2.125 ;
 RECT 3.735 1.525 3.865 1.655 ;
 RECT 2.985 0.88 3.115 1.01 ;
 RECT 5.675 0.93 5.805 1.06 ;
 RECT 3.34 0.525 3.47 0.655 ;
 RECT 6.605 1.995 6.735 2.125 ;
 RECT 6.16 0.88 6.29 1.01 ;
 RECT 1.93 1.495 2.06 1.625 ;
 RECT 8.405 0.875 8.535 1.005 ;
 RECT 2.525 1.825 2.655 1.955 ;
 RECT 7.67 1.28 7.8 1.41 ;
 RECT 5.675 2.015 5.805 2.145 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 6.605 0.88 6.735 1.01 ;
 RECT 8.405 1.945 8.535 2.075 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 7.495 0.575 7.625 0.705 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 19.64 0.26 19.77 0.39 ;
 RECT 21.975 1.035 22.105 1.165 ;
 RECT 20.22 0.635 20.35 0.765 ;
 RECT 6.93 1.28 7.06 1.41 ;
 RECT 10.93 0.495 11.06 0.625 ;
 RECT 10.205 0.625 10.335 0.755 ;
 RECT 9.525 0.925 9.655 1.055 ;
 RECT 14.105 0.67 14.235 0.8 ;
 RECT 13.18 1.7 13.31 1.83 ;
 RECT 13.735 0.265 13.865 0.395 ;
 RECT 13.43 1.29 13.56 1.42 ;
 RECT 12.215 0.64 12.345 0.77 ;
 RECT 11.785 0.665 11.915 0.795 ;
 RECT 20.48 1.075 20.61 1.205 ;
 RECT 23.24 0.26 23.37 0.39 ;
 RECT 10.005 2.37 10.135 2.5 ;
 RECT 24.415 2.31 24.545 2.44 ;
 RECT 21.53 1.075 21.66 1.205 ;
 RECT 24.38 1.03 24.51 1.16 ;
 RECT 22.455 0.975 22.585 1.105 ;
 RECT 10.125 1.445 10.255 1.575 ;
 RECT 5.48 0.54 5.61 0.67 ;
 RECT 6.49 1.45 6.62 1.58 ;
 RECT 5.345 1.63 5.475 1.76 ;
 RECT 14.675 0.975 14.805 1.105 ;
 RECT 9.435 0.595 9.565 0.725 ;
 RECT 9.435 1.87 9.565 2 ;
 RECT 8.93 0.595 9.06 0.725 ;
 RECT 8.93 1.9 9.06 2.03 ;
 RECT 18.13 0.63 18.26 0.76 ;
 RECT 18.13 1.71 18.26 1.84 ;
 RECT 17.545 2.64 17.675 2.77 ;
 RECT 15.165 0.36 15.295 0.49 ;
 RECT 15.08 2.64 15.21 2.77 ;
 RECT 14.675 1.705 14.805 1.835 ;
 RECT 17.07 1.725 17.2 1.855 ;
 RECT 17.35 1.25 17.48 1.38 ;
 RECT 17.63 0.62 17.76 0.75 ;
 RECT 21.355 0.135 21.485 0.265 ;
 RECT 17.07 0.62 17.2 0.75 ;
 RECT 15.68 1.705 15.81 1.835 ;
 RECT 15.68 0.975 15.81 1.105 ;
 RECT 11.355 0.745 11.485 0.875 ;
 RECT 13.76 0.83 13.89 0.96 ;
 LAYER M1 ;
 RECT 1.875 0.825 2.015 1.475 ;
 RECT 1.68 1.99 1.93 2.13 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.11 ;
 RECT 0.58 2.25 0.72 2.255 ;
 RECT 0.58 0.87 1.005 1.01 ;
 RECT 0.58 2.11 1.005 2.25 ;
 RECT 1.55 0.67 1.69 1.195 ;
 RECT 0.58 1.195 1.69 1.335 ;
 RECT 2.98 0.36 3.12 2.035 ;
 RECT 1.55 0.53 2.435 0.67 ;
 RECT 2.295 0.22 3.12 0.36 ;
 RECT 2.295 0.36 2.435 0.53 ;
 RECT 2.935 2.035 3.12 2.17 ;
 RECT 2.935 2.17 3.075 2.305 ;
 RECT 2.585 1.67 2.725 1.82 ;
 RECT 2.585 1.96 2.725 2.51 ;
 RECT 2.585 0.5 2.725 1.44 ;
 RECT 2.585 1.44 2.84 1.67 ;
 RECT 2.455 1.82 2.725 1.96 ;
 RECT 2.585 2.51 5.06 2.65 ;
 RECT 3.275 1.22 3.59 1.36 ;
 RECT 3.45 0.805 3.59 1.22 ;
 RECT 3.36 1.96 3.64 2.215 ;
 RECT 3.275 1.36 3.415 1.82 ;
 RECT 3.275 1.82 4.855 1.96 ;
 RECT 4.715 1.79 4.855 1.82 ;
 RECT 5.29 1.58 5.53 1.65 ;
 RECT 5.29 1.79 5.53 1.835 ;
 RECT 4.715 1.65 5.53 1.79 ;
 RECT 19.59 0.36 19.82 0.43 ;
 RECT 20.985 0.36 21.125 0.565 ;
 RECT 19.59 0.22 21.125 0.36 ;
 RECT 21.725 0.705 21.865 0.75 ;
 RECT 20.985 0.565 21.865 0.705 ;
 RECT 21.725 0.75 21.99 0.89 ;
 RECT 21.85 0.89 21.99 0.995 ;
 RECT 21.85 0.995 22.155 1.205 ;
 RECT 10.155 0.585 11.11 0.63 ;
 RECT 10.88 0.63 11.11 0.665 ;
 RECT 10.88 0.455 11.11 0.49 ;
 RECT 10.18 0.49 11.11 0.585 ;
 RECT 10.155 0.63 10.385 0.795 ;
 RECT 9.43 0.525 9.57 0.885 ;
 RECT 9.43 0.885 9.705 1.095 ;
 RECT 9.43 1.095 9.57 2.065 ;
 RECT 14.055 0.63 14.285 0.635 ;
 RECT 14.055 0.775 14.285 0.84 ;
 RECT 16.665 0.36 16.805 0.635 ;
 RECT 14.05 0.635 16.805 0.775 ;
 RECT 17.345 0.36 17.485 1.46 ;
 RECT 16.665 0.22 17.485 0.36 ;
 RECT 11.48 1.51 11.62 1.695 ;
 RECT 11.41 1.695 11.69 1.835 ;
 RECT 12.455 1.095 12.595 1.37 ;
 RECT 12.42 1.51 12.56 1.7 ;
 RECT 11.48 1.37 13.61 1.51 ;
 RECT 13.38 1.25 13.61 1.37 ;
 RECT 12.385 0.955 12.665 1.095 ;
 RECT 12.355 1.7 12.63 1.84 ;
 RECT 11.735 0.36 11.965 0.835 ;
 RECT 12.535 0.36 12.675 0.665 ;
 RECT 11.735 0.22 12.68 0.36 ;
 RECT 13.755 0.22 13.895 0.225 ;
 RECT 13.755 0.435 13.895 0.665 ;
 RECT 12.535 0.665 13.895 0.805 ;
 RECT 13.755 0.805 13.895 1.98 ;
 RECT 13.685 0.225 13.915 0.435 ;
 RECT 23.19 0.29 23.56 0.43 ;
 RECT 23.42 0.43 23.56 0.71 ;
 RECT 23.19 0.22 23.42 0.29 ;
 RECT 24.84 0.85 24.98 1.385 ;
 RECT 24.525 1.525 24.665 1.73 ;
 RECT 23.42 0.71 24.98 0.85 ;
 RECT 24.525 0.51 24.665 0.71 ;
 RECT 24.525 1.385 24.98 1.525 ;
 RECT 9.955 2.42 10.185 2.54 ;
 RECT 9.955 2.28 20.165 2.42 ;
 RECT 20.025 2.42 20.165 2.52 ;
 RECT 24.365 2.48 24.505 2.52 ;
 RECT 20.025 2.52 24.505 2.66 ;
 RECT 24.365 2.27 24.595 2.48 ;
 RECT 20.43 1.035 20.88 1.055 ;
 RECT 20.43 1.225 20.66 1.245 ;
 RECT 20.43 1.195 21.02 1.225 ;
 RECT 20.705 0.64 20.845 1.015 ;
 RECT 20.57 1.015 20.88 1.035 ;
 RECT 20.88 1.225 21.02 1.75 ;
 RECT 20.585 0.5 20.845 0.64 ;
 RECT 20.43 1.055 21.71 1.195 ;
 RECT 21.48 1.035 21.71 1.055 ;
 RECT 21.48 1.195 21.71 1.245 ;
 RECT 23.21 1.18 23.35 1.605 ;
 RECT 23.07 0.73 23.21 1.04 ;
 RECT 23.005 0.59 23.28 0.73 ;
 RECT 24.33 0.99 24.56 1.04 ;
 RECT 24.33 1.18 24.56 1.2 ;
 RECT 23.07 1.04 24.56 1.18 ;
 RECT 22.45 0.73 22.59 0.935 ;
 RECT 22.13 0.355 22.27 0.59 ;
 RECT 22.45 1.145 22.59 1.345 ;
 RECT 22.13 1.485 22.27 1.76 ;
 RECT 22.13 0.59 22.59 0.73 ;
 RECT 22.13 1.345 22.59 1.485 ;
 RECT 22.405 0.935 22.635 1.145 ;
 RECT 10.09 2.05 10.23 2.055 ;
 RECT 10.09 1.915 11.265 1.985 ;
 RECT 10.09 1.91 11.26 1.915 ;
 RECT 10.09 1.615 10.23 1.91 ;
 RECT 13.13 1.87 13.315 1.985 ;
 RECT 10.09 1.985 13.315 2.05 ;
 RECT 11.12 2.05 13.315 2.125 ;
 RECT 13.13 1.66 13.36 1.87 ;
 RECT 10.075 1.405 10.305 1.615 ;
 RECT 3.27 0.52 3.87 0.66 ;
 RECT 3.73 0.66 3.87 1.015 ;
 RECT 5.275 0.505 5.66 0.71 ;
 RECT 5.43 0.5 5.66 0.505 ;
 RECT 3.73 1.015 5.415 1.155 ;
 RECT 5.275 0.71 5.415 1.015 ;
 RECT 6.6 1.62 6.74 1.735 ;
 RECT 6.6 1.875 6.74 2.18 ;
 RECT 6.6 0.81 6.74 1.41 ;
 RECT 6.44 1.41 6.74 1.62 ;
 RECT 6.6 1.735 7.795 1.875 ;
 RECT 7.655 1.415 7.795 1.735 ;
 RECT 7.61 1.275 7.87 1.415 ;
 RECT 3.835 2.12 4.935 2.26 ;
 RECT 4.395 1.44 4.535 1.52 ;
 RECT 3.665 1.52 4.535 1.66 ;
 RECT 5.67 0.865 5.81 1.3 ;
 RECT 4.395 1.3 5.81 1.44 ;
 RECT 5.67 1.44 5.81 2.215 ;
 RECT 6.155 0.82 6.295 2.33 ;
 RECT 6.155 2.47 6.295 2.475 ;
 RECT 7.005 2.165 7.145 2.33 ;
 RECT 7.005 2.47 7.145 2.475 ;
 RECT 6.155 2.33 7.145 2.47 ;
 RECT 7.005 2.025 9.065 2.16 ;
 RECT 7.005 2.16 9.06 2.165 ;
 RECT 8.925 0.525 9.065 2.025 ;
 RECT 8.4 0.765 8.54 2.025 ;
 RECT 1.79 1.63 1.93 1.99 ;
 RECT 1.79 1.475 2.135 1.63 ;
 END
END RDFFNSRARX1

MACRO RDFFNSRARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 26.88 BY 2.88 ;
 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.055 0.46 4.195 0.485 ;
 RECT 9.875 1.09 12.245 1.23 ;
 RECT 4.055 0.755 5.13 0.875 ;
 RECT 4.01 0.485 4.235 0.735 ;
 RECT 4.01 0.735 5.13 0.755 ;
 RECT 4.99 0.22 7.225 0.36 ;
 RECT 4.99 0.36 5.13 0.735 ;
 RECT 7.085 0.875 8.005 1.015 ;
 RECT 7.86 0.245 10.01 0.255 ;
 RECT 7.86 0.255 10.015 0.385 ;
 RECT 9.875 0.385 10.015 1.09 ;
 RECT 12.105 0.81 12.245 1.09 ;
 RECT 12.105 0.6 12.395 0.81 ;
 RECT 7.085 0.36 7.225 0.875 ;
 RECT 7.865 0.385 8.005 0.875 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 26.88 0.08 ;
 RECT 23.7 0.08 23.94 0.26 ;
 RECT 7.425 0.59 7.7 0.73 ;
 RECT 15.105 0.335 15.37 0.495 ;
 RECT 16.11 0.335 16.375 0.495 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 2.015 0.08 2.155 0.39 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.615 0.08 4.85 0.595 ;
 RECT 11.35 0.08 11.49 0.945 ;
 RECT 12.855 0.08 12.995 0.525 ;
 RECT 21.35 0.08 21.49 0.36 ;
 RECT 18.69 0.08 18.83 0.82 ;
 RECT 17.625 0.08 17.765 0.82 ;
 RECT 22.565 0.08 22.705 0.35 ;
 RECT 7.49 0.08 7.63 0.59 ;
 RECT 15.16 0.08 15.3 0.335 ;
 RECT 16.165 0.08 16.305 0.335 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 26.88 2.96 ;
 RECT 1.945 2.34 2.195 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.27 1.98 1.41 2.8 ;
 RECT 5.2 2.07 5.34 2.8 ;
 RECT 7.3 2.375 7.44 2.8 ;
 RECT 11.95 2.57 12.09 2.8 ;
 RECT 15.075 2.57 15.215 2.8 ;
 RECT 12.85 2.57 12.99 2.8 ;
 RECT 16.08 2.57 16.22 2.8 ;
 RECT 18.605 2.57 18.745 2.8 ;
 RECT 17.54 2.57 17.68 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.475 1.65 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.765 0.22 1.13 0.615 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.465 1.205 14.82 1.445 ;
 RECT 14.67 0.915 14.81 1.205 ;
 RECT 14.67 1.84 14.81 1.885 ;
 RECT 14.67 1.445 14.81 1.7 ;
 RECT 15.675 1.84 15.815 1.885 ;
 RECT 15.675 0.915 15.815 1.7 ;
 RECT 16.65 1.84 16.79 1.885 ;
 RECT 16.65 0.915 16.79 1.7 ;
 RECT 14.67 1.7 16.79 1.84 ;
 END
 ANTENNADIFFAREA 1.145 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 16.945 1.095 17.205 1.335 ;
 RECT 17.065 0.51 17.205 1.095 ;
 RECT 18.125 1.905 18.265 1.91 ;
 RECT 18.125 0.56 18.265 1.765 ;
 RECT 19.19 1.905 19.33 1.91 ;
 RECT 19.19 0.56 19.33 1.765 ;
 RECT 17.065 1.905 17.205 1.915 ;
 RECT 17.065 1.335 17.205 1.765 ;
 RECT 17.065 1.765 19.33 1.905 ;
 END
 ANTENNADIFFAREA 1.043 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.88 1.155 7.165 1.49 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 25.26 1.435 25.6 1.8 ;
 RECT 23.58 1.99 25.445 2.13 ;
 RECT 21.35 2.22 23.72 2.36 ;
 RECT 23.58 1.435 23.72 1.99 ;
 RECT 25.305 1.8 25.445 1.99 ;
 RECT 21.35 1.39 21.49 2.22 ;
 RECT 22.735 1.37 22.875 2.22 ;
 RECT 23.58 2.13 23.72 2.22 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.03 0.59 20.4 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 OBS
 LAYER PO ;
 RECT 6.855 1.755 6.955 2.57 ;
 RECT 6.855 1.655 7.815 1.755 ;
 RECT 7.715 1.755 7.815 2.355 ;
 RECT 6.855 0.655 6.955 1.13 ;
 RECT 6.855 1.23 6.955 1.24 ;
 RECT 5.94 0.66 6.04 1.13 ;
 RECT 6.855 1.24 7.11 1.45 ;
 RECT 5.94 1.13 6.955 1.23 ;
 RECT 10.155 0.795 10.32 0.925 ;
 RECT 9.475 0.885 9.705 0.925 ;
 RECT 9.475 1.025 9.705 1.095 ;
 RECT 9.475 0.925 10.32 1.025 ;
 RECT 10.155 0.585 10.385 0.795 ;
 RECT 13.105 1.76 13.36 1.97 ;
 RECT 13.105 1.97 13.205 2.565 ;
 RECT 14.935 0.39 15.035 1.4 ;
 RECT 14.935 1.5 15.035 2.37 ;
 RECT 13.685 0.29 15.035 0.39 ;
 RECT 15.94 0.515 16.04 1.4 ;
 RECT 15.94 1.5 16.04 2.37 ;
 RECT 16.43 0.51 16.53 1.4 ;
 RECT 16.43 1.5 16.53 2.37 ;
 RECT 14.935 1.4 16.53 1.5 ;
 RECT 15.425 0.51 15.525 1.4 ;
 RECT 15.425 1.5 15.525 2.37 ;
 RECT 13.685 0.225 13.915 0.29 ;
 RECT 13.685 0.39 13.915 0.435 ;
 RECT 13.375 1.365 13.64 1.415 ;
 RECT 13.375 1.515 13.64 1.565 ;
 RECT 14.07 0.84 14.17 1.415 ;
 RECT 13.54 0.61 13.64 1.36 ;
 RECT 13.38 1.36 13.64 1.365 ;
 RECT 13.54 1.57 13.64 2.56 ;
 RECT 13.38 1.565 13.64 1.57 ;
 RECT 13.375 1.415 14.17 1.515 ;
 RECT 14.055 0.63 14.285 0.84 ;
 RECT 12.205 0.81 12.305 2.21 ;
 RECT 12.165 0.6 12.395 0.81 ;
 RECT 11.735 0.535 11.9 0.625 ;
 RECT 10.88 0.455 11.9 0.535 ;
 RECT 10.96 0.435 11.9 0.455 ;
 RECT 10.88 0.535 11.11 0.665 ;
 RECT 11.735 0.835 11.835 2.21 ;
 RECT 11.735 0.625 11.965 0.835 ;
 RECT 20.375 1.1 20.66 1.245 ;
 RECT 25.01 0.195 25.11 2.665 ;
 RECT 24 0.095 25.11 0.195 ;
 RECT 20.375 1.245 20.475 2.665 ;
 RECT 24 0.195 24.1 0.945 ;
 RECT 20.43 1.035 20.66 1.1 ;
 RECT 20.375 2.665 25.11 2.765 ;
 RECT 8.145 2.69 10.055 2.695 ;
 RECT 9.955 2.54 10.055 2.69 ;
 RECT 8.935 2.695 10.055 2.79 ;
 RECT 8.145 0.655 8.245 2.595 ;
 RECT 8.145 2.595 9.035 2.69 ;
 RECT 9.955 2.33 10.185 2.54 ;
 RECT 21.61 1.245 21.71 2.02 ;
 RECT 21.48 1.035 21.71 1.245 ;
 RECT 24.31 2.27 24.595 2.48 ;
 RECT 24.31 1.2 24.41 2.27 ;
 RECT 24.31 0.375 24.41 0.99 ;
 RECT 24.31 0.99 24.56 1.2 ;
 RECT 22.825 0.38 22.925 0.96 ;
 RECT 22.825 1.06 22.925 1.14 ;
 RECT 23.19 0.22 23.42 0.28 ;
 RECT 22.825 0.28 23.42 0.38 ;
 RECT 23.19 0.38 23.42 0.43 ;
 RECT 22.825 1.14 23.095 1.24 ;
 RECT 22.995 1.24 23.095 1.84 ;
 RECT 22.405 0.935 22.635 0.96 ;
 RECT 22.405 1.06 22.635 1.145 ;
 RECT 22.405 0.96 22.925 1.06 ;
 RECT 2.305 1.62 2.405 2.675 ;
 RECT 2.37 0.185 9.28 0.195 ;
 RECT 9.18 0.195 9.28 1.29 ;
 RECT 2.37 0.195 4.525 0.285 ;
 RECT 2.37 0.285 2.47 1.52 ;
 RECT 10.075 1.39 10.27 1.405 ;
 RECT 3.19 1.565 3.29 2.675 ;
 RECT 1.87 1.44 2.115 1.52 ;
 RECT 1.87 1.62 2.115 1.69 ;
 RECT 1.87 1.52 2.47 1.62 ;
 RECT 4.425 0.285 4.525 1.24 ;
 RECT 4.425 0.095 9.28 0.185 ;
 RECT 9.18 1.29 10.27 1.39 ;
 RECT 2.305 2.675 3.29 2.775 ;
 RECT 10.075 1.405 10.305 1.615 ;
 RECT 5.475 0.475 5.66 0.5 ;
 RECT 13.11 0.205 13.21 1.18 ;
 RECT 10.57 0.105 13.21 0.205 ;
 RECT 10.57 0.205 10.67 1.91 ;
 RECT 9.75 1.71 9.85 1.91 ;
 RECT 8.665 0.475 8.765 1.61 ;
 RECT 8.665 1.61 9.85 1.71 ;
 RECT 8.665 1.71 8.765 1.725 ;
 RECT 9.215 1.71 9.315 2.445 ;
 RECT 9.75 1.91 10.67 2.01 ;
 RECT 5.475 0.375 8.765 0.475 ;
 RECT 5.43 0.5 5.66 0.71 ;
 RECT 5.93 1.575 6.03 2.485 ;
 RECT 6.44 1.41 6.67 1.475 ;
 RECT 6.44 1.575 6.67 1.62 ;
 RECT 5.93 1.475 6.67 1.575 ;
 RECT 7.75 0.655 7.85 1.24 ;
 RECT 7.62 1.24 7.85 1.475 ;
 RECT 1.53 0.655 1.63 1.495 ;
 RECT 1.335 1.495 1.63 1.745 ;
 RECT 1.53 1.745 1.63 2.37 ;
 RECT 0.815 0.27 1.155 0.52 ;
 RECT 1.055 0.52 1.155 2.465 ;
 RECT 3.685 1.33 3.825 1.475 ;
 RECT 3.685 1.71 3.785 2.475 ;
 RECT 3.725 0.65 3.825 1.33 ;
 RECT 3.685 1.475 3.915 1.71 ;
 RECT 4.77 2.465 5.085 2.71 ;
 RECT 4.985 1.79 5.085 2.465 ;
 RECT 4.125 0.715 4.225 1.61 ;
 RECT 4.16 1.71 4.26 2.48 ;
 RECT 4.125 1.61 4.26 1.71 ;
 RECT 4.005 0.485 4.245 0.715 ;
 RECT 5.29 1.61 5.555 1.82 ;
 RECT 5.455 1.82 5.555 2.49 ;
 RECT 5.085 0.66 5.185 1.51 ;
 RECT 5.085 1.51 5.555 1.61 ;
 RECT 3.235 0.705 3.335 1.165 ;
 RECT 2.795 1.27 2.895 1.445 ;
 RECT 3.235 0.47 3.52 0.705 ;
 RECT 2.795 1.17 3.335 1.265 ;
 RECT 2.795 1.265 3.17 1.27 ;
 RECT 3.025 1.165 3.335 1.17 ;
 RECT 2.65 1.445 2.895 1.69 ;
 RECT 17.905 0.385 18.005 1.33 ;
 RECT 17.905 1.43 18.005 2.575 ;
 RECT 17.325 1.22 17.59 1.33 ;
 RECT 17.325 0.385 17.425 1.22 ;
 RECT 18.97 0.365 19.07 1.33 ;
 RECT 17.325 1.33 19.07 1.43 ;
 RECT 18.39 0.385 18.49 1.33 ;
 RECT 18.39 1.43 18.49 2.575 ;
 RECT 18.97 1.43 19.07 2.575 ;
 RECT 19.59 0.22 19.82 0.265 ;
 RECT 19.59 0.365 19.82 0.43 ;
 RECT 17.325 1.43 17.425 2.575 ;
 RECT 18.97 0.265 19.82 0.365 ;
 RECT 21.915 0.215 22.015 0.995 ;
 RECT 21.915 0.995 22.155 1.205 ;
 RECT 21.915 1.205 22.015 2 ;
 RECT 21.135 0.855 21.235 2.2 ;
 RECT 24 1.125 24.1 2.2 ;
 RECT 20.17 0.755 21.705 0.84 ;
 RECT 20.17 0.84 21.7 0.855 ;
 RECT 21.605 0.215 21.705 0.755 ;
 RECT 21.135 0.21 21.235 0.755 ;
 RECT 20.17 0.595 20.4 0.755 ;
 RECT 21.135 2.2 24.1 2.3 ;
 RECT 6.855 1.45 6.955 1.655 ;
 LAYER CO ;
 RECT 6.16 2.07 6.29 2.2 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.805 2.115 0.935 2.245 ;
 RECT 3.905 2.125 4.035 2.255 ;
 RECT 2.59 0.905 2.72 1.035 ;
 RECT 2.94 2.105 3.07 2.235 ;
 RECT 1.88 0.875 2.01 1.005 ;
 RECT 1.275 2.05 1.405 2.18 ;
 RECT 4.385 1.825 4.515 1.955 ;
 RECT 1.395 1.55 1.525 1.68 ;
 RECT 2.02 0.21 2.15 0.34 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 4.735 2.125 4.865 2.255 ;
 RECT 1.75 1.995 1.88 2.125 ;
 RECT 3.735 1.525 3.865 1.655 ;
 RECT 2.985 0.88 3.115 1.01 ;
 RECT 5.675 0.93 5.805 1.06 ;
 RECT 3.34 0.525 3.47 0.655 ;
 RECT 6.605 1.995 6.735 2.125 ;
 RECT 6.16 0.88 6.29 1.01 ;
 RECT 1.93 1.495 2.06 1.625 ;
 RECT 8.405 0.875 8.535 1.005 ;
 RECT 5.345 1.63 5.475 1.76 ;
 RECT 14.675 0.975 14.805 1.105 ;
 RECT 9.435 0.595 9.565 0.725 ;
 RECT 9.435 1.87 9.565 2 ;
 RECT 8.93 0.595 9.06 0.725 ;
 RECT 8.93 1.9 9.06 2.03 ;
 RECT 18.13 0.63 18.26 0.76 ;
 RECT 18.13 1.71 18.26 1.84 ;
 RECT 17.545 2.64 17.675 2.77 ;
 RECT 2.525 1.825 2.655 1.955 ;
 RECT 7.67 1.28 7.8 1.41 ;
 RECT 5.675 2.015 5.805 2.145 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 6.605 0.88 6.735 1.01 ;
 RECT 8.405 1.945 8.535 2.075 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 7.495 0.595 7.625 0.725 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 4.06 0.53 4.19 0.66 ;
 RECT 3.435 2.07 3.565 2.2 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 4.665 0.455 4.795 0.585 ;
 RECT 2.705 1.49 2.835 1.62 ;
 RECT 4.81 2.515 4.94 2.645 ;
 RECT 3.455 0.88 3.585 1.01 ;
 RECT 0.875 0.325 1.005 0.455 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 5.205 2.135 5.335 2.265 ;
 RECT 17.41 1.26 17.54 1.39 ;
 RECT 19.64 0.26 19.77 0.39 ;
 RECT 21.975 1.035 22.105 1.165 ;
 RECT 20.22 0.635 20.35 0.765 ;
 RECT 6.93 1.28 7.06 1.41 ;
 RECT 10.93 0.495 11.06 0.625 ;
 RECT 10.205 0.625 10.335 0.755 ;
 RECT 9.525 0.925 9.655 1.055 ;
 RECT 14.105 0.67 14.235 0.8 ;
 RECT 13.18 1.8 13.31 1.93 ;
 RECT 13.735 0.265 13.865 0.395 ;
 RECT 13.43 1.4 13.56 1.53 ;
 RECT 12.215 0.64 12.345 0.77 ;
 RECT 11.785 0.665 11.915 0.795 ;
 RECT 20.48 1.075 20.61 1.205 ;
 RECT 23.24 0.26 23.37 0.39 ;
 RECT 10.005 2.37 10.135 2.5 ;
 RECT 24.415 2.31 24.545 2.44 ;
 RECT 21.53 1.075 21.66 1.205 ;
 RECT 24.38 1.03 24.51 1.16 ;
 RECT 22.455 0.975 22.585 1.105 ;
 RECT 10.125 1.445 10.255 1.575 ;
 RECT 5.48 0.54 5.61 0.67 ;
 RECT 6.49 1.45 6.62 1.58 ;
 RECT 15.165 0.36 15.295 0.49 ;
 RECT 15.08 2.64 15.21 2.77 ;
 RECT 14.675 1.705 14.805 1.835 ;
 RECT 17.07 1.725 17.2 1.855 ;
 RECT 17.63 0.62 17.76 0.75 ;
 RECT 21.355 0.135 21.485 0.265 ;
 RECT 19.195 1.71 19.325 1.84 ;
 RECT 18.61 2.64 18.74 2.77 ;
 RECT 18.695 0.62 18.825 0.75 ;
 RECT 19.195 0.63 19.325 0.76 ;
 RECT 16.655 1.705 16.785 1.835 ;
 RECT 16.655 0.975 16.785 1.105 ;
 RECT 16.17 0.36 16.3 0.49 ;
 RECT 16.085 2.64 16.215 2.77 ;
 RECT 17.07 0.62 17.2 0.75 ;
 RECT 15.68 1.705 15.81 1.835 ;
 RECT 15.68 0.975 15.81 1.105 ;
 RECT 11.355 0.745 11.485 0.875 ;
 RECT 13.76 0.83 13.89 0.96 ;
 RECT 12.86 0.33 12.99 0.46 ;
 RECT 13.76 1.78 13.89 1.91 ;
 RECT 12.855 2.64 12.985 2.77 ;
 RECT 12.46 0.96 12.59 1.09 ;
 RECT 12.425 1.705 12.555 1.835 ;
 RECT 11.955 2.64 12.085 2.77 ;
 RECT 11.485 1.7 11.615 1.83 ;
 RECT 7.305 2.445 7.435 2.575 ;
 RECT 25.31 1.475 25.44 1.605 ;
 RECT 23.75 0.12 23.88 0.25 ;
 RECT 23.585 1.49 23.715 1.62 ;
 RECT 24.53 1.465 24.66 1.595 ;
 RECT 24.53 0.595 24.66 0.725 ;
 RECT 22.57 0.12 22.7 0.25 ;
 RECT 22.74 1.445 22.87 1.575 ;
 RECT 23.215 1.405 23.345 1.535 ;
 RECT 23.075 0.595 23.205 0.725 ;
 RECT 22.135 1.485 22.265 1.615 ;
 RECT 22.135 0.435 22.265 0.565 ;
 RECT 21.355 1.475 21.485 1.605 ;
 RECT 20.885 1.425 21.015 1.555 ;
 RECT 20.635 0.505 20.765 0.635 ;
 RECT 2.015 2.345 2.145 2.475 ;
 LAYER M1 ;
 RECT 5.67 1.44 5.81 2.215 ;
 RECT 3.275 1.22 3.59 1.36 ;
 RECT 3.45 0.805 3.59 1.22 ;
 RECT 3.36 1.96 3.64 2.215 ;
 RECT 3.275 1.36 3.415 1.82 ;
 RECT 3.275 1.82 4.855 1.96 ;
 RECT 4.715 1.79 4.855 1.82 ;
 RECT 5.29 1.58 5.53 1.65 ;
 RECT 5.29 1.79 5.53 1.835 ;
 RECT 4.715 1.65 5.53 1.79 ;
 RECT 6.6 1.62 6.74 1.735 ;
 RECT 6.6 1.875 6.74 2.18 ;
 RECT 6.6 0.81 6.74 1.41 ;
 RECT 6.44 1.41 6.74 1.62 ;
 RECT 7.665 1.415 7.805 1.735 ;
 RECT 6.6 1.735 7.805 1.875 ;
 RECT 7.605 1.275 7.87 1.415 ;
 RECT 1.79 1.63 1.93 1.99 ;
 RECT 1.79 1.475 2.135 1.63 ;
 RECT 1.875 0.825 2.015 1.475 ;
 RECT 1.68 1.99 1.93 2.13 ;
 RECT 23.07 0.73 23.21 1.04 ;
 RECT 23.21 1.18 23.35 1.605 ;
 RECT 23.005 0.59 23.28 0.73 ;
 RECT 24.33 0.99 24.56 1.04 ;
 RECT 23.07 1.04 24.56 1.18 ;
 RECT 24.33 1.18 24.56 1.2 ;
 RECT 23.19 0.29 23.56 0.43 ;
 RECT 23.42 0.43 23.56 0.71 ;
 RECT 23.19 0.22 23.42 0.29 ;
 RECT 24.84 0.85 24.98 1.385 ;
 RECT 24.525 1.525 24.665 1.73 ;
 RECT 23.42 0.71 24.98 0.85 ;
 RECT 24.525 0.51 24.665 0.71 ;
 RECT 24.525 1.385 24.98 1.525 ;
 RECT 22.45 1.145 22.59 1.345 ;
 RECT 22.13 1.485 22.27 1.76 ;
 RECT 22.45 0.73 22.59 0.935 ;
 RECT 22.13 0.355 22.27 0.59 ;
 RECT 22.13 1.345 22.59 1.485 ;
 RECT 22.405 0.935 22.635 1.145 ;
 RECT 22.13 0.59 22.59 0.73 ;
 RECT 20.43 1.225 20.66 1.245 ;
 RECT 20.43 1.195 21.02 1.225 ;
 RECT 20.57 1.015 20.88 1.035 ;
 RECT 20.43 1.035 20.88 1.055 ;
 RECT 20.705 0.64 20.845 1.015 ;
 RECT 20.88 1.225 21.02 1.75 ;
 RECT 20.585 0.5 20.845 0.64 ;
 RECT 21.48 1.035 21.71 1.055 ;
 RECT 21.48 1.195 21.71 1.245 ;
 RECT 20.43 1.055 21.71 1.195 ;
 RECT 19.59 0.36 19.82 0.43 ;
 RECT 20.985 0.36 21.125 0.565 ;
 RECT 19.59 0.22 21.125 0.36 ;
 RECT 21.725 0.705 21.865 0.75 ;
 RECT 21.85 0.995 22.155 1.205 ;
 RECT 21.85 0.89 21.99 0.995 ;
 RECT 21.725 0.75 21.99 0.89 ;
 RECT 20.985 0.565 21.865 0.705 ;
 RECT 14.055 0.63 14.285 0.635 ;
 RECT 14.055 0.775 14.285 0.84 ;
 RECT 14.05 0.635 16.805 0.775 ;
 RECT 16.665 0.36 16.805 0.635 ;
 RECT 17.345 0.36 17.485 1.22 ;
 RECT 17.345 1.22 17.59 1.43 ;
 RECT 17.345 1.43 17.485 1.435 ;
 RECT 16.665 0.22 17.485 0.36 ;
 RECT 9.43 0.525 9.57 0.885 ;
 RECT 9.43 1.095 9.57 2.065 ;
 RECT 9.43 0.885 9.705 1.095 ;
 RECT 6.155 0.82 6.295 2.33 ;
 RECT 6.155 2.47 6.295 2.475 ;
 RECT 7.005 2.165 7.145 2.33 ;
 RECT 7.005 2.47 7.145 2.475 ;
 RECT 6.155 2.33 7.145 2.47 ;
 RECT 8.085 2.165 8.225 2.295 ;
 RECT 8.4 0.765 8.54 2.295 ;
 RECT 8.4 2.435 8.54 2.44 ;
 RECT 8.925 0.525 9.065 2.295 ;
 RECT 8.925 2.435 9.065 2.44 ;
 RECT 7.005 2.025 8.225 2.165 ;
 RECT 8.085 2.295 9.065 2.435 ;
 RECT 11.735 0.36 11.965 0.835 ;
 RECT 12.535 0.36 12.675 0.665 ;
 RECT 11.735 0.22 12.68 0.36 ;
 RECT 13.755 0.22 13.895 0.225 ;
 RECT 13.755 0.435 13.895 0.665 ;
 RECT 12.535 0.665 13.895 0.805 ;
 RECT 13.755 0.805 13.895 1.98 ;
 RECT 13.685 0.225 13.915 0.435 ;
 RECT 10.155 0.585 11.11 0.63 ;
 RECT 10.88 0.63 11.11 0.665 ;
 RECT 10.88 0.455 11.11 0.49 ;
 RECT 10.18 0.49 11.11 0.585 ;
 RECT 10.155 0.63 10.385 0.795 ;
 RECT 3.27 0.52 3.87 0.66 ;
 RECT 3.73 0.66 3.87 1.015 ;
 RECT 5.275 0.505 5.66 0.71 ;
 RECT 3.73 1.015 5.415 1.155 ;
 RECT 5.275 0.71 5.415 1.015 ;
 RECT 5.43 0.5 5.66 0.505 ;
 RECT 2.585 1.67 2.725 1.82 ;
 RECT 2.585 1.96 2.725 2.51 ;
 RECT 2.585 0.5 2.725 1.44 ;
 RECT 2.585 1.44 2.84 1.67 ;
 RECT 2.455 1.82 2.725 1.96 ;
 RECT 2.585 2.51 5.06 2.65 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.11 ;
 RECT 0.58 2.25 0.72 2.255 ;
 RECT 0.58 0.87 1.005 1.01 ;
 RECT 0.58 2.11 1.005 2.25 ;
 RECT 0.58 1.195 1.69 1.335 ;
 RECT 1.55 0.67 1.69 1.195 ;
 RECT 2.98 0.36 3.12 2.035 ;
 RECT 2.295 0.22 3.12 0.36 ;
 RECT 1.55 0.53 2.435 0.67 ;
 RECT 2.935 2.17 3.075 2.305 ;
 RECT 2.935 2.035 3.12 2.17 ;
 RECT 2.295 0.36 2.435 0.53 ;
 RECT 9.955 2.42 10.185 2.54 ;
 RECT 20.025 2.42 20.165 2.52 ;
 RECT 9.955 2.28 20.165 2.42 ;
 RECT 24.365 2.48 24.505 2.52 ;
 RECT 20.025 2.52 24.505 2.66 ;
 RECT 24.365 2.27 24.595 2.48 ;
 RECT 11.48 1.51 11.62 1.695 ;
 RECT 11.41 1.695 11.69 1.835 ;
 RECT 12.455 1.095 12.595 1.37 ;
 RECT 12.42 1.51 12.56 1.7 ;
 RECT 13.38 1.36 13.61 1.37 ;
 RECT 13.38 1.51 13.61 1.57 ;
 RECT 11.48 1.37 13.61 1.51 ;
 RECT 12.385 0.955 12.665 1.095 ;
 RECT 12.355 1.7 12.63 1.84 ;
 RECT 10.09 2.05 10.23 2.055 ;
 RECT 10.09 1.915 11.265 1.985 ;
 RECT 10.09 1.91 11.26 1.915 ;
 RECT 10.09 1.615 10.23 1.91 ;
 RECT 13.13 1.97 13.315 1.985 ;
 RECT 10.09 1.985 13.315 2.05 ;
 RECT 11.12 2.05 13.315 2.125 ;
 RECT 13.13 1.76 13.36 1.97 ;
 RECT 10.075 1.405 10.305 1.615 ;
 RECT 3.835 2.12 4.935 2.26 ;
 RECT 4.395 1.44 4.535 1.52 ;
 RECT 3.665 1.52 4.535 1.66 ;
 RECT 5.67 0.865 5.81 1.3 ;
 RECT 4.395 1.3 5.81 1.44 ;
 END
END RDFFNSRARX2

MACRO RDFFNSRASRNX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.84 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.895 0.59 21.265 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.125 1.435 26.465 1.8 ;
 RECT 24.445 1.99 26.31 2.13 ;
 RECT 22.215 2.22 24.585 2.36 ;
 RECT 26.17 1.8 26.31 1.99 ;
 RECT 24.445 1.435 24.585 1.99 ;
 RECT 22.215 1.39 22.355 2.22 ;
 RECT 23.6 1.37 23.74 2.22 ;
 RECT 24.445 2.13 24.585 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.8 0.22 1.165 0.525 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.825 0.08 2.105 0.295 ;
 RECT 24.565 0.08 24.805 0.26 ;
 RECT 5.755 0.31 6.045 0.45 ;
 RECT 13.365 0.275 14.39 0.415 ;
 RECT 14.25 0.75 15.195 0.89 ;
 RECT 0 -0.08 27.84 0.08 ;
 RECT 0.335 0.08 0.475 0.775 ;
 RECT 1.305 0.08 1.445 0.97 ;
 RECT 4.65 0.08 4.885 0.46 ;
 RECT 9.505 0.08 9.645 0.815 ;
 RECT 19.37 0.08 19.51 0.82 ;
 RECT 22.215 0.08 22.355 0.36 ;
 RECT 23.43 0.08 23.57 0.35 ;
 RECT 5.835 0.08 5.975 0.31 ;
 RECT 13.365 0.415 13.505 0.945 ;
 RECT 13.365 0.08 13.505 0.275 ;
 RECT 15.055 0.89 15.195 1.11 ;
 RECT 14.25 0.415 14.39 0.75 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 19.225 2.6 19.49 2.8 ;
 RECT 9.25 2.215 9.525 2.355 ;
 RECT 0 2.8 27.84 2.96 ;
 RECT 0.335 1.74 0.475 2.8 ;
 RECT 1.98 2.34 2.23 2.8 ;
 RECT 1.305 1.98 1.445 2.8 ;
 RECT 5.835 1.98 5.975 2.8 ;
 RECT 6.865 2 7.005 2.8 ;
 RECT 5.355 2.07 5.495 2.8 ;
 RECT 12.275 2.335 12.545 2.8 ;
 RECT 9.315 2.355 9.455 2.8 ;
 RECT 9.315 2.195 9.455 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.355 1.475 1.685 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.74 1.095 20.15 1.335 ;
 RECT 19.87 0.56 20.01 1.095 ;
 RECT 18.81 1.905 18.95 1.915 ;
 RECT 18.81 0.78 18.95 1.765 ;
 RECT 19.87 1.905 20.01 1.91 ;
 RECT 18.795 1.765 20.01 1.905 ;
 RECT 19.87 1.335 20.01 1.765 ;
 END
 ANTENNADIFFAREA 0.723 ;
 END QN

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.72 2.12 10.04 2.485 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.045 0.485 4.36 0.605 ;
 RECT 9.88 1.095 10.02 1.1 ;
 RECT 8.965 0.955 10.02 1.095 ;
 RECT 9.88 0.22 10.02 0.245 ;
 RECT 9.875 0.245 12.025 0.255 ;
 RECT 9.875 0.255 12.03 0.385 ;
 RECT 11.89 1.09 13.88 1.23 ;
 RECT 14.085 1.56 14.315 1.6 ;
 RECT 13.74 1.42 14.315 1.56 ;
 RECT 14.085 1.39 14.315 1.42 ;
 RECT 4.045 0.605 9.105 0.745 ;
 RECT 8.965 0.745 9.105 0.955 ;
 RECT 9.88 0.385 10.02 0.955 ;
 RECT 11.89 0.385 12.03 1.09 ;
 RECT 13.74 1.23 13.88 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.21 2.12 7.495 2.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 OBS
 LAYER PO ;
 RECT 6.09 1.825 6.19 2.51 ;
 RECT 17.655 0.195 17.755 2.055 ;
 RECT 16.19 0.77 16.29 2.055 ;
 RECT 17.655 0.095 20.49 0.195 ;
 RECT 16.19 0.55 16.29 0.56 ;
 RECT 16.19 0.56 16.445 0.77 ;
 RECT 16.19 2.055 17.755 2.155 ;
 RECT 20.255 0.195 20.49 0.43 ;
 RECT 14.22 0.73 14.32 1.39 ;
 RECT 14.085 1.39 14.32 1.6 ;
 RECT 14.22 1.6 14.32 2.39 ;
 RECT 2.405 0.285 2.505 1.52 ;
 RECT 1.905 1.52 2.505 1.62 ;
 RECT 2.405 0.185 11.295 0.195 ;
 RECT 4.46 0.095 11.295 0.185 ;
 RECT 2.405 0.195 4.56 0.285 ;
 RECT 11.195 0.195 11.295 1.29 ;
 RECT 12.09 1.39 12.285 1.405 ;
 RECT 3.225 1.565 3.325 2.675 ;
 RECT 2.34 1.62 2.44 2.675 ;
 RECT 1.905 1.44 2.15 1.52 ;
 RECT 1.905 1.62 2.15 1.69 ;
 RECT 4.46 0.285 4.56 1.24 ;
 RECT 11.195 1.29 12.285 1.39 ;
 RECT 2.34 2.675 3.325 2.775 ;
 RECT 12.09 1.405 12.32 1.615 ;
 RECT 22.475 1.245 22.575 2.02 ;
 RECT 22.345 1.035 22.575 1.245 ;
 RECT 12.585 0.105 15.41 0.205 ;
 RECT 12.585 0.205 12.685 1.91 ;
 RECT 15.31 0.205 15.41 1.265 ;
 RECT 11.765 1.71 11.865 1.91 ;
 RECT 10.68 1.61 11.865 1.71 ;
 RECT 10.68 0.475 10.78 1.61 ;
 RECT 11.23 1.71 11.33 2.425 ;
 RECT 7.345 0.475 7.445 0.895 ;
 RECT 11.765 1.91 12.685 2.01 ;
 RECT 7.345 0.375 10.78 0.475 ;
 RECT 7.22 0.895 7.45 1.105 ;
 RECT 12.895 0.455 14.825 0.535 ;
 RECT 14.595 0.535 14.825 0.6 ;
 RECT 14.595 0.39 14.825 0.435 ;
 RECT 12.975 0.435 14.825 0.455 ;
 RECT 12.895 0.535 13.125 0.665 ;
 RECT 13.75 0.535 13.98 0.835 ;
 RECT 13.75 0.835 13.85 2.39 ;
 RECT 22.78 0.215 22.88 0.995 ;
 RECT 22.78 0.995 23.02 1.205 ;
 RECT 22.78 1.205 22.88 2 ;
 RECT 25.175 0.375 25.275 0.99 ;
 RECT 25.175 0.99 25.425 1.2 ;
 RECT 25.175 1.2 25.275 2.27 ;
 RECT 25.175 2.27 25.46 2.48 ;
 RECT 10.16 0.655 10.26 2.305 ;
 RECT 10.465 2.3 10.695 2.305 ;
 RECT 10.465 2.405 10.695 2.51 ;
 RECT 10.16 2.305 10.695 2.405 ;
 RECT 22 0.21 22.1 0.755 ;
 RECT 22 0.855 22.1 2.2 ;
 RECT 24.865 1.125 24.965 2.2 ;
 RECT 21.035 0.755 22.57 0.84 ;
 RECT 21.035 0.84 22.565 0.855 ;
 RECT 22.47 0.215 22.57 0.755 ;
 RECT 21.035 0.595 21.265 0.755 ;
 RECT 22 2.2 24.965 2.3 ;
 RECT 23.69 1.06 23.79 1.14 ;
 RECT 23.69 0.38 23.79 0.96 ;
 RECT 23.69 1.14 23.96 1.24 ;
 RECT 23.86 1.24 23.96 1.84 ;
 RECT 23.27 0.935 23.5 0.96 ;
 RECT 23.27 0.96 23.79 1.06 ;
 RECT 23.27 1.06 23.5 1.145 ;
 RECT 24.055 0.22 24.285 0.28 ;
 RECT 24.055 0.38 24.285 0.43 ;
 RECT 23.69 0.28 24.285 0.38 ;
 RECT 7.945 1.575 8.045 2.485 ;
 RECT 8.455 1.575 8.685 1.685 ;
 RECT 7.945 1.475 8.685 1.575 ;
 RECT 25.875 0.195 25.975 2.665 ;
 RECT 24.865 0.095 25.975 0.195 ;
 RECT 21.24 1.245 21.34 2.665 ;
 RECT 24.865 0.195 24.965 0.945 ;
 RECT 21.24 1.2 21.525 1.245 ;
 RECT 21.295 1.035 21.525 1.1 ;
 RECT 21.24 2.665 25.975 2.765 ;
 RECT 21.24 1.1 21.57 1.2 ;
 RECT 12.17 0.795 12.335 0.925 ;
 RECT 11.49 0.885 11.72 0.925 ;
 RECT 11.49 1.025 11.72 1.095 ;
 RECT 11.49 0.925 12.335 1.025 ;
 RECT 12.17 0.585 12.4 0.795 ;
 RECT 3.27 0.705 3.37 1.165 ;
 RECT 2.83 1.27 2.93 1.445 ;
 RECT 3.27 0.47 3.555 0.705 ;
 RECT 2.83 1.17 3.37 1.265 ;
 RECT 2.83 1.265 3.205 1.27 ;
 RECT 3.06 1.165 3.37 1.17 ;
 RECT 2.685 1.445 2.93 1.69 ;
 RECT 4.16 0.715 4.26 1.61 ;
 RECT 4.195 1.71 4.295 2.48 ;
 RECT 4.16 1.61 4.295 1.71 ;
 RECT 4.04 0.485 4.28 0.715 ;
 RECT 0.85 0.27 1.19 0.52 ;
 RECT 1.09 0.52 1.19 2.465 ;
 RECT 9.765 0.655 9.865 1.155 ;
 RECT 9.355 1.255 9.585 1.44 ;
 RECT 9.355 1.155 9.865 1.255 ;
 RECT 1.565 0.49 1.665 1.495 ;
 RECT 1.37 1.495 1.665 1.745 ;
 RECT 1.565 1.745 1.665 2.37 ;
 RECT 3.72 1.33 3.86 1.475 ;
 RECT 3.72 1.71 3.82 2.475 ;
 RECT 3.76 0.65 3.86 1.33 ;
 RECT 3.72 1.475 3.95 1.71 ;
 RECT 8.87 0.655 8.97 1.18 ;
 RECT 8.87 1.28 8.97 1.655 ;
 RECT 7.955 0.66 8.055 1.18 ;
 RECT 8.87 1.655 9.83 1.755 ;
 RECT 9.73 1.755 9.83 2.255 ;
 RECT 8.87 1.755 8.97 2.51 ;
 RECT 9.73 2.255 9.965 2.355 ;
 RECT 9.735 2.355 9.965 2.465 ;
 RECT 7.955 1.18 8.97 1.28 ;
 RECT 15.72 0.55 15.82 2.69 ;
 RECT 6.65 1.58 6.75 2.69 ;
 RECT 6.39 1.01 6.49 1.48 ;
 RECT 7.25 2.445 7.48 2.69 ;
 RECT 6.39 1.48 6.75 1.58 ;
 RECT 6.65 2.69 15.82 2.79 ;
 RECT 19.07 0.49 19.17 1.275 ;
 RECT 19.65 0.385 19.75 1.275 ;
 RECT 19.65 1.375 19.75 2.73 ;
 RECT 19.07 1.375 19.17 2.74 ;
 RECT 18.27 0.49 18.5 0.62 ;
 RECT 18.27 0.39 19.17 0.49 ;
 RECT 19.07 1.275 19.75 1.375 ;
 RECT 16.825 0.43 16.925 1.245 ;
 RECT 16.775 1.245 17.005 1.455 ;
 RECT 16.76 0.22 16.99 0.43 ;
 RECT 4.98 2.445 5.24 2.655 ;
 RECT 5.14 1.79 5.24 2.445 ;
 RECT 15.25 1.445 15.35 2.035 ;
 RECT 15.235 2.035 15.465 2.245 ;
 RECT 6.09 0.98 6.19 1.615 ;
 RECT 5.95 1.615 6.19 1.825 ;
 LAYER CO ;
 RECT 0.84 0.74 0.97 0.87 ;
 RECT 2.56 1.825 2.69 1.955 ;
 RECT 10.42 1.945 10.55 2.075 ;
 RECT 1.31 2.05 1.44 2.18 ;
 RECT 21.5 0.505 21.63 0.635 ;
 RECT 7.695 2.015 7.825 2.145 ;
 RECT 23.435 0.12 23.565 0.25 ;
 RECT 23 1.485 23.13 1.615 ;
 RECT 25.395 1.465 25.525 1.595 ;
 RECT 15.94 1.705 16.07 1.835 ;
 RECT 25.395 0.595 25.525 0.725 ;
 RECT 3.77 1.525 3.9 1.655 ;
 RECT 9.32 2.225 9.45 2.355 ;
 RECT 19.29 2.64 19.42 2.77 ;
 RECT 0.84 2.115 0.97 2.245 ;
 RECT 19.875 0.63 20.005 0.76 ;
 RECT 23.94 0.595 24.07 0.725 ;
 RECT 3.375 0.525 3.505 0.655 ;
 RECT 4.42 1.825 4.55 1.955 ;
 RECT 16.415 1.705 16.545 1.835 ;
 RECT 24.08 1.405 24.21 1.535 ;
 RECT 7.7 0.905 7.83 1.035 ;
 RECT 0.91 0.325 1.04 0.455 ;
 RECT 5.84 0.315 5.97 0.445 ;
 RECT 8.175 0.905 8.305 1.035 ;
 RECT 11.45 0.595 11.58 0.725 ;
 RECT 9.51 0.62 9.64 0.75 ;
 RECT 23.605 1.445 23.735 1.575 ;
 RECT 0.34 1.825 0.47 1.955 ;
 RECT 14.475 1.035 14.605 1.165 ;
 RECT 15.06 0.91 15.19 1.04 ;
 RECT 6.87 2.11 7 2.24 ;
 RECT 19.375 0.62 19.505 0.75 ;
 RECT 5.36 2.135 5.49 2.265 ;
 RECT 2.975 2.105 3.105 2.235 ;
 RECT 3.94 2.11 4.07 2.24 ;
 RECT 1.895 0.145 2.025 0.275 ;
 RECT 10.945 1.9 11.075 2.03 ;
 RECT 0.34 2.345 0.47 2.475 ;
 RECT 2.05 2.345 2.18 2.475 ;
 RECT 23 0.435 23.13 0.565 ;
 RECT 6.65 1.23 6.78 1.36 ;
 RECT 15.47 1.705 15.6 1.835 ;
 RECT 5.84 2.075 5.97 2.205 ;
 RECT 3.49 0.88 3.62 1.01 ;
 RECT 9.785 2.295 9.915 2.425 ;
 RECT 7.3 2.485 7.43 2.615 ;
 RECT 18.32 0.45 18.45 0.58 ;
 RECT 16.825 1.285 16.955 1.415 ;
 RECT 14.645 0.43 14.775 0.56 ;
 RECT 16.265 0.6 16.395 0.73 ;
 RECT 16.81 0.26 16.94 0.39 ;
 RECT 5.03 2.485 5.16 2.615 ;
 RECT 15.285 2.075 15.415 2.205 ;
 RECT 6 1.655 6.13 1.785 ;
 RECT 20.305 0.26 20.435 0.39 ;
 RECT 25.245 1.03 25.375 1.16 ;
 RECT 12.945 0.495 13.075 0.625 ;
 RECT 14.135 1.43 14.265 1.56 ;
 RECT 12.22 0.625 12.35 0.755 ;
 RECT 12.14 1.445 12.27 1.575 ;
 RECT 22.395 1.075 22.525 1.205 ;
 RECT 7.27 0.935 7.4 1.065 ;
 RECT 23.32 0.975 23.45 1.105 ;
 RECT 13.8 0.665 13.93 0.795 ;
 RECT 22.84 1.035 22.97 1.165 ;
 RECT 25.28 2.31 25.41 2.44 ;
 RECT 10.515 2.34 10.645 2.47 ;
 RECT 21.085 0.635 21.215 0.765 ;
 RECT 24.105 0.26 24.235 0.39 ;
 RECT 8.505 1.515 8.635 1.645 ;
 RECT 21.345 1.075 21.475 1.205 ;
 RECT 11.54 0.925 11.67 1.055 ;
 RECT 24.45 1.49 24.58 1.62 ;
 RECT 3.02 0.88 3.15 1.01 ;
 RECT 11.45 1.87 11.58 2 ;
 RECT 4.89 2.11 5.02 2.24 ;
 RECT 4.705 0.32 4.835 0.45 ;
 RECT 22.22 0.135 22.35 0.265 ;
 RECT 1.965 1.495 2.095 1.625 ;
 RECT 1.915 0.745 2.045 0.875 ;
 RECT 1.785 1.995 1.915 2.125 ;
 RECT 8.62 1.995 8.75 2.125 ;
 RECT 0.34 0.59 0.47 0.72 ;
 RECT 8.175 2.07 8.305 2.2 ;
 RECT 10.945 0.595 11.075 0.725 ;
 RECT 2.74 1.49 2.87 1.62 ;
 RECT 9.405 1.245 9.535 1.375 ;
 RECT 18.815 1.725 18.945 1.855 ;
 RECT 0.34 2.085 0.47 2.215 ;
 RECT 6.38 2.045 6.51 2.175 ;
 RECT 1.43 1.55 1.56 1.68 ;
 RECT 13.5 1.835 13.63 1.965 ;
 RECT 13.37 0.765 13.5 0.895 ;
 RECT 1.31 0.74 1.44 0.87 ;
 RECT 24.615 0.12 24.745 0.25 ;
 RECT 4.095 0.53 4.225 0.66 ;
 RECT 18.815 0.85 18.945 0.98 ;
 RECT 12.345 2.38 12.475 2.51 ;
 RECT 8.62 0.905 8.75 1.035 ;
 RECT 21.75 1.425 21.88 1.555 ;
 RECT 0.34 0.33 0.47 0.46 ;
 RECT 16.535 0.92 16.665 1.05 ;
 RECT 22.22 1.475 22.35 1.605 ;
 RECT 10.42 0.875 10.55 1.005 ;
 RECT 2.625 0.79 2.755 0.92 ;
 RECT 14.44 1.835 14.57 1.965 ;
 RECT 3.47 2.07 3.6 2.2 ;
 RECT 26.175 1.475 26.305 1.605 ;
 RECT 19.875 1.71 20.005 1.84 ;
 LAYER M1 ;
 RECT 8.615 1.685 9.185 1.775 ;
 RECT 8.455 1.635 9.185 1.685 ;
 RECT 9.045 1.24 9.585 1.38 ;
 RECT 3.87 2.105 5.09 2.245 ;
 RECT 6.375 1.365 6.515 2.25 ;
 RECT 4.43 1.365 4.57 1.5 ;
 RECT 3.6 1.64 4.105 1.675 ;
 RECT 3.6 1.5 4.57 1.64 ;
 RECT 4.43 1.225 7.08 1.25 ;
 RECT 7.69 1.04 7.83 1.25 ;
 RECT 7.69 1.39 7.83 2.215 ;
 RECT 7.69 0.885 7.83 0.9 ;
 RECT 4.43 1.25 7.83 1.365 ;
 RECT 6.94 1.365 7.83 1.39 ;
 RECT 7.625 0.9 7.9 1.04 ;
 RECT 23.935 0.73 24.075 1.04 ;
 RECT 24.075 1.18 24.215 1.605 ;
 RECT 23.87 0.59 24.145 0.73 ;
 RECT 25.195 0.99 25.425 1.04 ;
 RECT 23.935 1.04 25.425 1.18 ;
 RECT 25.195 1.18 25.425 1.2 ;
 RECT 24.055 0.29 24.425 0.43 ;
 RECT 24.285 0.43 24.425 0.71 ;
 RECT 24.055 0.22 24.285 0.29 ;
 RECT 25.705 0.85 25.845 1.385 ;
 RECT 25.39 1.525 25.53 1.73 ;
 RECT 24.285 0.71 25.845 0.85 ;
 RECT 25.39 0.51 25.53 0.71 ;
 RECT 25.39 1.385 25.845 1.525 ;
 RECT 21.295 1.225 21.525 1.245 ;
 RECT 21.295 1.195 21.885 1.225 ;
 RECT 21.435 1.015 21.745 1.035 ;
 RECT 21.295 1.035 21.745 1.055 ;
 RECT 21.57 0.64 21.71 1.015 ;
 RECT 21.745 1.225 21.885 1.75 ;
 RECT 21.45 0.5 21.71 0.64 ;
 RECT 22.345 1.035 22.575 1.055 ;
 RECT 22.345 1.195 22.575 1.245 ;
 RECT 21.295 1.055 22.575 1.195 ;
 RECT 23.315 1.145 23.455 1.345 ;
 RECT 22.995 1.485 23.135 1.76 ;
 RECT 23.315 0.73 23.455 0.935 ;
 RECT 22.995 0.355 23.135 0.59 ;
 RECT 22.995 1.345 23.455 1.485 ;
 RECT 23.27 0.935 23.5 1.145 ;
 RECT 22.995 0.59 23.455 0.73 ;
 RECT 20.255 0.36 20.485 0.43 ;
 RECT 21.85 0.36 21.99 0.565 ;
 RECT 20.255 0.22 21.99 0.36 ;
 RECT 22.59 0.705 22.73 0.75 ;
 RECT 22.715 0.995 23.02 1.205 ;
 RECT 22.715 0.89 22.855 0.995 ;
 RECT 22.59 0.75 22.855 0.89 ;
 RECT 21.85 0.565 22.73 0.705 ;
 RECT 14.47 1.545 14.61 1.83 ;
 RECT 14.47 1.17 14.61 1.405 ;
 RECT 13.425 1.83 14.675 1.97 ;
 RECT 14.4 1.03 14.68 1.17 ;
 RECT 15.49 0.775 15.63 1.405 ;
 RECT 16.215 0.56 16.445 0.635 ;
 RECT 14.47 1.405 15.63 1.545 ;
 RECT 15.49 0.635 16.445 0.775 ;
 RECT 14.595 0.28 18.5 0.42 ;
 RECT 18.27 0.42 18.5 0.62 ;
 RECT 14.595 0.42 14.825 0.6 ;
 RECT 16.76 0.22 16.99 0.28 ;
 RECT 16.76 0.42 16.99 0.43 ;
 RECT 11.445 0.525 11.585 0.885 ;
 RECT 11.445 1.095 11.585 2.065 ;
 RECT 11.445 0.885 11.72 1.095 ;
 RECT 8.965 2.055 9.105 2.34 ;
 RECT 8.17 2.34 9.105 2.48 ;
 RECT 9.325 1.66 9.465 1.915 ;
 RECT 8.965 1.915 9.465 2.055 ;
 RECT 8.17 1.04 8.31 2.34 ;
 RECT 8.17 0.895 8.31 0.9 ;
 RECT 8.1 0.9 8.375 1.04 ;
 RECT 9.325 1.52 11.08 1.66 ;
 RECT 10.94 0.525 11.08 1.52 ;
 RECT 10.94 1.66 11.08 2.11 ;
 RECT 10.415 0.765 10.555 1.52 ;
 RECT 10.415 1.66 10.555 2.145 ;
 RECT 12.17 0.585 13.125 0.63 ;
 RECT 12.895 0.63 13.125 0.665 ;
 RECT 12.895 0.455 13.125 0.49 ;
 RECT 12.195 0.49 13.125 0.585 ;
 RECT 12.17 0.63 12.4 0.795 ;
 RECT 13.75 0.57 13.98 0.95 ;
 RECT 0.615 1.335 0.755 2.11 ;
 RECT 0.615 2.25 0.755 2.255 ;
 RECT 0.615 0.875 0.755 1.195 ;
 RECT 0.615 2.11 1.04 2.25 ;
 RECT 0.615 0.735 1.04 0.875 ;
 RECT 0.615 1.195 1.725 1.335 ;
 RECT 1.585 0.6 1.725 1.195 ;
 RECT 3.015 0.36 3.155 2.035 ;
 RECT 2.33 0.36 2.47 0.46 ;
 RECT 2.33 0.22 3.155 0.36 ;
 RECT 2.97 2.17 3.11 2.305 ;
 RECT 1.585 0.46 2.47 0.6 ;
 RECT 2.97 2.035 3.155 2.17 ;
 RECT 3.765 0.66 3.905 0.895 ;
 RECT 3.305 0.52 3.905 0.66 ;
 RECT 3.765 0.895 7.45 1.035 ;
 RECT 7.22 1.035 7.45 1.105 ;
 RECT 1.865 0.88 2.005 1.475 ;
 RECT 1.825 1.63 1.965 1.99 ;
 RECT 1.825 1.475 2.17 1.63 ;
 RECT 1.715 1.99 1.965 2.13 ;
 RECT 1.865 0.74 2.185 0.88 ;
 RECT 3.31 1.82 4.89 1.96 ;
 RECT 4.75 1.79 4.89 1.82 ;
 RECT 3.395 1.96 3.675 2.215 ;
 RECT 3.485 0.805 3.625 1.22 ;
 RECT 3.31 1.22 3.625 1.36 ;
 RECT 3.31 1.36 3.45 1.82 ;
 RECT 5.95 1.615 6.18 1.65 ;
 RECT 5.95 1.79 6.18 1.825 ;
 RECT 4.75 1.65 6.185 1.79 ;
 RECT 2.62 1.67 2.76 1.82 ;
 RECT 2.62 1.96 2.76 2.51 ;
 RECT 2.62 0.5 2.76 1.44 ;
 RECT 2.62 1.44 2.875 1.67 ;
 RECT 2.49 1.82 2.76 1.96 ;
 RECT 4.98 2.445 5.21 2.51 ;
 RECT 4.98 2.65 5.21 2.655 ;
 RECT 2.62 2.51 5.21 2.65 ;
 RECT 16.3 1.7 16.595 1.84 ;
 RECT 16.3 1.84 16.44 2.075 ;
 RECT 15.605 1.84 15.745 2.075 ;
 RECT 15.41 1.7 15.745 1.84 ;
 RECT 15.605 2.075 16.44 2.215 ;
 RECT 16.495 1.055 16.635 1.245 ;
 RECT 15.935 1.385 16.075 1.625 ;
 RECT 16.775 1.385 17.005 1.455 ;
 RECT 15.935 1.245 17.005 1.385 ;
 RECT 16.465 0.915 16.765 1.055 ;
 RECT 15.905 1.625 16.16 1.92 ;
 RECT 13.14 1.56 13.28 2.11 ;
 RECT 12.09 1.405 12.32 1.42 ;
 RECT 12.09 1.56 12.32 1.615 ;
 RECT 12.09 1.42 13.28 1.56 ;
 RECT 13.14 2.11 15.465 2.245 ;
 RECT 13.14 2.245 15.46 2.25 ;
 RECT 15.235 2.035 15.465 2.11 ;
 RECT 17.005 2.205 17.145 2.39 ;
 RECT 12.86 1.895 13 2.39 ;
 RECT 12.86 2.39 17.145 2.53 ;
 RECT 11.735 1.755 13 1.895 ;
 RECT 11.735 1.895 11.875 2.34 ;
 RECT 10.465 2.3 10.695 2.34 ;
 RECT 10.465 2.48 10.695 2.51 ;
 RECT 10.465 2.34 11.875 2.48 ;
 RECT 17.005 2.065 21.03 2.205 ;
 RECT 20.89 2.205 21.03 2.52 ;
 RECT 25.23 2.48 25.37 2.52 ;
 RECT 20.89 2.52 25.37 2.66 ;
 RECT 25.23 2.27 25.46 2.48 ;
 RECT 8.615 1.04 8.755 1.475 ;
 RECT 8.455 1.475 8.755 1.635 ;
 RECT 8.615 1.775 8.755 2.18 ;
 RECT 8.545 0.9 8.82 1.04 ;
 RECT 9.045 1.38 9.185 1.635 ;
 END
END RDFFNSRASRNX1

MACRO RDFFNSRASRNX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.84 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.895 0.59 21.265 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.125 1.435 26.465 1.8 ;
 RECT 24.445 1.99 26.31 2.13 ;
 RECT 22.215 2.22 24.585 2.36 ;
 RECT 26.17 1.8 26.31 1.99 ;
 RECT 24.445 1.435 24.585 1.99 ;
 RECT 22.215 1.39 22.355 2.22 ;
 RECT 23.6 1.37 23.74 2.22 ;
 RECT 24.445 2.13 24.585 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.8 0.22 1.165 0.525 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.825 0.08 2.105 0.295 ;
 RECT 24.565 0.08 24.805 0.26 ;
 RECT 5.755 0.31 6.045 0.45 ;
 RECT 13.365 0.275 14.39 0.415 ;
 RECT 9.44 0.615 9.71 0.755 ;
 RECT 14.25 0.75 15.195 0.89 ;
 RECT 0 -0.08 27.84 0.08 ;
 RECT 1.305 0.08 1.445 0.97 ;
 RECT 4.65 0.08 4.885 0.46 ;
 RECT 0.335 0.08 0.475 0.775 ;
 RECT 18.325 0.08 18.465 0.82 ;
 RECT 19.37 0.08 19.51 0.82 ;
 RECT 22.215 0.08 22.355 0.36 ;
 RECT 23.43 0.08 23.57 0.35 ;
 RECT 5.835 0.08 5.975 0.31 ;
 RECT 13.365 0.415 13.505 0.945 ;
 RECT 13.365 0.08 13.505 0.275 ;
 RECT 9.505 0.08 9.645 0.615 ;
 RECT 15.055 0.89 15.195 1.11 ;
 RECT 14.25 0.415 14.39 0.75 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 18.225 2.6 18.49 2.8 ;
 RECT 19.225 2.6 19.49 2.8 ;
 RECT 9.25 2.215 9.525 2.355 ;
 RECT 0 2.8 27.84 2.96 ;
 RECT 1.98 2.34 2.23 2.8 ;
 RECT 0.335 1.74 0.475 2.8 ;
 RECT 1.305 1.98 1.445 2.8 ;
 RECT 5.355 2.07 5.495 2.8 ;
 RECT 5.835 1.98 5.975 2.8 ;
 RECT 6.865 2 7.005 2.8 ;
 RECT 12.275 2.335 12.545 2.8 ;
 RECT 9.315 2.355 9.455 2.8 ;
 RECT 9.315 2.195 9.455 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.355 1.475 1.685 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.87 1.095 20.24 1.335 ;
 RECT 19.87 0.56 20.01 1.095 ;
 RECT 17.76 1.905 17.9 1.915 ;
 RECT 17.76 0.51 17.9 1.765 ;
 RECT 18.81 1.905 18.95 1.915 ;
 RECT 18.81 0.51 18.95 1.765 ;
 RECT 19.87 1.905 20.01 1.91 ;
 RECT 17.725 1.765 20.01 1.905 ;
 RECT 19.87 1.335 20.01 1.765 ;
 END
 ANTENNADIFFAREA 1.102 ;
 END QN

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.73 2.255 10.045 2.465 ;
 RECT 9.765 2.12 10.045 2.255 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.045 0.485 4.36 0.605 ;
 RECT 8.965 0.905 10.02 1.045 ;
 RECT 9.875 0.245 12.025 0.255 ;
 RECT 9.875 0.255 12.03 0.385 ;
 RECT 11.89 1.09 13.88 1.23 ;
 RECT 14.085 1.56 14.315 1.6 ;
 RECT 13.74 1.42 14.315 1.56 ;
 RECT 14.085 1.39 14.315 1.42 ;
 RECT 4.045 0.605 9.105 0.745 ;
 RECT 8.965 0.745 9.105 0.905 ;
 RECT 9.88 0.385 10.02 0.905 ;
 RECT 11.89 0.385 12.03 1.09 ;
 RECT 13.74 1.23 13.88 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.24 2.12 7.48 2.66 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 OBS
 LAYER PO ;
 RECT 6.09 0.98 6.19 1.615 ;
 RECT 5.95 1.615 6.19 1.825 ;
 RECT 6.09 1.825 6.19 2.51 ;
 RECT 20.255 0.195 20.355 0.22 ;
 RECT 16.19 0.095 20.355 0.195 ;
 RECT 16.19 0.77 16.29 2.155 ;
 RECT 16.19 0.195 16.29 0.56 ;
 RECT 16.19 0.56 16.445 0.77 ;
 RECT 16.19 0.09 16.29 0.095 ;
 RECT 20.255 0.22 20.485 0.43 ;
 RECT 14.22 0.73 14.32 1.39 ;
 RECT 14.085 1.39 14.32 1.6 ;
 RECT 14.22 1.6 14.32 2.39 ;
 RECT 2.405 0.285 2.505 1.52 ;
 RECT 1.905 1.52 2.505 1.62 ;
 RECT 2.405 0.185 11.295 0.195 ;
 RECT 4.46 0.095 11.295 0.185 ;
 RECT 2.405 0.195 4.56 0.285 ;
 RECT 11.195 0.195 11.295 1.29 ;
 RECT 12.09 1.39 12.285 1.405 ;
 RECT 3.225 1.565 3.325 2.675 ;
 RECT 2.34 1.62 2.44 2.675 ;
 RECT 1.905 1.44 2.15 1.52 ;
 RECT 1.905 1.62 2.15 1.69 ;
 RECT 4.46 0.285 4.56 1.24 ;
 RECT 11.195 1.29 12.285 1.39 ;
 RECT 2.34 2.675 3.325 2.775 ;
 RECT 12.09 1.405 12.32 1.615 ;
 RECT 22.475 1.245 22.575 2.02 ;
 RECT 22.345 1.035 22.575 1.245 ;
 RECT 12.585 0.105 15.41 0.205 ;
 RECT 12.585 0.205 12.685 1.91 ;
 RECT 15.31 0.205 15.41 1.265 ;
 RECT 11.765 1.71 11.865 1.91 ;
 RECT 10.68 1.61 11.865 1.71 ;
 RECT 10.68 0.475 10.78 1.61 ;
 RECT 11.23 1.71 11.33 2.425 ;
 RECT 7.345 0.475 7.445 0.895 ;
 RECT 11.765 1.91 12.685 2.01 ;
 RECT 7.345 0.375 10.78 0.475 ;
 RECT 7.22 0.895 7.45 1.105 ;
 RECT 12.895 0.455 14.825 0.535 ;
 RECT 14.595 0.535 14.825 0.6 ;
 RECT 14.595 0.39 14.825 0.435 ;
 RECT 12.975 0.435 14.825 0.455 ;
 RECT 12.895 0.535 13.125 0.665 ;
 RECT 13.75 0.535 13.98 0.835 ;
 RECT 13.75 0.835 13.85 2.39 ;
 RECT 22.78 0.215 22.88 0.995 ;
 RECT 22.78 0.995 23.02 1.205 ;
 RECT 22.78 1.205 22.88 2 ;
 RECT 25.175 0.375 25.275 0.99 ;
 RECT 25.175 0.99 25.425 1.2 ;
 RECT 25.175 1.2 25.275 2.27 ;
 RECT 25.175 2.27 25.46 2.48 ;
 RECT 10.16 0.655 10.26 2.305 ;
 RECT 10.465 2.3 10.695 2.305 ;
 RECT 10.465 2.405 10.695 2.51 ;
 RECT 10.16 2.305 10.695 2.405 ;
 RECT 22 0.21 22.1 0.755 ;
 RECT 22 0.855 22.1 2.2 ;
 RECT 24.865 1.125 24.965 2.2 ;
 RECT 21.035 0.755 22.57 0.84 ;
 RECT 21.035 0.84 22.565 0.855 ;
 RECT 22.47 0.215 22.57 0.755 ;
 RECT 21.035 0.595 21.265 0.755 ;
 RECT 22 2.2 24.965 2.3 ;
 RECT 23.69 1.06 23.79 1.14 ;
 RECT 23.69 0.38 23.79 0.96 ;
 RECT 23.69 1.14 23.96 1.24 ;
 RECT 23.86 1.24 23.96 1.84 ;
 RECT 23.27 0.935 23.5 0.96 ;
 RECT 23.27 0.96 23.79 1.06 ;
 RECT 23.27 1.06 23.5 1.145 ;
 RECT 24.055 0.22 24.285 0.28 ;
 RECT 24.055 0.38 24.285 0.43 ;
 RECT 23.69 0.28 24.285 0.38 ;
 RECT 7.945 1.575 8.045 2.485 ;
 RECT 8.455 1.575 8.685 1.685 ;
 RECT 7.945 1.475 8.685 1.575 ;
 RECT 25.875 0.195 25.975 2.665 ;
 RECT 24.865 0.095 25.975 0.195 ;
 RECT 21.24 1.245 21.34 2.665 ;
 RECT 24.865 0.195 24.965 0.945 ;
 RECT 21.24 1.2 21.525 1.245 ;
 RECT 21.295 1.035 21.525 1.1 ;
 RECT 21.24 2.665 25.975 2.765 ;
 RECT 21.24 1.1 21.57 1.2 ;
 RECT 12.17 0.795 12.335 0.925 ;
 RECT 11.49 0.885 11.72 0.925 ;
 RECT 11.49 1.025 11.72 1.095 ;
 RECT 11.49 0.925 12.335 1.025 ;
 RECT 12.17 0.585 12.4 0.795 ;
 RECT 3.27 0.705 3.37 1.165 ;
 RECT 2.83 1.27 2.93 1.445 ;
 RECT 3.27 0.47 3.555 0.705 ;
 RECT 2.83 1.17 3.37 1.265 ;
 RECT 2.83 1.265 3.205 1.27 ;
 RECT 3.06 1.165 3.37 1.17 ;
 RECT 2.685 1.445 2.93 1.69 ;
 RECT 4.16 0.715 4.26 1.61 ;
 RECT 4.195 1.71 4.295 2.48 ;
 RECT 4.16 1.61 4.295 1.71 ;
 RECT 4.04 0.485 4.28 0.715 ;
 RECT 9.765 0.655 9.865 1.155 ;
 RECT 9.15 1.255 9.38 1.475 ;
 RECT 9.15 1.155 9.865 1.255 ;
 RECT 1.565 0.49 1.665 1.495 ;
 RECT 1.37 1.495 1.665 1.745 ;
 RECT 1.565 1.745 1.665 2.37 ;
 RECT 3.72 1.33 3.86 1.475 ;
 RECT 3.72 1.71 3.82 2.475 ;
 RECT 3.76 0.65 3.86 1.33 ;
 RECT 3.72 1.475 3.95 1.71 ;
 RECT 1.09 0.52 1.19 2.465 ;
 RECT 0.85 0.27 1.19 0.52 ;
 RECT 15.72 0.55 15.82 2.69 ;
 RECT 6.65 1.58 6.75 2.69 ;
 RECT 6.39 1.01 6.49 1.48 ;
 RECT 7.245 2.45 7.475 2.69 ;
 RECT 6.39 1.48 6.75 1.58 ;
 RECT 6.65 2.69 15.82 2.79 ;
 RECT 8.87 0.655 8.97 1.18 ;
 RECT 8.87 1.28 8.97 1.655 ;
 RECT 7.955 0.66 8.055 1.18 ;
 RECT 8.87 1.655 9.83 1.755 ;
 RECT 9.73 1.755 9.83 2.255 ;
 RECT 8.87 1.755 8.97 2.51 ;
 RECT 7.955 1.18 8.97 1.28 ;
 RECT 9.73 2.255 9.96 2.465 ;
 RECT 16.775 1.33 19.75 1.43 ;
 RECT 16.825 0.615 16.925 1.245 ;
 RECT 19.65 0.385 19.75 1.33 ;
 RECT 19.65 1.43 19.75 2.73 ;
 RECT 19.07 0.385 19.17 1.33 ;
 RECT 19.07 1.43 19.17 2.74 ;
 RECT 18.595 1.43 18.695 2.73 ;
 RECT 18.595 0.385 18.695 1.33 ;
 RECT 18.015 0.385 18.115 1.33 ;
 RECT 18.015 1.43 18.115 2.74 ;
 RECT 16.775 1.245 17.005 1.33 ;
 RECT 16.775 1.43 17.005 1.455 ;
 RECT 16.76 0.405 16.99 0.615 ;
 RECT 4.98 2.445 5.24 2.655 ;
 RECT 5.14 1.79 5.24 2.445 ;
 RECT 15.25 1.445 15.35 2.035 ;
 RECT 15.235 2.035 15.465 2.245 ;
 LAYER CO ;
 RECT 7.695 2.015 7.825 2.145 ;
 RECT 23.435 0.12 23.565 0.25 ;
 RECT 23 1.485 23.13 1.615 ;
 RECT 25.395 1.465 25.525 1.595 ;
 RECT 15.94 1.705 16.07 1.835 ;
 RECT 25.395 0.595 25.525 0.725 ;
 RECT 3.77 1.525 3.9 1.655 ;
 RECT 9.32 2.225 9.45 2.355 ;
 RECT 19.29 2.64 19.42 2.77 ;
 RECT 0.84 2.115 0.97 2.245 ;
 RECT 19.875 0.63 20.005 0.76 ;
 RECT 23.94 0.595 24.07 0.725 ;
 RECT 3.375 0.525 3.505 0.655 ;
 RECT 4.42 1.825 4.55 1.955 ;
 RECT 24.45 1.49 24.58 1.62 ;
 RECT 3.02 0.88 3.15 1.01 ;
 RECT 11.45 1.87 11.58 2 ;
 RECT 4.89 2.11 5.02 2.24 ;
 RECT 4.705 0.32 4.835 0.45 ;
 RECT 16.415 1.705 16.545 1.835 ;
 RECT 24.08 1.405 24.21 1.535 ;
 RECT 7.7 0.905 7.83 1.035 ;
 RECT 0.91 0.325 1.04 0.455 ;
 RECT 5.84 0.315 5.97 0.445 ;
 RECT 8.175 0.905 8.305 1.035 ;
 RECT 11.45 0.595 11.58 0.725 ;
 RECT 9.51 0.62 9.64 0.75 ;
 RECT 23.605 1.445 23.735 1.575 ;
 RECT 0.34 1.825 0.47 1.955 ;
 RECT 14.475 1.035 14.605 1.165 ;
 RECT 15.06 0.91 15.19 1.04 ;
 RECT 6.87 2.11 7 2.24 ;
 RECT 19.375 0.62 19.505 0.75 ;
 RECT 5.36 2.135 5.49 2.265 ;
 RECT 2.975 2.105 3.105 2.235 ;
 RECT 3.94 2.11 4.07 2.24 ;
 RECT 1.895 0.145 2.025 0.275 ;
 RECT 10.945 1.9 11.075 2.03 ;
 RECT 0.34 2.345 0.47 2.475 ;
 RECT 2.05 2.345 2.18 2.475 ;
 RECT 23 0.435 23.13 0.565 ;
 RECT 6.65 1.23 6.78 1.36 ;
 RECT 15.47 1.705 15.6 1.835 ;
 RECT 5.84 2.075 5.97 2.205 ;
 RECT 3.49 0.88 3.62 1.01 ;
 RECT 13.5 1.835 13.63 1.965 ;
 RECT 7.295 2.49 7.425 2.62 ;
 RECT 9.78 2.295 9.91 2.425 ;
 RECT 16.825 1.285 16.955 1.415 ;
 RECT 14.645 0.43 14.775 0.56 ;
 RECT 16.265 0.6 16.395 0.73 ;
 RECT 16.81 0.445 16.94 0.575 ;
 RECT 5.03 2.485 5.16 2.615 ;
 RECT 15.285 2.075 15.415 2.205 ;
 RECT 6 1.655 6.13 1.785 ;
 RECT 20.305 0.26 20.435 0.39 ;
 RECT 25.245 1.03 25.375 1.16 ;
 RECT 12.945 0.495 13.075 0.625 ;
 RECT 14.135 1.43 14.265 1.56 ;
 RECT 12.22 0.625 12.35 0.755 ;
 RECT 12.14 1.445 12.27 1.575 ;
 RECT 22.395 1.075 22.525 1.205 ;
 RECT 7.27 0.935 7.4 1.065 ;
 RECT 23.32 0.975 23.45 1.105 ;
 RECT 13.8 0.665 13.93 0.795 ;
 RECT 22.84 1.035 22.97 1.165 ;
 RECT 25.28 2.31 25.41 2.44 ;
 RECT 10.515 2.34 10.645 2.47 ;
 RECT 21.085 0.635 21.215 0.765 ;
 RECT 24.105 0.26 24.235 0.39 ;
 RECT 8.505 1.515 8.635 1.645 ;
 RECT 21.345 1.075 21.475 1.205 ;
 RECT 11.54 0.925 11.67 1.055 ;
 RECT 22.22 0.135 22.35 0.265 ;
 RECT 1.965 1.495 2.095 1.625 ;
 RECT 1.915 0.745 2.045 0.875 ;
 RECT 1.785 1.995 1.915 2.125 ;
 RECT 8.62 1.995 8.75 2.125 ;
 RECT 0.34 0.59 0.47 0.72 ;
 RECT 8.175 2.07 8.305 2.2 ;
 RECT 10.945 0.595 11.075 0.725 ;
 RECT 2.74 1.49 2.87 1.62 ;
 RECT 9.2 1.28 9.33 1.41 ;
 RECT 18.815 1.725 18.945 1.855 ;
 RECT 0.34 2.085 0.47 2.215 ;
 RECT 6.38 2.045 6.51 2.175 ;
 RECT 1.43 1.55 1.56 1.68 ;
 RECT 18.29 2.64 18.42 2.77 ;
 RECT 18.33 0.62 18.46 0.75 ;
 RECT 17.765 1.725 17.895 1.855 ;
 RECT 17.765 0.62 17.895 0.75 ;
 RECT 13.37 0.765 13.5 0.895 ;
 RECT 1.31 0.74 1.44 0.87 ;
 RECT 24.615 0.12 24.745 0.25 ;
 RECT 4.095 0.53 4.225 0.66 ;
 RECT 18.815 0.62 18.945 0.75 ;
 RECT 12.345 2.38 12.475 2.51 ;
 RECT 8.62 0.905 8.75 1.035 ;
 RECT 21.75 1.425 21.88 1.555 ;
 RECT 0.34 0.33 0.47 0.46 ;
 RECT 16.535 0.92 16.665 1.05 ;
 RECT 22.22 1.475 22.35 1.605 ;
 RECT 10.42 0.875 10.55 1.005 ;
 RECT 2.625 0.79 2.755 0.92 ;
 RECT 14.44 1.835 14.57 1.965 ;
 RECT 3.47 2.07 3.6 2.2 ;
 RECT 26.175 1.475 26.305 1.605 ;
 RECT 19.875 1.71 20.005 1.84 ;
 RECT 0.84 0.74 0.97 0.87 ;
 RECT 2.56 1.825 2.69 1.955 ;
 RECT 10.42 1.945 10.55 2.075 ;
 RECT 1.31 2.05 1.44 2.18 ;
 RECT 21.5 0.505 21.63 0.635 ;
 LAYER M1 ;
 RECT 8.545 0.9 8.82 1.04 ;
 RECT 8.615 1.685 9.335 1.775 ;
 RECT 8.455 1.635 9.335 1.685 ;
 RECT 9.195 1.205 9.335 1.635 ;
 RECT 3.87 2.105 5.09 2.245 ;
 RECT 6.375 1.365 6.515 2.25 ;
 RECT 4.43 1.365 4.57 1.5 ;
 RECT 3.6 1.64 4.105 1.675 ;
 RECT 3.6 1.5 4.57 1.64 ;
 RECT 4.43 1.225 7.08 1.25 ;
 RECT 7.69 1.04 7.83 1.25 ;
 RECT 7.69 1.39 7.83 2.215 ;
 RECT 7.69 0.885 7.83 0.9 ;
 RECT 4.43 1.25 7.83 1.365 ;
 RECT 6.94 1.365 7.83 1.39 ;
 RECT 7.625 0.9 7.9 1.04 ;
 RECT 3.31 1.82 4.89 1.96 ;
 RECT 4.75 1.79 4.89 1.82 ;
 RECT 3.395 1.96 3.675 2.215 ;
 RECT 3.485 0.805 3.625 1.22 ;
 RECT 3.31 1.22 3.625 1.36 ;
 RECT 3.31 1.36 3.45 1.82 ;
 RECT 5.95 1.615 6.18 1.65 ;
 RECT 5.95 1.79 6.18 1.825 ;
 RECT 4.75 1.65 6.185 1.79 ;
 RECT 23.935 0.73 24.075 1.04 ;
 RECT 24.075 1.18 24.215 1.605 ;
 RECT 23.87 0.59 24.145 0.73 ;
 RECT 25.195 0.99 25.425 1.04 ;
 RECT 23.935 1.04 25.425 1.18 ;
 RECT 25.195 1.18 25.425 1.2 ;
 RECT 24.055 0.29 24.425 0.43 ;
 RECT 24.285 0.43 24.425 0.71 ;
 RECT 24.055 0.22 24.285 0.29 ;
 RECT 25.705 0.85 25.845 1.385 ;
 RECT 25.39 1.525 25.53 1.73 ;
 RECT 24.285 0.71 25.845 0.85 ;
 RECT 25.39 0.51 25.53 0.71 ;
 RECT 25.39 1.385 25.845 1.525 ;
 RECT 21.295 1.225 21.525 1.245 ;
 RECT 21.295 1.195 21.885 1.225 ;
 RECT 21.435 1.015 21.745 1.035 ;
 RECT 21.295 1.035 21.745 1.055 ;
 RECT 21.57 0.64 21.71 1.015 ;
 RECT 21.745 1.225 21.885 1.75 ;
 RECT 21.45 0.5 21.71 0.64 ;
 RECT 22.345 1.035 22.575 1.055 ;
 RECT 22.345 1.195 22.575 1.245 ;
 RECT 21.295 1.055 22.575 1.195 ;
 RECT 23.315 1.145 23.455 1.345 ;
 RECT 22.995 1.485 23.135 1.76 ;
 RECT 23.315 0.73 23.455 0.935 ;
 RECT 22.995 0.355 23.135 0.59 ;
 RECT 22.995 1.345 23.455 1.485 ;
 RECT 23.27 0.935 23.5 1.145 ;
 RECT 22.995 0.59 23.455 0.73 ;
 RECT 20.255 0.36 20.485 0.43 ;
 RECT 21.85 0.36 21.99 0.565 ;
 RECT 20.255 0.22 21.99 0.36 ;
 RECT 22.59 0.705 22.73 0.75 ;
 RECT 22.715 0.995 23.02 1.205 ;
 RECT 22.715 0.89 22.855 0.995 ;
 RECT 22.59 0.75 22.855 0.89 ;
 RECT 21.85 0.565 22.73 0.705 ;
 RECT 14.47 1.545 14.61 1.83 ;
 RECT 14.47 1.17 14.61 1.405 ;
 RECT 13.425 1.83 14.675 1.97 ;
 RECT 14.4 1.03 14.68 1.17 ;
 RECT 15.49 0.775 15.63 1.405 ;
 RECT 16.215 0.56 16.445 0.635 ;
 RECT 14.47 1.405 15.63 1.545 ;
 RECT 15.49 0.635 16.445 0.775 ;
 RECT 14.595 0.405 16.99 0.42 ;
 RECT 14.595 0.28 16.94 0.405 ;
 RECT 14.595 0.42 14.825 0.6 ;
 RECT 16.76 0.42 16.99 0.615 ;
 RECT 11.445 0.525 11.585 0.885 ;
 RECT 11.445 1.095 11.585 2.065 ;
 RECT 11.445 0.885 11.72 1.095 ;
 RECT 8.965 2.055 9.105 2.34 ;
 RECT 8.17 2.34 9.105 2.48 ;
 RECT 9.48 1.66 9.62 1.915 ;
 RECT 8.965 1.915 9.62 2.055 ;
 RECT 8.17 1.04 8.31 2.34 ;
 RECT 8.17 0.895 8.31 0.9 ;
 RECT 8.1 0.9 8.375 1.04 ;
 RECT 9.48 1.52 11.08 1.66 ;
 RECT 10.94 0.525 11.08 1.52 ;
 RECT 10.94 1.66 11.08 2.11 ;
 RECT 10.415 0.765 10.555 1.52 ;
 RECT 10.415 1.66 10.555 2.145 ;
 RECT 12.17 0.585 13.125 0.63 ;
 RECT 12.895 0.63 13.125 0.665 ;
 RECT 12.895 0.455 13.125 0.49 ;
 RECT 12.195 0.49 13.125 0.585 ;
 RECT 12.17 0.63 12.4 0.795 ;
 RECT 13.75 0.57 13.98 0.95 ;
 RECT 2.62 1.67 2.76 1.82 ;
 RECT 2.62 1.96 2.76 2.51 ;
 RECT 2.62 0.5 2.76 1.44 ;
 RECT 2.62 1.44 2.875 1.67 ;
 RECT 2.49 1.82 2.76 1.96 ;
 RECT 4.98 2.445 5.21 2.51 ;
 RECT 4.98 2.65 5.21 2.655 ;
 RECT 2.62 2.51 5.21 2.65 ;
 RECT 0.615 1.335 0.755 2.11 ;
 RECT 0.615 2.25 0.755 2.255 ;
 RECT 0.615 0.875 0.755 1.195 ;
 RECT 0.615 2.11 1.04 2.25 ;
 RECT 0.615 0.735 1.04 0.875 ;
 RECT 0.615 1.195 1.725 1.335 ;
 RECT 1.585 0.6 1.725 1.195 ;
 RECT 3.015 0.36 3.155 2.035 ;
 RECT 2.33 0.36 2.47 0.46 ;
 RECT 2.33 0.22 3.155 0.36 ;
 RECT 2.97 2.17 3.11 2.305 ;
 RECT 1.585 0.46 2.47 0.6 ;
 RECT 2.97 2.035 3.155 2.17 ;
 RECT 3.765 0.66 3.905 0.895 ;
 RECT 3.305 0.52 3.905 0.66 ;
 RECT 3.765 0.895 7.45 1.035 ;
 RECT 7.22 1.035 7.45 1.105 ;
 RECT 1.865 0.88 2.005 1.475 ;
 RECT 1.825 1.63 1.965 1.99 ;
 RECT 1.825 1.475 2.17 1.63 ;
 RECT 1.715 1.99 1.965 2.13 ;
 RECT 1.865 0.74 2.185 0.88 ;
 RECT 16.3 1.7 16.595 1.84 ;
 RECT 16.3 1.84 16.44 2.075 ;
 RECT 15.605 1.84 15.745 2.075 ;
 RECT 15.41 1.7 15.745 1.84 ;
 RECT 15.605 2.075 16.44 2.215 ;
 RECT 16.495 1.055 16.635 1.245 ;
 RECT 15.935 1.385 16.075 1.625 ;
 RECT 16.775 1.385 17.005 1.455 ;
 RECT 15.935 1.245 17.005 1.385 ;
 RECT 16.465 0.915 16.765 1.055 ;
 RECT 15.905 1.625 16.16 1.92 ;
 RECT 13.14 1.56 13.28 2.11 ;
 RECT 12.09 1.405 12.32 1.42 ;
 RECT 12.09 1.56 12.32 1.615 ;
 RECT 12.09 1.42 13.28 1.56 ;
 RECT 13.14 2.11 15.465 2.245 ;
 RECT 13.14 2.245 15.46 2.25 ;
 RECT 15.235 2.035 15.465 2.11 ;
 RECT 17.005 2.205 17.145 2.39 ;
 RECT 12.86 1.895 13 2.39 ;
 RECT 12.86 2.39 17.145 2.53 ;
 RECT 11.735 1.755 13 1.895 ;
 RECT 11.735 1.895 11.875 2.34 ;
 RECT 10.465 2.3 10.695 2.34 ;
 RECT 10.465 2.48 10.695 2.51 ;
 RECT 10.465 2.34 11.875 2.48 ;
 RECT 17.005 2.065 21.03 2.205 ;
 RECT 20.89 2.205 21.03 2.52 ;
 RECT 25.23 2.48 25.37 2.52 ;
 RECT 20.89 2.52 25.37 2.66 ;
 RECT 25.23 2.27 25.46 2.48 ;
 RECT 8.615 1.775 8.755 2.18 ;
 RECT 8.615 1.04 8.755 1.475 ;
 RECT 8.455 1.475 8.755 1.635 ;
 END
END RDFFNSRASRNX2

MACRO RDFFNX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 20.8 BY 2.88 ;
 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.43 1.145 6.715 1.415 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.3 1.09 9.72 1.5 ;
 RECT 9.3 1.5 9.44 1.855 ;
 RECT 9.3 0.525 9.44 1.09 ;
 END
 ANTENNADIFFAREA 0.626 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.35 1 10.715 1.345 ;
 RECT 10.35 1.345 10.49 1.855 ;
 RECT 10.35 0.48 10.49 1 ;
 END
 ANTENNADIFFAREA 0.604 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 20.8 2.96 ;
 RECT 4.99 2.615 5.225 2.8 ;
 RECT 3.035 2.51 3.265 2.65 ;
 RECT 6.455 2.37 6.725 2.51 ;
 RECT 1.34 2.51 1.61 2.65 ;
 RECT 8.82 2.275 8.96 2.8 ;
 RECT 10.83 2.275 10.97 2.8 ;
 RECT 0.525 1.64 0.685 2.8 ;
 RECT 12.555 2.025 12.695 2.8 ;
 RECT 9.87 2.275 10.01 2.8 ;
 RECT 7.695 1.94 7.835 2.8 ;
 RECT 3.08 2.65 3.22 2.8 ;
 RECT 6.52 2.51 6.66 2.8 ;
 RECT 1.405 2.65 1.545 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 20.8 0.08 ;
 RECT 15.515 0.22 15.765 0.36 ;
 RECT 6.445 0.565 6.715 0.705 ;
 RECT 3.045 0.555 3.295 0.695 ;
 RECT 0.525 0.08 0.685 0.84 ;
 RECT 12.555 0.08 12.695 0.815 ;
 RECT 8.74 0.08 8.88 0.575 ;
 RECT 1.405 0.08 1.545 0.32 ;
 RECT 10.835 0.08 10.975 0.575 ;
 RECT 5.055 0.08 5.195 0.78 ;
 RECT 9.87 0.08 10.01 0.575 ;
 RECT 7.695 0.08 7.835 0.785 ;
 RECT 18.28 0.08 18.42 0.65 ;
 RECT 15.56 0.08 15.7 0.22 ;
 RECT 6.51 0.08 6.65 0.565 ;
 RECT 3.11 0.08 3.25 0.555 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 19.135 1.4 19.475 1.765 ;
 RECT 15.56 2.225 19.3 2.385 ;
 RECT 15.515 1.47 15.745 1.61 ;
 RECT 18.235 1.395 18.375 2.225 ;
 RECT 19.15 1.765 19.29 2.225 ;
 RECT 15.56 1.61 15.7 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.71 0.81 14.09 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.77 0.825 2.17 1.135 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 11.505 0.385 11.605 1.325 ;
 RECT 11.505 1.325 12.14 1.425 ;
 RECT 12.34 0.385 12.44 1.215 ;
 RECT 12.34 1.215 12.615 1.27 ;
 RECT 12.34 1.425 12.44 2.425 ;
 RECT 12.34 1.37 12.615 1.425 ;
 RECT 15.265 0.145 15.365 0.945 ;
 RECT 15.265 1.045 15.365 1.76 ;
 RECT 12.815 1.045 12.915 1.27 ;
 RECT 12.815 1.37 12.915 2.425 ;
 RECT 12.34 1.27 12.915 1.37 ;
 RECT 17.455 1.145 17.555 2.09 ;
 RECT 16.42 1.86 16.52 2.09 ;
 RECT 16.29 1.545 16.52 1.76 ;
 RECT 13.8 0.84 14.03 0.945 ;
 RECT 13.8 1.045 14.03 1.07 ;
 RECT 12.815 0.385 12.915 0.945 ;
 RECT 12.815 0.945 15.365 1.045 ;
 RECT 16.42 2.09 17.555 2.19 ;
 RECT 15.265 1.76 16.52 1.86 ;
 RECT 4.785 0.37 4.885 1.21 ;
 RECT 4.785 1.21 5.07 1.42 ;
 RECT 4.785 1.42 4.885 2.16 ;
 RECT 11.2 0.385 11.3 2.405 ;
 RECT 11.1 2.405 11.33 2.635 ;
 RECT 18.535 0.27 18.635 0.745 ;
 RECT 18.535 0.975 18.635 1.855 ;
 RECT 18.39 0.745 18.635 0.975 ;
 RECT 2.06 0.38 2.16 0.89 ;
 RECT 2.06 1.12 2.16 2.36 ;
 RECT 1.94 0.89 2.17 1.12 ;
 RECT 6.79 0.33 6.89 1.175 ;
 RECT 6.79 1.395 6.89 2.235 ;
 RECT 6.53 1.175 6.89 1.395 ;
 RECT 6.25 0.33 6.35 2.135 ;
 RECT 6.13 2.135 6.36 2.365 ;
 RECT 4.18 1.445 4.28 2.285 ;
 RECT 4.095 2.285 4.325 2.515 ;
 RECT 2.585 1.34 2.815 1.45 ;
 RECT 2.585 0.38 2.685 1.24 ;
 RECT 2.585 1.45 2.685 2.345 ;
 RECT 3.68 0.38 3.78 1.24 ;
 RECT 3.68 1.34 3.78 2.67 ;
 RECT 2.585 1.24 3.78 1.34 ;
 RECT 2.89 0.84 3.135 0.87 ;
 RECT 2.89 0.97 3.135 1.06 ;
 RECT 2.89 0.38 2.99 0.84 ;
 RECT 3.365 0.38 3.465 0.87 ;
 RECT 2.89 0.87 3.465 0.97 ;
 RECT 9.555 1.04 9.655 1.22 ;
 RECT 7.79 1.22 9.655 1.32 ;
 RECT 9.555 1.32 9.655 2.75 ;
 RECT 7.985 0.365 8.085 1.16 ;
 RECT 7.79 1.16 8.085 1.22 ;
 RECT 7.985 1.39 8.085 2.47 ;
 RECT 7.79 1.32 8.085 1.39 ;
 RECT 9.08 0.1 9.18 0.94 ;
 RECT 9.555 0.105 9.655 0.94 ;
 RECT 9.08 0.94 9.655 1.04 ;
 RECT 9.08 1.32 9.18 2.765 ;
 RECT 3.355 1.75 3.455 2.67 ;
 RECT 2.885 1.73 2.985 2.34 ;
 RECT 3.225 1.53 3.455 1.63 ;
 RECT 3.225 1.73 3.455 1.75 ;
 RECT 2.885 1.63 3.455 1.73 ;
 RECT 1.2 0.38 1.3 1.23 ;
 RECT 1.2 1.46 1.3 2.34 ;
 RECT 1.2 1.23 1.435 1.46 ;
 RECT 17.93 0.275 18.03 1.025 ;
 RECT 17.93 1.255 18.03 1.86 ;
 RECT 17.93 1.025 18.21 1.255 ;
 RECT 15.845 0.965 15.945 1.145 ;
 RECT 17.455 0.275 17.555 0.865 ;
 RECT 17.175 0.965 17.275 1.145 ;
 RECT 15.845 1.145 17.275 1.245 ;
 RECT 16.985 1.245 17.085 1.86 ;
 RECT 15.845 0.735 16.075 0.965 ;
 RECT 17.175 0.865 17.555 0.965 ;
 RECT 11.51 1.835 11.61 2.425 ;
 RECT 11.5 1.605 11.73 1.835 ;
 RECT 1.75 1.76 1.85 2.34 ;
 RECT 1.63 1.53 1.86 1.76 ;
 RECT 5.335 0.37 5.435 2.68 ;
 RECT 7.205 2.475 7.435 2.68 ;
 RECT 5.335 2.68 7.435 2.78 ;
 RECT 1.66 0.1 4.355 0.2 ;
 RECT 4.255 0.42 4.355 0.95 ;
 RECT 4.055 0.2 4.355 0.42 ;
 RECT 1.66 0.2 1.76 0.97 ;
 RECT 9.98 0.99 10.235 1.085 ;
 RECT 10.135 1.085 10.235 1.24 ;
 RECT 10.135 0.105 10.235 0.87 ;
 RECT 9.98 0.87 10.235 0.89 ;
 RECT 10.615 0.1 13.465 0.2 ;
 RECT 10.615 0.2 10.715 0.89 ;
 RECT 11.995 0.2 12.095 0.925 ;
 RECT 10.135 1.34 10.235 2.755 ;
 RECT 10.605 1.34 10.705 2.765 ;
 RECT 9.98 0.89 10.715 0.99 ;
 RECT 13.235 0.2 13.465 0.4 ;
 RECT 10.135 1.24 10.705 1.34 ;
 RECT 11.87 0.925 12.1 1.135 ;
 RECT 16.27 0.865 16.995 0.965 ;
 RECT 16.27 0.735 16.5 0.865 ;
 RECT 16.895 0.275 16.995 0.865 ;
 RECT 12.04 2.605 13.39 2.695 ;
 RECT 13.16 2.475 13.39 2.605 ;
 RECT 12.04 1.425 12.14 2.605 ;
 RECT 12.045 2.695 13.39 2.705 ;
 LAYER CO ;
 RECT 18.285 0.47 18.415 0.6 ;
 RECT 18.24 1.455 18.37 1.585 ;
 RECT 10.355 1.675 10.485 1.805 ;
 RECT 9.875 0.395 10.005 0.525 ;
 RECT 9.305 0.585 9.435 0.715 ;
 RECT 9.875 2.34 10.005 2.47 ;
 RECT 10.84 0.395 10.97 0.525 ;
 RECT 10.835 2.34 10.965 2.47 ;
 RECT 8.745 0.395 8.875 0.525 ;
 RECT 6.18 2.185 6.31 2.315 ;
 RECT 16.34 1.595 16.47 1.725 ;
 RECT 19.185 1.44 19.315 1.57 ;
 RECT 0.54 0.36 0.67 0.49 ;
 RECT 0.54 1.71 0.67 1.84 ;
 RECT 0.54 1.97 0.67 2.1 ;
 RECT 0.54 2.23 0.67 2.36 ;
 RECT 12.435 1.255 12.565 1.385 ;
 RECT 7.84 1.21 7.97 1.34 ;
 RECT 7.7 0.605 7.83 0.735 ;
 RECT 8.26 2.025 8.39 2.155 ;
 RECT 8.26 0.605 8.39 0.735 ;
 RECT 6.58 1.215 6.71 1.345 ;
 RECT 4.145 2.335 4.275 2.465 ;
 RECT 3.275 1.57 3.405 1.7 ;
 RECT 2.945 0.89 3.075 1.02 ;
 RECT 1.68 1.58 1.81 1.71 ;
 RECT 1.99 0.94 2.12 1.07 ;
 RECT 7.14 0.57 7.27 0.7 ;
 RECT 7.14 1.87 7.27 2 ;
 RECT 6.515 0.57 6.645 0.7 ;
 RECT 5.045 2.63 5.175 2.76 ;
 RECT 0.94 1.935 1.07 2.065 ;
 RECT 0.94 0.6 1.07 0.73 ;
 RECT 3.085 2.515 3.215 2.645 ;
 RECT 2.315 1.52 2.445 1.65 ;
 RECT 5.62 1.705 5.75 1.835 ;
 RECT 5.62 0.6 5.75 0.73 ;
 RECT 2.315 0.6 2.445 0.73 ;
 RECT 13.285 0.225 13.415 0.355 ;
 RECT 11.92 0.965 12.05 1.095 ;
 RECT 4.89 1.25 5.02 1.38 ;
 RECT 17.68 1.435 17.81 1.565 ;
 RECT 17.68 0.505 17.81 0.635 ;
 RECT 17.205 1.415 17.335 1.545 ;
 RECT 17.205 0.505 17.335 0.635 ;
 RECT 16.645 1.415 16.775 1.545 ;
 RECT 16.645 0.505 16.775 0.635 ;
 RECT 10.355 0.555 10.485 0.685 ;
 RECT 7.7 2.01 7.83 2.14 ;
 RECT 11.745 2.05 11.875 2.18 ;
 RECT 11.745 0.615 11.875 0.745 ;
 RECT 13.04 2.065 13.17 2.195 ;
 RECT 9.305 1.675 9.435 1.805 ;
 RECT 7.255 2.525 7.385 2.655 ;
 RECT 10.03 0.915 10.16 1.045 ;
 RECT 4.105 0.24 4.235 0.37 ;
 RECT 8.825 2.34 8.955 2.47 ;
 RECT 2.635 1.28 2.765 1.41 ;
 RECT 13.85 0.89 13.98 1.02 ;
 RECT 1.255 1.28 1.385 1.41 ;
 RECT 15.895 0.785 16.025 0.915 ;
 RECT 1.41 0.12 1.54 0.25 ;
 RECT 6 0.57 6.13 0.7 ;
 RECT 6 1.48 6.13 1.61 ;
 RECT 6.525 2.375 6.655 2.505 ;
 RECT 0.54 0.62 0.67 0.75 ;
 RECT 3.925 1.67 4.055 1.8 ;
 RECT 1.41 2.515 1.54 2.645 ;
 RECT 15.565 0.225 15.695 0.355 ;
 RECT 5.06 0.6 5.19 0.73 ;
 RECT 4.485 0.6 4.615 0.73 ;
 RECT 4.485 1.48 4.615 1.61 ;
 RECT 3.925 0.6 4.055 0.73 ;
 RECT 3.115 0.555 3.245 0.685 ;
 RECT 15.565 1.475 15.695 1.605 ;
 RECT 14.96 1.255 15.09 1.385 ;
 RECT 14.915 0.505 15.045 0.635 ;
 RECT 13.21 2.525 13.34 2.655 ;
 RECT 11.15 2.455 11.28 2.585 ;
 RECT 11.55 1.655 11.68 1.785 ;
 RECT 13.04 0.615 13.17 0.745 ;
 RECT 12.56 0.615 12.69 0.745 ;
 RECT 12.56 2.075 12.69 2.205 ;
 RECT 16.32 0.785 16.45 0.915 ;
 RECT 18.44 0.795 18.57 0.925 ;
 RECT 18.03 1.075 18.16 1.205 ;
 RECT 18.765 0.505 18.895 0.635 ;
 RECT 18.765 1.44 18.895 1.57 ;
 LAYER M1 ;
 RECT 12.34 1.17 12.68 1.51 ;
 RECT 1.25 1.21 1.39 1.275 ;
 RECT 1.25 1.415 1.39 1.48 ;
 RECT 2.31 0.55 2.45 1.275 ;
 RECT 2.31 1.415 2.45 1.71 ;
 RECT 1.25 1.275 2.45 1.415 ;
 RECT 4.48 0.55 4.62 1.475 ;
 RECT 4.415 1.475 4.685 1.615 ;
 RECT 14.955 0.64 15.095 0.78 ;
 RECT 14.955 0.92 15.095 1.455 ;
 RECT 14.85 0.5 15.095 0.64 ;
 RECT 14.955 0.78 16.09 0.92 ;
 RECT 12.18 1.845 12.32 2.45 ;
 RECT 11.145 2.385 11.285 2.45 ;
 RECT 11.145 2.45 12.32 2.59 ;
 RECT 11.145 2.59 11.285 2.65 ;
 RECT 13.035 0.55 13.175 1.705 ;
 RECT 12.18 1.705 13.175 1.845 ;
 RECT 13.035 1.845 13.175 2.265 ;
 RECT 18.76 0.435 18.9 1.07 ;
 RECT 18.76 1.21 18.9 1.64 ;
 RECT 17.96 1.07 18.9 1.21 ;
 RECT 16.335 0.92 16.475 1.785 ;
 RECT 16.25 0.78 16.5 0.92 ;
 RECT 9.02 0.385 9.16 0.87 ;
 RECT 8.255 0.87 9.16 1.01 ;
 RECT 8.255 0.55 8.395 0.87 ;
 RECT 8.255 1.01 8.395 2.21 ;
 RECT 9.58 0.385 9.72 0.75 ;
 RECT 9.02 0.245 9.72 0.385 ;
 RECT 10.025 0.89 10.165 1.095 ;
 RECT 9.58 0.75 10.165 0.89 ;
 RECT 11.545 1.095 11.685 1.835 ;
 RECT 11.87 0.925 12.1 0.955 ;
 RECT 11.87 1.095 12.1 1.135 ;
 RECT 11.545 0.955 12.1 1.095 ;
 RECT 15.235 0.36 15.375 0.5 ;
 RECT 13.185 0.22 15.375 0.36 ;
 RECT 16.64 0.435 16.78 0.5 ;
 RECT 16.64 0.64 16.78 1.61 ;
 RECT 15.235 0.5 16.78 0.64 ;
 RECT 17.2 0.36 17.34 1.41 ;
 RECT 18 0.36 18.14 0.79 ;
 RECT 17.135 1.41 17.405 1.55 ;
 RECT 17.2 0.22 18.14 0.36 ;
 RECT 18 0.79 18.62 0.93 ;
 RECT 15.235 1.33 15.375 2.52 ;
 RECT 13.13 2.52 15.375 2.66 ;
 RECT 17.675 0.64 17.815 1.925 ;
 RECT 15.885 1.33 16.025 1.925 ;
 RECT 17.61 0.5 17.86 0.64 ;
 RECT 15.885 1.925 17.815 2.065 ;
 RECT 15.235 1.19 16.025 1.33 ;
 RECT 0.935 0.6 1.075 2.13 ;
 RECT 1.87 0.41 2.01 0.46 ;
 RECT 2.63 0.41 2.77 1.475 ;
 RECT 1.87 0.27 2.77 0.41 ;
 RECT 0.935 0.46 2.01 0.6 ;
 RECT 7.415 1.775 7.555 2.52 ;
 RECT 7.185 2.52 7.555 2.66 ;
 RECT 8.535 2.135 8.675 2.435 ;
 RECT 7.975 1.775 8.115 2.435 ;
 RECT 7.415 1.635 8.115 1.775 ;
 RECT 7.975 2.435 8.675 2.575 ;
 RECT 10.76 1.86 10.9 1.995 ;
 RECT 11.26 2.045 11.925 2.185 ;
 RECT 11.26 1.86 11.4 2.045 ;
 RECT 11.26 0.75 11.4 1.72 ;
 RECT 10.76 1.72 11.4 1.86 ;
 RECT 8.535 1.995 10.9 2.135 ;
 RECT 11.26 0.61 11.97 0.75 ;
 RECT 3.44 0.375 3.58 1.26 ;
 RECT 4.77 0.375 4.91 0.93 ;
 RECT 3.27 1.26 3.58 1.4 ;
 RECT 3.27 1.4 3.41 1.77 ;
 RECT 3.44 0.235 4.91 0.375 ;
 RECT 5.335 0.24 6.135 0.38 ;
 RECT 5.995 0.38 6.135 1.66 ;
 RECT 5.335 0.38 5.475 0.93 ;
 RECT 4.77 0.93 5.475 1.07 ;
 RECT 6.175 2.23 6.315 2.33 ;
 RECT 3.805 2.33 6.315 2.47 ;
 RECT 3.805 2.085 3.945 2.33 ;
 RECT 1.675 1.945 3.945 2.085 ;
 RECT 2.94 0.835 3.08 1.945 ;
 RECT 1.675 1.715 1.815 1.945 ;
 RECT 1.605 1.575 1.88 1.715 ;
 RECT 6.175 2.09 7.275 2.23 ;
 RECT 7.135 0.52 7.275 2.09 ;
 RECT 5.895 1.94 6.035 2.05 ;
 RECT 4.135 2.05 6.035 2.19 ;
 RECT 4.135 1.805 4.275 2.05 ;
 RECT 3.92 0.545 4.06 1.665 ;
 RECT 3.855 1.665 4.275 1.805 ;
 RECT 6.855 0.365 6.995 1.8 ;
 RECT 7.415 0.365 7.555 1.205 ;
 RECT 6.855 0.225 7.555 0.365 ;
 RECT 5.895 1.8 6.995 1.94 ;
 RECT 7.415 1.205 8.04 1.345 ;
 RECT 5.615 0.55 5.755 1.245 ;
 RECT 5.615 1.385 5.755 1.9 ;
 RECT 4.84 1.245 5.755 1.385 ;
 RECT 4.84 1.21 5.07 1.245 ;
 RECT 4.84 1.385 5.07 1.42 ;
 END
END RDFFNX2

MACRO RDFFX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 20.16 BY 2.88 ;
 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.31 0.835 6.72 1.12 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.645 1.5 8.785 2.295 ;
 RECT 8.645 1.09 9.065 1.5 ;
 RECT 8.645 0.525 8.785 1.09 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.695 1.12 10.07 1.465 ;
 RECT 9.695 1.465 9.835 1.79 ;
 RECT 9.695 0.48 9.835 1.12 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 20.16 2.96 ;
 RECT 4.995 2.615 5.23 2.8 ;
 RECT 3.04 2.51 3.27 2.65 ;
 RECT 1.345 2.51 1.615 2.65 ;
 RECT 6.505 2.37 6.775 2.51 ;
 RECT 9.215 2.275 9.355 2.8 ;
 RECT 7.7 1.94 7.84 2.8 ;
 RECT 10.255 2 10.395 2.8 ;
 RECT 0.485 1.64 0.645 2.8 ;
 RECT 11.945 2.025 12.085 2.8 ;
 RECT 3.085 2.65 3.225 2.8 ;
 RECT 1.41 2.65 1.55 2.8 ;
 RECT 6.57 2.51 6.71 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 20.16 0.08 ;
 RECT 6.45 0.555 6.72 0.695 ;
 RECT 14.905 0.22 15.155 0.36 ;
 RECT 3.05 0.555 3.3 0.695 ;
 RECT 9.215 0.08 9.355 0.575 ;
 RECT 7.7 0.08 7.84 0.785 ;
 RECT 1.41 0.08 1.55 0.32 ;
 RECT 5.06 0.08 5.2 0.78 ;
 RECT 10.305 0.08 10.445 0.865 ;
 RECT 11.945 0.08 12.085 0.815 ;
 RECT 0.485 0.08 0.645 0.84 ;
 RECT 17.67 0.08 17.81 0.65 ;
 RECT 6.515 0.08 6.655 0.555 ;
 RECT 14.95 0.08 15.09 0.22 ;
 RECT 3.115 0.08 3.255 0.555 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 18.525 1.4 18.865 1.765 ;
 RECT 14.94 2.225 18.69 2.385 ;
 RECT 14.905 1.47 15.135 1.61 ;
 RECT 17.625 1.395 17.765 2.225 ;
 RECT 18.54 1.765 18.68 2.225 ;
 RECT 14.95 1.61 15.09 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.075 0.81 13.455 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.78 0.83 2.175 1.135 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 14.655 1.76 15.91 1.86 ;
 RECT 7.99 0.365 8.09 1.16 ;
 RECT 7.795 1.16 8.09 1.22 ;
 RECT 7.99 1.39 8.09 2.47 ;
 RECT 7.795 1.32 8.09 1.39 ;
 RECT 8.9 0.105 9 1.22 ;
 RECT 8.9 1.32 9 2.75 ;
 RECT 7.795 1.22 9 1.32 ;
 RECT 6.835 0.33 6.935 1.27 ;
 RECT 6.835 1.49 6.935 2.235 ;
 RECT 6.535 1.27 6.935 1.49 ;
 RECT 11.385 0.205 11.485 0.925 ;
 RECT 9.48 0.105 12.855 0.205 ;
 RECT 12.625 0.205 12.855 0.4 ;
 RECT 9.48 0.205 9.58 0.87 ;
 RECT 9.335 0.87 9.58 1.085 ;
 RECT 9.48 1.085 9.58 2.755 ;
 RECT 11.26 0.925 11.49 1.135 ;
 RECT 10.59 0.385 10.69 2.405 ;
 RECT 10.49 2.405 10.72 2.635 ;
 RECT 17.925 0.27 18.025 0.745 ;
 RECT 17.925 0.975 18.025 1.855 ;
 RECT 17.78 0.745 18.025 0.975 ;
 RECT 10.9 1.835 11 2.425 ;
 RECT 10.89 1.605 11.12 1.835 ;
 RECT 2.065 0.38 2.165 0.93 ;
 RECT 2.065 1.16 2.165 2.36 ;
 RECT 1.945 0.93 2.175 1.16 ;
 RECT 1.755 1.76 1.855 2.34 ;
 RECT 1.635 1.53 1.865 1.76 ;
 RECT 6.255 0.33 6.355 0.865 ;
 RECT 6.255 1.08 6.355 2.235 ;
 RECT 6.255 0.865 6.545 1.08 ;
 RECT 1.17 0.38 1.27 1.23 ;
 RECT 1.17 1.46 1.27 2.34 ;
 RECT 1.17 1.23 1.4 1.46 ;
 RECT 4.185 1.445 4.285 2.285 ;
 RECT 4.1 2.285 4.33 2.515 ;
 RECT 2.59 1.34 2.82 1.45 ;
 RECT 2.59 0.38 2.69 1.24 ;
 RECT 2.59 1.45 2.69 2.345 ;
 RECT 3.685 0.38 3.785 1.24 ;
 RECT 3.685 1.34 3.785 2.435 ;
 RECT 2.59 1.24 3.785 1.34 ;
 RECT 3.36 1.75 3.46 2.44 ;
 RECT 3.23 1.53 3.46 1.63 ;
 RECT 3.23 1.73 3.46 1.75 ;
 RECT 2.89 1.73 2.99 2.34 ;
 RECT 2.89 1.63 3.46 1.73 ;
 RECT 2.895 0.84 3.14 0.87 ;
 RECT 2.895 0.97 3.14 1.06 ;
 RECT 2.895 0.38 2.995 0.84 ;
 RECT 3.37 0.38 3.47 0.87 ;
 RECT 2.895 0.87 3.47 0.97 ;
 RECT 1.665 0.1 4.36 0.2 ;
 RECT 4.06 0.2 4.36 0.42 ;
 RECT 1.665 0.2 1.765 0.97 ;
 RECT 4.26 0.42 4.36 0.95 ;
 RECT 4.79 0.37 4.89 1.21 ;
 RECT 4.79 1.21 5.075 1.42 ;
 RECT 4.79 1.42 4.89 2.16 ;
 RECT 11.43 2.605 12.78 2.695 ;
 RECT 11.43 1.425 11.53 2.605 ;
 RECT 11.435 2.695 12.78 2.705 ;
 RECT 10.895 0.385 10.995 1.325 ;
 RECT 12.55 2.475 12.78 2.605 ;
 RECT 10.895 1.325 11.53 1.425 ;
 RECT 17.32 0.275 17.42 1.025 ;
 RECT 17.32 1.255 17.42 1.86 ;
 RECT 17.32 1.025 17.6 1.255 ;
 RECT 5.34 0.37 5.44 2.68 ;
 RECT 7.21 2.475 7.44 2.68 ;
 RECT 5.34 2.68 7.44 2.78 ;
 RECT 15.235 0.965 15.335 1.145 ;
 RECT 16.845 0.275 16.945 0.865 ;
 RECT 16.565 0.965 16.665 1.145 ;
 RECT 15.235 1.145 16.665 1.245 ;
 RECT 16.375 1.245 16.475 1.86 ;
 RECT 15.235 0.735 15.465 0.965 ;
 RECT 16.565 0.865 16.945 0.965 ;
 RECT 15.66 0.865 16.385 0.965 ;
 RECT 15.66 0.735 15.89 0.865 ;
 RECT 16.285 0.275 16.385 0.865 ;
 RECT 11.73 1.215 12.005 1.27 ;
 RECT 11.73 1.37 12.005 1.425 ;
 RECT 11.73 1.27 12.305 1.37 ;
 RECT 12.205 1.045 12.305 1.27 ;
 RECT 12.205 1.37 12.305 2.425 ;
 RECT 14.655 1.045 14.755 1.76 ;
 RECT 16.845 1.145 16.945 2.09 ;
 RECT 15.81 1.86 15.91 2.09 ;
 RECT 11.73 0.385 11.83 1.215 ;
 RECT 11.73 1.425 11.83 2.425 ;
 RECT 15.68 1.545 15.91 1.76 ;
 RECT 13.165 0.84 13.395 0.945 ;
 RECT 13.165 1.045 13.395 1.07 ;
 RECT 12.205 0.385 12.305 0.945 ;
 RECT 12.205 0.945 14.755 1.045 ;
 RECT 14.655 0.145 14.755 0.945 ;
 RECT 15.81 2.09 16.945 2.19 ;
 LAYER CO ;
 RECT 0.9 0.6 1.03 0.73 ;
 RECT 3.93 1.67 4.06 1.8 ;
 RECT 1.415 2.515 1.545 2.645 ;
 RECT 3.09 2.515 3.22 2.645 ;
 RECT 2.32 1.52 2.45 1.65 ;
 RECT 5.625 1.705 5.755 1.835 ;
 RECT 5.625 0.6 5.755 0.73 ;
 RECT 5.065 0.6 5.195 0.73 ;
 RECT 4.49 0.6 4.62 0.73 ;
 RECT 4.49 1.48 4.62 1.61 ;
 RECT 3.93 0.6 4.06 0.73 ;
 RECT 3.12 0.555 3.25 0.685 ;
 RECT 2.32 0.6 2.45 0.73 ;
 RECT 12.675 0.225 12.805 0.355 ;
 RECT 14.955 1.475 15.085 1.605 ;
 RECT 14.35 1.255 14.48 1.385 ;
 RECT 14.305 0.505 14.435 0.635 ;
 RECT 12.6 2.525 12.73 2.655 ;
 RECT 10.54 2.455 10.67 2.585 ;
 RECT 10.94 1.655 11.07 1.785 ;
 RECT 12.43 0.635 12.56 0.765 ;
 RECT 15.71 0.785 15.84 0.915 ;
 RECT 17.83 0.795 17.96 0.925 ;
 RECT 17.42 1.075 17.55 1.205 ;
 RECT 18.155 0.505 18.285 0.635 ;
 RECT 18.155 1.44 18.285 1.57 ;
 RECT 17.675 0.47 17.805 0.6 ;
 RECT 17.63 1.455 17.76 1.585 ;
 RECT 17.07 1.435 17.2 1.565 ;
 RECT 17.07 0.505 17.2 0.635 ;
 RECT 7.26 2.525 7.39 2.655 ;
 RECT 9.385 0.915 9.515 1.045 ;
 RECT 9.7 1.6 9.83 1.73 ;
 RECT 9.22 0.395 9.35 0.525 ;
 RECT 8.65 0.585 8.78 0.715 ;
 RECT 8.65 2.105 8.78 2.235 ;
 RECT 9.22 2.34 9.35 2.47 ;
 RECT 11.825 1.255 11.955 1.385 ;
 RECT 11.31 0.965 11.44 1.095 ;
 RECT 6.365 0.91 6.495 1.04 ;
 RECT 6.585 1.31 6.715 1.44 ;
 RECT 4.15 2.335 4.28 2.465 ;
 RECT 4.11 0.24 4.24 0.37 ;
 RECT 3.28 1.57 3.41 1.7 ;
 RECT 4.895 1.25 5.025 1.38 ;
 RECT 13.215 0.89 13.345 1.02 ;
 RECT 15.73 1.595 15.86 1.725 ;
 RECT 15.285 0.785 15.415 0.915 ;
 RECT 1.415 0.12 1.545 0.25 ;
 RECT 18.575 1.44 18.705 1.57 ;
 RECT 0.5 0.36 0.63 0.49 ;
 RECT 0.5 0.62 0.63 0.75 ;
 RECT 0.5 1.71 0.63 1.84 ;
 RECT 0.5 1.97 0.63 2.1 ;
 RECT 0.5 2.23 0.63 2.36 ;
 RECT 14.955 0.225 15.085 0.355 ;
 RECT 16.595 1.415 16.725 1.545 ;
 RECT 16.595 0.505 16.725 0.635 ;
 RECT 16.035 1.415 16.165 1.545 ;
 RECT 16.035 0.505 16.165 0.635 ;
 RECT 9.7 0.555 9.83 0.685 ;
 RECT 7.705 2.01 7.835 2.14 ;
 RECT 7.845 1.21 7.975 1.34 ;
 RECT 7.705 0.605 7.835 0.735 ;
 RECT 8.265 2.025 8.395 2.155 ;
 RECT 8.265 0.605 8.395 0.735 ;
 RECT 11.95 0.635 12.08 0.765 ;
 RECT 11.95 2.075 12.08 2.205 ;
 RECT 11.135 2.05 11.265 2.18 ;
 RECT 11.135 0.635 11.265 0.765 ;
 RECT 10.31 0.635 10.44 0.765 ;
 RECT 10.26 2.06 10.39 2.19 ;
 RECT 12.43 2.065 12.56 2.195 ;
 RECT 8.65 1.715 8.78 1.845 ;
 RECT 2.95 0.89 3.08 1.02 ;
 RECT 2.64 1.28 2.77 1.41 ;
 RECT 1.685 1.58 1.815 1.71 ;
 RECT 1.995 0.98 2.125 1.11 ;
 RECT 1.22 1.28 1.35 1.41 ;
 RECT 7.145 0.57 7.275 0.7 ;
 RECT 7.145 1.64 7.275 1.77 ;
 RECT 6.52 0.56 6.65 0.69 ;
 RECT 6.005 0.57 6.135 0.7 ;
 RECT 6.005 1.48 6.135 1.61 ;
 RECT 6.575 2.375 6.705 2.505 ;
 RECT 5.05 2.63 5.18 2.76 ;
 RECT 0.9 1.935 1.03 2.065 ;
 LAYER M1 ;
 RECT 11.73 1.17 12.07 1.51 ;
 RECT 4.485 0.55 4.625 1.475 ;
 RECT 4.42 1.475 4.69 1.615 ;
 RECT 1.215 1.21 1.355 1.275 ;
 RECT 1.215 1.415 1.355 1.48 ;
 RECT 2.315 0.55 2.455 1.275 ;
 RECT 2.315 1.415 2.455 1.71 ;
 RECT 1.215 1.275 2.455 1.415 ;
 RECT 14.345 0.64 14.485 0.78 ;
 RECT 14.345 0.92 14.485 1.455 ;
 RECT 14.24 0.5 14.485 0.64 ;
 RECT 14.345 0.78 15.48 0.92 ;
 RECT 15.725 0.92 15.865 1.785 ;
 RECT 15.64 0.78 15.89 0.92 ;
 RECT 14.625 0.36 14.765 0.5 ;
 RECT 12.575 0.22 14.765 0.36 ;
 RECT 16.03 0.435 16.17 0.5 ;
 RECT 16.03 0.64 16.17 1.61 ;
 RECT 14.625 0.5 16.17 0.64 ;
 RECT 5.9 1.94 6.04 2.05 ;
 RECT 4.14 2.05 6.04 2.19 ;
 RECT 4.14 1.805 4.28 2.05 ;
 RECT 3.855 1.665 4.28 1.805 ;
 RECT 3.925 0.545 4.065 1.665 ;
 RECT 7.42 0.365 7.56 1.205 ;
 RECT 6.86 0.365 7 1.8 ;
 RECT 6.86 0.225 7.56 0.365 ;
 RECT 5.9 1.8 7 1.94 ;
 RECT 7.42 1.205 8.045 1.345 ;
 RECT 11.26 0.925 11.49 0.955 ;
 RECT 10.935 0.955 11.49 1.095 ;
 RECT 11.26 1.095 11.49 1.135 ;
 RECT 10.935 1.095 11.075 1.835 ;
 RECT 0.895 0.6 1.035 2.13 ;
 RECT 1.875 0.41 2.015 0.46 ;
 RECT 0.895 0.46 2.015 0.6 ;
 RECT 1.875 0.275 2.775 0.41 ;
 RECT 2.635 0.41 2.775 1.475 ;
 RECT 1.875 0.27 2.71 0.275 ;
 RECT 1.875 0.6 2.015 0.61 ;
 RECT 8.26 0.24 8.4 0.245 ;
 RECT 8.26 0.385 8.4 2.21 ;
 RECT 8.925 0.385 9.065 0.75 ;
 RECT 8.26 0.245 9.065 0.385 ;
 RECT 9.38 0.89 9.52 1.095 ;
 RECT 8.925 0.75 9.52 0.89 ;
 RECT 5.34 0.24 6.14 0.38 ;
 RECT 6 0.38 6.14 1.305 ;
 RECT 5.34 0.38 5.48 0.93 ;
 RECT 6 1.445 6.14 1.66 ;
 RECT 4.775 0.93 5.48 1.07 ;
 RECT 3.445 0.375 3.585 1.26 ;
 RECT 4.775 0.375 4.915 0.93 ;
 RECT 3.275 1.26 3.585 1.4 ;
 RECT 3.275 1.4 3.415 1.77 ;
 RECT 3.445 0.235 4.915 0.375 ;
 RECT 6.58 1.26 6.72 1.305 ;
 RECT 6.58 1.445 6.72 1.495 ;
 RECT 6 1.305 6.72 1.445 ;
 RECT 17.39 0.36 17.53 0.79 ;
 RECT 16.59 0.36 16.73 1.41 ;
 RECT 16.525 1.41 16.795 1.55 ;
 RECT 16.59 0.22 17.53 0.36 ;
 RECT 17.39 0.79 18.01 0.93 ;
 RECT 11.57 1.845 11.71 2.45 ;
 RECT 10.535 2.385 10.675 2.45 ;
 RECT 10.535 2.45 11.71 2.59 ;
 RECT 10.535 2.59 10.675 2.65 ;
 RECT 12.425 0.585 12.565 1.705 ;
 RECT 11.57 1.705 12.565 1.845 ;
 RECT 12.425 1.845 12.565 2.265 ;
 RECT 12.52 2.52 14.765 2.65 ;
 RECT 12.52 2.65 14.755 2.66 ;
 RECT 14.625 1.33 14.765 2.52 ;
 RECT 17.065 0.64 17.205 1.925 ;
 RECT 15.275 1.33 15.415 1.925 ;
 RECT 17 0.5 17.25 0.64 ;
 RECT 15.275 1.925 17.205 2.065 ;
 RECT 14.625 1.19 15.415 1.33 ;
 RECT 18.15 0.435 18.29 1.07 ;
 RECT 17.35 1.07 18.29 1.21 ;
 RECT 18.15 1.21 18.29 1.64 ;
 RECT 3.81 2.085 3.95 2.33 ;
 RECT 1.675 1.945 3.95 2.085 ;
 RECT 2.945 0.835 3.085 1.945 ;
 RECT 1.68 1.715 1.82 1.945 ;
 RECT 1.61 1.575 1.885 1.715 ;
 RECT 3.81 2.33 6.32 2.47 ;
 RECT 6.18 2.23 6.32 2.33 ;
 RECT 7.14 0.52 7.28 2.09 ;
 RECT 6.18 2.09 7.28 2.23 ;
 RECT 7.98 1.775 8.12 2.435 ;
 RECT 7.42 1.635 8.12 1.775 ;
 RECT 7.42 1.775 7.56 2.52 ;
 RECT 7.19 2.52 7.56 2.66 ;
 RECT 9.975 1.86 10.115 1.995 ;
 RECT 8.935 1.995 10.115 2.135 ;
 RECT 8.935 2.135 9.075 2.435 ;
 RECT 7.98 2.435 9.075 2.575 ;
 RECT 10.65 2.045 11.315 2.185 ;
 RECT 10.65 1.86 10.79 2.045 ;
 RECT 10.65 0.63 11.315 0.77 ;
 RECT 10.65 0.77 10.79 1.72 ;
 RECT 9.975 1.72 10.79 1.86 ;
 RECT 5.62 0.55 5.76 1.245 ;
 RECT 5.62 1.385 5.76 1.9 ;
 RECT 4.845 1.245 5.76 1.385 ;
 RECT 4.845 1.21 5.075 1.245 ;
 RECT 4.845 1.385 5.075 1.42 ;
 END
END RDFFX1

MACRO RDFFX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 20.48 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.985 1.09 9.405 1.5 ;
 RECT 8.985 1.5 9.125 1.855 ;
 RECT 8.985 0.525 9.125 1.09 ;
 END
 ANTENNADIFFAREA 0.584 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.96 1.12 10.24 1.465 ;
 RECT 10.035 1.465 10.175 1.855 ;
 RECT 10.035 0.48 10.175 1.12 ;
 END
 ANTENNADIFFAREA 0.6 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 20.48 2.96 ;
 RECT 9.51 2.275 9.65 2.8 ;
 RECT 4.675 2.615 4.91 2.8 ;
 RECT 6.14 2.37 6.41 2.51 ;
 RECT 2.72 2.51 2.95 2.65 ;
 RECT 1.025 2.51 1.295 2.65 ;
 RECT 7.38 1.94 7.52 2.8 ;
 RECT 12.27 2.025 12.41 2.8 ;
 RECT 10.515 2.275 10.655 2.8 ;
 RECT 0.185 1.64 0.345 2.8 ;
 RECT 8.505 2.275 8.645 2.8 ;
 RECT 6.205 2.51 6.345 2.8 ;
 RECT 2.765 2.65 2.905 2.8 ;
 RECT 1.09 2.65 1.23 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 20.48 0.08 ;
 RECT 9.555 0.08 9.695 0.575 ;
 RECT 6.13 0.56 6.4 0.7 ;
 RECT 2.73 0.555 2.98 0.695 ;
 RECT 15.23 0.22 15.48 0.36 ;
 RECT 0.185 0.08 0.345 0.84 ;
 RECT 12.27 0.08 12.41 0.815 ;
 RECT 8.425 0.08 8.565 0.575 ;
 RECT 10.51 0.08 10.65 0.575 ;
 RECT 7.38 0.08 7.52 0.785 ;
 RECT 17.995 0.08 18.135 0.65 ;
 RECT 4.74 0.08 4.88 0.78 ;
 RECT 1.09 0.08 1.23 0.32 ;
 RECT 6.195 0.08 6.335 0.56 ;
 RECT 2.795 0.08 2.935 0.555 ;
 RECT 15.275 0.08 15.415 0.22 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 18.85 1.4 19.19 1.765 ;
 RECT 15.265 2.225 19.015 2.385 ;
 RECT 15.23 1.47 15.46 1.61 ;
 RECT 17.95 1.395 18.09 2.225 ;
 RECT 18.865 1.765 19.005 2.225 ;
 RECT 15.275 1.61 15.415 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.4 0.81 13.78 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.02 0.84 6.385 1.115 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 0.84 1.855 1.135 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 9.635 0.87 9.92 0.88 ;
 RECT 11.71 0.205 11.81 0.925 ;
 RECT 10.29 0.205 10.39 0.88 ;
 RECT 9.635 0.88 10.39 0.98 ;
 RECT 9.82 1.23 10.39 1.33 ;
 RECT 9.82 1.33 9.92 2.755 ;
 RECT 10.29 1.33 10.39 2.77 ;
 RECT 12.95 0.205 13.18 0.4 ;
 RECT 10.29 0.105 13.18 0.205 ;
 RECT 11.585 0.925 11.815 1.135 ;
 RECT 5.02 0.37 5.12 2.68 ;
 RECT 6.89 2.475 7.12 2.68 ;
 RECT 5.02 2.68 7.12 2.78 ;
 RECT 2.575 0.87 3.15 0.97 ;
 RECT 3.05 0.38 3.15 0.87 ;
 RECT 2.575 0.84 2.82 0.87 ;
 RECT 2.575 0.97 2.82 1.06 ;
 RECT 2.575 0.38 2.675 0.84 ;
 RECT 10.915 0.385 11.015 2.405 ;
 RECT 10.815 2.405 11.045 2.635 ;
 RECT 1.745 0.38 1.845 0.945 ;
 RECT 1.745 1.175 1.845 2.36 ;
 RECT 1.625 0.945 1.855 1.175 ;
 RECT 0.85 0.38 0.95 1.23 ;
 RECT 0.85 1.46 0.95 2.34 ;
 RECT 0.85 1.23 1.08 1.46 ;
 RECT 4.47 0.37 4.57 1.21 ;
 RECT 4.47 1.21 4.755 1.42 ;
 RECT 4.47 1.42 4.57 2.16 ;
 RECT 17.645 0.275 17.745 1.025 ;
 RECT 17.645 1.255 17.745 1.86 ;
 RECT 17.645 1.025 17.925 1.255 ;
 RECT 11.225 1.835 11.325 2.425 ;
 RECT 11.215 1.605 11.445 1.835 ;
 RECT 1.345 0.1 4.04 0.2 ;
 RECT 3.74 0.2 4.04 0.42 ;
 RECT 1.345 0.2 1.445 0.97 ;
 RECT 3.94 0.42 4.04 0.95 ;
 RECT 1.435 1.76 1.535 2.34 ;
 RECT 1.315 1.53 1.545 1.76 ;
 RECT 6.475 0.33 6.575 1.27 ;
 RECT 6.475 1.49 6.575 2.235 ;
 RECT 6.215 1.27 6.575 1.49 ;
 RECT 3.865 1.445 3.965 2.285 ;
 RECT 3.78 2.285 4.01 2.515 ;
 RECT 7.67 0.365 7.77 1.16 ;
 RECT 7.475 1.16 7.77 1.22 ;
 RECT 7.67 1.39 7.77 2.47 ;
 RECT 7.475 1.32 7.77 1.39 ;
 RECT 9.24 0.98 9.34 1.22 ;
 RECT 9.24 1.32 9.34 2.75 ;
 RECT 7.475 1.22 9.34 1.32 ;
 RECT 8.77 1.32 8.87 2.77 ;
 RECT 9.24 0.105 9.34 0.88 ;
 RECT 8.77 0.095 8.87 0.88 ;
 RECT 8.77 0.88 9.34 0.98 ;
 RECT 3.04 1.75 3.14 2.47 ;
 RECT 2.91 1.53 3.14 1.63 ;
 RECT 2.91 1.73 3.14 1.75 ;
 RECT 2.57 1.73 2.67 2.34 ;
 RECT 2.57 1.63 3.14 1.73 ;
 RECT 17.17 0.275 17.27 0.865 ;
 RECT 16.89 0.965 16.99 1.145 ;
 RECT 15.56 0.965 15.66 1.145 ;
 RECT 15.56 1.145 16.99 1.245 ;
 RECT 16.7 1.245 16.8 1.86 ;
 RECT 16.89 0.865 17.27 0.965 ;
 RECT 15.56 0.735 15.79 0.965 ;
 RECT 18.25 0.27 18.35 0.745 ;
 RECT 18.25 0.975 18.35 1.855 ;
 RECT 18.105 0.745 18.35 0.975 ;
 RECT 5.935 0.33 6.035 0.86 ;
 RECT 5.935 1.09 6.035 2.235 ;
 RECT 5.935 0.86 6.245 1.09 ;
 RECT 15.985 0.865 16.71 0.965 ;
 RECT 15.985 0.735 16.215 0.865 ;
 RECT 16.61 0.275 16.71 0.865 ;
 RECT 2.27 1.34 2.5 1.45 ;
 RECT 2.27 0.38 2.37 1.24 ;
 RECT 2.27 1.45 2.37 2.345 ;
 RECT 3.365 0.38 3.465 1.24 ;
 RECT 2.27 1.24 3.465 1.34 ;
 RECT 3.365 1.34 3.465 2.47 ;
 RECT 12.055 1.27 12.63 1.37 ;
 RECT 14.98 0.145 15.08 0.945 ;
 RECT 14.98 1.045 15.08 1.76 ;
 RECT 12.53 1.045 12.63 1.27 ;
 RECT 12.53 1.37 12.63 2.425 ;
 RECT 12.055 0.385 12.155 1.215 ;
 RECT 12.055 1.215 12.33 1.27 ;
 RECT 17.17 1.145 17.27 2.09 ;
 RECT 16.135 1.86 16.235 2.09 ;
 RECT 16.005 1.545 16.235 1.76 ;
 RECT 13.49 0.84 13.72 0.945 ;
 RECT 13.49 1.045 13.72 1.07 ;
 RECT 12.53 0.385 12.63 0.945 ;
 RECT 12.53 0.945 15.08 1.045 ;
 RECT 12.055 1.425 12.155 2.425 ;
 RECT 12.055 1.37 12.33 1.425 ;
 RECT 16.135 2.09 17.27 2.19 ;
 RECT 14.98 1.76 16.235 1.86 ;
 RECT 11.755 2.605 13.105 2.695 ;
 RECT 12.875 2.475 13.105 2.605 ;
 RECT 11.755 1.425 11.855 2.605 ;
 RECT 11.76 2.695 13.105 2.705 ;
 RECT 11.22 0.385 11.32 1.325 ;
 RECT 11.22 1.325 11.855 1.425 ;
 RECT 9.82 1.085 9.92 1.23 ;
 RECT 9.635 0.98 9.92 1.085 ;
 RECT 9.82 0.105 9.92 0.87 ;
 LAYER CO ;
 RECT 6.265 1.31 6.395 1.44 ;
 RECT 3.83 2.335 3.96 2.465 ;
 RECT 9.685 0.915 9.815 1.045 ;
 RECT 10.04 1.675 10.17 1.805 ;
 RECT 2.96 1.57 3.09 1.7 ;
 RECT 1.365 1.58 1.495 1.71 ;
 RECT 1.675 0.995 1.805 1.125 ;
 RECT 0.9 1.28 1.03 1.41 ;
 RECT 4.73 2.63 4.86 2.76 ;
 RECT 0.6 1.935 0.73 2.065 ;
 RECT 0.6 0.6 0.73 0.73 ;
 RECT 3.61 1.67 3.74 1.8 ;
 RECT 1.095 2.515 1.225 2.645 ;
 RECT 3.61 0.6 3.74 0.73 ;
 RECT 2.8 0.555 2.93 0.685 ;
 RECT 2 0.6 2.13 0.73 ;
 RECT 13 0.225 13.13 0.355 ;
 RECT 10.865 2.455 10.995 2.585 ;
 RECT 11.265 1.655 11.395 1.785 ;
 RECT 12.755 0.615 12.885 0.745 ;
 RECT 12.275 0.615 12.405 0.745 ;
 RECT 12.275 2.075 12.405 2.205 ;
 RECT 17.745 1.075 17.875 1.205 ;
 RECT 18.48 0.505 18.61 0.635 ;
 RECT 18.48 1.44 18.61 1.57 ;
 RECT 18 0.47 18.13 0.6 ;
 RECT 17.955 1.455 18.085 1.585 ;
 RECT 17.395 1.435 17.525 1.565 ;
 RECT 9.56 0.395 9.69 0.525 ;
 RECT 10.515 0.395 10.645 0.525 ;
 RECT 10.52 2.34 10.65 2.47 ;
 RECT 8.43 0.395 8.56 0.525 ;
 RECT 7.945 2.025 8.075 2.155 ;
 RECT 3.79 0.24 3.92 0.37 ;
 RECT 12.15 1.255 12.28 1.385 ;
 RECT 2.63 0.89 2.76 1.02 ;
 RECT 2.32 1.28 2.45 1.41 ;
 RECT 8.51 2.34 8.64 2.47 ;
 RECT 13.54 0.89 13.67 1.02 ;
 RECT 6.825 0.57 6.955 0.7 ;
 RECT 6.825 1.845 6.955 1.975 ;
 RECT 6.2 0.565 6.33 0.695 ;
 RECT 5.685 0.57 5.815 0.7 ;
 RECT 5.685 1.48 5.815 1.61 ;
 RECT 6.21 2.375 6.34 2.505 ;
 RECT 0.2 0.36 0.33 0.49 ;
 RECT 0.2 0.62 0.33 0.75 ;
 RECT 0.2 1.71 0.33 1.84 ;
 RECT 2.77 2.515 2.9 2.645 ;
 RECT 2 1.52 2.13 1.65 ;
 RECT 5.305 1.705 5.435 1.835 ;
 RECT 5.305 0.6 5.435 0.73 ;
 RECT 4.745 0.6 4.875 0.73 ;
 RECT 4.17 0.6 4.3 0.73 ;
 RECT 4.17 1.48 4.3 1.61 ;
 RECT 15.28 1.475 15.41 1.605 ;
 RECT 14.675 1.255 14.805 1.385 ;
 RECT 14.63 0.505 14.76 0.635 ;
 RECT 12.925 2.525 13.055 2.655 ;
 RECT 16.035 0.785 16.165 0.915 ;
 RECT 18.155 0.795 18.285 0.925 ;
 RECT 17.395 0.505 17.525 0.635 ;
 RECT 16.92 1.415 17.05 1.545 ;
 RECT 16.92 0.505 17.05 0.635 ;
 RECT 16.36 1.415 16.49 1.545 ;
 RECT 8.99 0.575 9.12 0.705 ;
 RECT 9.515 2.34 9.645 2.47 ;
 RECT 6.065 0.91 6.195 1.04 ;
 RECT 11.46 2.05 11.59 2.18 ;
 RECT 11.46 0.615 11.59 0.745 ;
 RECT 12.755 2.065 12.885 2.195 ;
 RECT 8.99 1.675 9.12 1.805 ;
 RECT 6.94 2.525 7.07 2.655 ;
 RECT 16.055 1.595 16.185 1.725 ;
 RECT 15.61 0.785 15.74 0.915 ;
 RECT 1.095 0.12 1.225 0.25 ;
 RECT 18.9 1.44 19.03 1.57 ;
 RECT 11.635 0.965 11.765 1.095 ;
 RECT 0.2 1.97 0.33 2.1 ;
 RECT 0.2 2.23 0.33 2.36 ;
 RECT 15.28 0.225 15.41 0.355 ;
 RECT 4.575 1.25 4.705 1.38 ;
 RECT 16.36 0.505 16.49 0.635 ;
 RECT 10.04 0.555 10.17 0.685 ;
 RECT 7.385 2.01 7.515 2.14 ;
 RECT 7.525 1.21 7.655 1.34 ;
 RECT 7.385 0.605 7.515 0.735 ;
 RECT 7.945 0.605 8.075 0.735 ;
 LAYER M1 ;
 RECT 16.05 0.92 16.19 1.785 ;
 RECT 15.965 0.78 16.215 0.92 ;
 RECT 4.525 1.21 4.755 1.245 ;
 RECT 4.525 1.385 4.755 1.42 ;
 RECT 4.525 1.245 5.44 1.385 ;
 RECT 5.3 0.55 5.44 1.245 ;
 RECT 5.3 1.385 5.44 1.9 ;
 RECT 4.165 0.55 4.305 1.475 ;
 RECT 4.1 1.475 4.37 1.615 ;
 RECT 14.95 0.36 15.09 0.5 ;
 RECT 12.9 0.22 15.09 0.36 ;
 RECT 14.95 0.5 16.495 0.64 ;
 RECT 16.355 0.435 16.495 0.5 ;
 RECT 16.355 0.64 16.495 1.61 ;
 RECT 0.595 0.6 0.735 2.13 ;
 RECT 1.555 0.41 1.695 0.46 ;
 RECT 2.315 0.41 2.455 1.475 ;
 RECT 1.555 0.27 2.455 0.41 ;
 RECT 0.595 0.46 1.695 0.6 ;
 RECT 5.58 1.94 5.72 2.05 ;
 RECT 3.82 2.05 5.72 2.19 ;
 RECT 3.82 1.805 3.96 2.05 ;
 RECT 3.605 0.545 3.745 1.665 ;
 RECT 3.54 1.665 3.96 1.805 ;
 RECT 7.1 0.365 7.24 1.205 ;
 RECT 6.54 0.365 6.68 1.8 ;
 RECT 6.54 0.225 7.24 0.365 ;
 RECT 5.58 1.8 6.68 1.94 ;
 RECT 7.1 1.205 7.725 1.345 ;
 RECT 17.715 0.36 17.855 0.79 ;
 RECT 16.915 0.36 17.055 1.41 ;
 RECT 16.85 1.41 17.12 1.55 ;
 RECT 16.915 0.22 17.855 0.36 ;
 RECT 17.715 0.79 18.335 0.93 ;
 RECT 0.895 1.21 1.035 1.275 ;
 RECT 0.895 1.415 1.035 1.48 ;
 RECT 0.895 1.275 2.135 1.415 ;
 RECT 1.995 0.55 2.135 1.275 ;
 RECT 1.995 1.415 2.135 1.71 ;
 RECT 12.055 1.17 12.395 1.51 ;
 RECT 12.845 2.52 15.09 2.65 ;
 RECT 12.845 2.65 15.08 2.66 ;
 RECT 14.95 1.33 15.09 2.52 ;
 RECT 17.39 0.64 17.53 1.925 ;
 RECT 15.6 1.33 15.74 1.925 ;
 RECT 17.325 0.5 17.575 0.64 ;
 RECT 15.6 1.925 17.53 2.065 ;
 RECT 14.95 1.19 15.74 1.33 ;
 RECT 3.49 2.33 6 2.47 ;
 RECT 5.86 2.23 6 2.33 ;
 RECT 3.49 2.085 3.63 2.33 ;
 RECT 1.355 1.945 3.63 2.085 ;
 RECT 2.625 0.835 2.765 1.945 ;
 RECT 1.36 1.715 1.5 1.945 ;
 RECT 1.29 1.575 1.565 1.715 ;
 RECT 5.86 2.09 6.96 2.23 ;
 RECT 6.82 0.52 6.96 2.09 ;
 RECT 18.475 0.435 18.615 1.07 ;
 RECT 17.675 1.07 18.615 1.21 ;
 RECT 18.475 1.21 18.615 1.64 ;
 RECT 11.895 1.845 12.035 2.45 ;
 RECT 10.86 2.385 11 2.45 ;
 RECT 10.86 2.45 12.035 2.59 ;
 RECT 10.86 2.59 11 2.65 ;
 RECT 12.75 0.55 12.89 1.705 ;
 RECT 11.895 1.705 12.89 1.845 ;
 RECT 12.75 1.845 12.89 2.265 ;
 RECT 8.705 0.385 8.845 0.88 ;
 RECT 7.94 0.88 8.845 1.02 ;
 RECT 7.94 0.55 8.08 0.88 ;
 RECT 7.94 1.02 8.08 2.21 ;
 RECT 8.705 0.245 9.405 0.385 ;
 RECT 9.265 0.385 9.405 0.75 ;
 RECT 9.68 0.89 9.82 1.095 ;
 RECT 9.265 0.75 9.86 0.89 ;
 RECT 11.26 1.095 11.4 1.835 ;
 RECT 11.585 0.925 11.815 0.955 ;
 RECT 11.26 0.955 11.815 1.095 ;
 RECT 11.585 1.095 11.815 1.135 ;
 RECT 5.68 0.38 5.82 1.305 ;
 RECT 5.02 0.38 5.16 0.93 ;
 RECT 5.68 1.445 5.82 1.66 ;
 RECT 5.02 0.24 5.82 0.38 ;
 RECT 4.455 0.93 5.16 1.07 ;
 RECT 4.455 0.375 4.595 0.93 ;
 RECT 3.125 0.375 3.265 1.26 ;
 RECT 3.125 0.235 4.595 0.375 ;
 RECT 2.955 1.26 3.265 1.4 ;
 RECT 2.955 1.4 3.095 1.77 ;
 RECT 5.68 1.305 6.4 1.445 ;
 RECT 6.26 1.26 6.4 1.305 ;
 RECT 6.26 1.445 6.4 1.51 ;
 RECT 8.22 2.135 8.36 2.435 ;
 RECT 7.66 1.775 7.8 2.435 ;
 RECT 7.1 1.635 7.8 1.775 ;
 RECT 7.66 2.435 8.36 2.575 ;
 RECT 7.1 1.775 7.24 2.52 ;
 RECT 6.87 2.52 7.24 2.66 ;
 RECT 10.315 1.86 10.455 1.995 ;
 RECT 8.22 1.995 10.455 2.135 ;
 RECT 10.975 2.045 11.64 2.185 ;
 RECT 10.975 1.86 11.115 2.045 ;
 RECT 10.975 0.75 11.115 1.72 ;
 RECT 10.315 1.72 11.115 1.86 ;
 RECT 10.975 0.61 11.66 0.75 ;
 RECT 14.67 0.64 14.81 0.78 ;
 RECT 14.67 0.92 14.81 1.455 ;
 RECT 14.565 0.5 14.81 0.64 ;
 RECT 14.67 0.78 15.805 0.92 ;
 END
END RDFFX2

MACRO RSDFFX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 23.04 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 1.13 1.39 1.47 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.79 1.42 2.095 1.805 ;
 RECT 1.63 0.92 1.93 1.06 ;
 RECT 1.79 1.06 1.93 1.42 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.63 2.25 2.08 2.575 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.16 0.835 9.595 1.08 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.475 1.09 11.845 1.5 ;
 RECT 11.525 1.5 11.665 2.295 ;
 RECT 11.525 0.525 11.665 1.09 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.305 1.27 12.715 1.66 ;
 RECT 12.575 1.66 12.715 1.79 ;
 RECT 12.575 0.48 12.715 1.27 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 23.04 2.96 ;
 RECT 7.875 2.615 8.11 2.8 ;
 RECT 5.92 2.51 6.15 2.65 ;
 RECT 4.225 2.51 4.495 2.65 ;
 RECT 2.565 1.97 2.965 2.11 ;
 RECT 9.385 2.37 9.655 2.51 ;
 RECT 0.185 1.64 0.345 2.8 ;
 RECT 13.135 2 13.275 2.8 ;
 RECT 10.58 1.94 10.72 2.8 ;
 RECT 14.825 2.025 14.965 2.8 ;
 RECT 1.07 1.985 1.21 2.8 ;
 RECT 12.095 2.275 12.235 2.8 ;
 RECT 5.965 2.65 6.105 2.8 ;
 RECT 4.29 2.65 4.43 2.8 ;
 RECT 2.825 2.11 2.965 2.8 ;
 RECT 9.45 2.51 9.59 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 23.04 0.08 ;
 RECT 5.93 0.555 6.18 0.695 ;
 RECT 17.785 0.22 18.035 0.36 ;
 RECT 9.33 0.555 9.6 0.695 ;
 RECT 4.29 0.08 4.43 0.32 ;
 RECT 13.185 0.08 13.325 0.865 ;
 RECT 12.095 0.08 12.235 0.575 ;
 RECT 1.07 0.08 1.21 0.4 ;
 RECT 20.55 0.08 20.69 0.65 ;
 RECT 0.185 0.08 0.345 0.84 ;
 RECT 10.58 0.08 10.72 0.785 ;
 RECT 7.94 0.08 8.08 0.78 ;
 RECT 14.825 0.08 14.965 0.815 ;
 RECT 5.995 0.08 6.135 0.555 ;
 RECT 17.83 0.08 17.97 0.22 ;
 RECT 9.395 0.08 9.535 0.555 ;
 RECT 2.81 0.73 2.95 0.735 ;
 RECT 2.565 0.59 2.95 0.73 ;
 RECT 2.81 0.08 2.95 0.59 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 21.405 1.4 21.745 1.765 ;
 RECT 17.82 2.225 21.57 2.385 ;
 RECT 17.785 1.47 18.015 1.61 ;
 RECT 20.505 1.395 20.645 2.225 ;
 RECT 21.42 1.765 21.56 2.225 ;
 RECT 17.83 1.61 17.97 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 15.955 0.81 16.335 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 13.47 0.385 13.57 2.405 ;
 RECT 13.37 2.405 13.6 2.635 ;
 RECT 1.91 1.565 2.2 1.795 ;
 RECT 2.1 1.795 2.2 2.385 ;
 RECT 4.945 0.38 5.045 0.945 ;
 RECT 4.945 1.175 5.045 2.36 ;
 RECT 4.825 0.945 5.055 1.175 ;
 RECT 13.78 1.835 13.88 2.425 ;
 RECT 13.77 1.605 14 1.835 ;
 RECT 20.805 0.27 20.905 0.745 ;
 RECT 20.805 0.975 20.905 1.855 ;
 RECT 20.66 0.745 20.905 0.975 ;
 RECT 8.22 0.37 8.32 2.68 ;
 RECT 10.09 2.475 10.32 2.68 ;
 RECT 8.22 2.68 10.32 2.78 ;
 RECT 9.715 0.33 9.815 1.265 ;
 RECT 9.715 1.485 9.815 2.235 ;
 RECT 9.415 1.265 9.815 1.485 ;
 RECT 7.67 0.37 7.77 1.21 ;
 RECT 7.67 1.42 7.77 2.16 ;
 RECT 7.67 1.21 7.955 1.42 ;
 RECT 1.63 0.335 1.73 0.875 ;
 RECT 1.63 0.875 1.86 1.105 ;
 RECT 9.135 0.33 9.235 0.865 ;
 RECT 9.135 1.08 9.235 2.235 ;
 RECT 9.135 0.865 9.425 1.08 ;
 RECT 5.775 0.38 5.875 0.84 ;
 RECT 5.775 0.87 6.35 0.97 ;
 RECT 6.25 0.38 6.35 0.87 ;
 RECT 5.775 0.84 6.02 0.87 ;
 RECT 5.775 0.97 6.02 1.06 ;
 RECT 2.885 0.35 2.985 1.205 ;
 RECT 2.885 1.415 2.985 2.395 ;
 RECT 2.735 1.205 2.985 1.415 ;
 RECT 5.47 1.45 5.57 2.345 ;
 RECT 6.565 0.38 6.665 1.24 ;
 RECT 5.47 1.24 6.665 1.34 ;
 RECT 6.565 1.34 6.665 2.435 ;
 RECT 5.47 1.34 5.7 1.45 ;
 RECT 5.47 0.38 5.57 1.24 ;
 RECT 2.405 0.45 2.505 2.385 ;
 RECT 2.395 0.24 2.625 0.45 ;
 RECT 6.24 1.75 6.34 2.44 ;
 RECT 5.77 1.73 5.87 2.34 ;
 RECT 6.11 1.53 6.34 1.63 ;
 RECT 6.11 1.73 6.34 1.75 ;
 RECT 5.77 1.63 6.34 1.73 ;
 RECT 10.87 0.365 10.97 1.16 ;
 RECT 10.675 1.16 10.97 1.22 ;
 RECT 10.87 1.39 10.97 2.47 ;
 RECT 10.675 1.32 10.97 1.39 ;
 RECT 10.675 1.22 11.88 1.32 ;
 RECT 11.78 0.105 11.88 1.22 ;
 RECT 11.78 1.32 11.88 2.75 ;
 RECT 4.545 0.1 7.24 0.2 ;
 RECT 7.14 0.42 7.24 0.95 ;
 RECT 6.94 0.2 7.24 0.42 ;
 RECT 4.545 0.2 4.645 0.97 ;
 RECT 7.065 1.445 7.165 2.285 ;
 RECT 6.98 2.285 7.21 2.515 ;
 RECT 4.635 1.76 4.735 2.34 ;
 RECT 4.515 1.53 4.745 1.76 ;
 RECT 14.31 2.605 15.66 2.695 ;
 RECT 15.43 2.475 15.66 2.605 ;
 RECT 14.31 1.425 14.41 2.605 ;
 RECT 13.775 0.385 13.875 1.325 ;
 RECT 14.315 2.695 15.66 2.705 ;
 RECT 13.775 1.325 14.41 1.425 ;
 RECT 1.195 1.165 1.425 1.23 ;
 RECT 1.195 1.33 1.425 1.395 ;
 RECT 0.855 1.23 1.425 1.33 ;
 RECT 1.325 0.345 1.425 1.165 ;
 RECT 1.325 1.395 1.425 2.385 ;
 RECT 0.855 0.345 0.955 1.23 ;
 RECT 0.855 1.33 0.955 2.385 ;
 RECT 4.05 0.38 4.15 1.23 ;
 RECT 4.05 1.46 4.15 2.34 ;
 RECT 4.05 1.23 4.28 1.46 ;
 RECT 14.61 0.385 14.71 1.215 ;
 RECT 14.61 1.215 14.885 1.27 ;
 RECT 14.61 1.425 14.71 2.425 ;
 RECT 14.61 1.37 14.885 1.425 ;
 RECT 15.085 1.045 15.185 1.27 ;
 RECT 15.085 1.37 15.185 2.425 ;
 RECT 14.61 1.27 15.185 1.37 ;
 RECT 17.535 1.045 17.635 1.76 ;
 RECT 16.045 0.84 16.275 0.945 ;
 RECT 16.045 1.045 16.275 1.07 ;
 RECT 15.085 0.385 15.185 0.945 ;
 RECT 15.085 0.945 17.635 1.045 ;
 RECT 17.535 0.145 17.635 0.945 ;
 RECT 19.725 1.145 19.825 2.09 ;
 RECT 18.69 1.86 18.79 2.09 ;
 RECT 18.56 1.545 18.79 1.76 ;
 RECT 17.535 1.76 18.79 1.86 ;
 RECT 18.69 2.09 19.825 2.19 ;
 RECT 20.2 0.275 20.3 1.025 ;
 RECT 20.2 1.255 20.3 1.86 ;
 RECT 20.2 1.025 20.48 1.255 ;
 RECT 18.115 0.965 18.215 1.145 ;
 RECT 18.115 1.145 19.545 1.245 ;
 RECT 19.445 0.965 19.545 1.145 ;
 RECT 19.255 1.245 19.355 1.86 ;
 RECT 19.725 0.275 19.825 0.865 ;
 RECT 18.115 0.735 18.345 0.965 ;
 RECT 19.445 0.865 19.825 0.965 ;
 RECT 18.54 0.865 19.265 0.965 ;
 RECT 18.54 0.735 18.77 0.865 ;
 RECT 19.165 0.275 19.265 0.865 ;
 RECT 14.265 0.205 14.365 0.925 ;
 RECT 12.36 0.205 12.46 0.87 ;
 RECT 12.215 0.87 12.46 1.085 ;
 RECT 12.36 1.085 12.46 2.755 ;
 RECT 12.36 0.105 15.735 0.205 ;
 RECT 15.505 0.205 15.735 0.4 ;
 RECT 14.14 0.925 14.37 1.135 ;
 RECT 1.63 1.385 1.73 2.365 ;
 RECT 2.1 0.365 2.2 1.285 ;
 RECT 1.63 1.285 2.2 1.385 ;
 RECT 1.63 2.365 1.86 2.575 ;
 LAYER CO ;
 RECT 0.2 0.62 0.33 0.75 ;
 RECT 0.2 1.71 0.33 1.84 ;
 RECT 0.2 1.97 0.33 2.1 ;
 RECT 0.2 2.23 0.33 2.36 ;
 RECT 17.835 0.225 17.965 0.355 ;
 RECT 1.68 2.405 1.81 2.535 ;
 RECT 6.81 1.67 6.94 1.8 ;
 RECT 4.295 2.515 4.425 2.645 ;
 RECT 5.97 2.515 6.1 2.645 ;
 RECT 5.2 1.52 5.33 1.65 ;
 RECT 6 0.555 6.13 0.685 ;
 RECT 5.2 0.6 5.33 0.73 ;
 RECT 3.11 1.975 3.24 2.105 ;
 RECT 3.11 0.595 3.24 0.725 ;
 RECT 2.635 0.595 2.765 0.725 ;
 RECT 2.635 1.975 2.765 2.105 ;
 RECT 17.835 1.475 17.965 1.605 ;
 RECT 17.23 1.255 17.36 1.385 ;
 RECT 17.185 0.505 17.315 0.635 ;
 RECT 15.48 2.525 15.61 2.655 ;
 RECT 13.42 2.455 13.55 2.585 ;
 RECT 14.015 0.635 14.145 0.765 ;
 RECT 13.19 0.635 13.32 0.765 ;
 RECT 13.14 2.06 13.27 2.19 ;
 RECT 15.31 2.065 15.44 2.195 ;
 RECT 11.53 1.715 11.66 1.845 ;
 RECT 10.14 2.525 10.27 2.655 ;
 RECT 11.53 0.585 11.66 0.715 ;
 RECT 11.53 2.105 11.66 2.235 ;
 RECT 12.1 2.34 12.23 2.47 ;
 RECT 14.705 1.255 14.835 1.385 ;
 RECT 14.19 0.965 14.32 1.095 ;
 RECT 18.59 0.785 18.72 0.915 ;
 RECT 20.71 0.795 20.84 0.925 ;
 RECT 20.3 1.075 20.43 1.205 ;
 RECT 21.035 0.505 21.165 0.635 ;
 RECT 21.035 1.44 21.165 1.57 ;
 RECT 20.555 0.47 20.685 0.6 ;
 RECT 20.51 1.455 20.64 1.585 ;
 RECT 19.95 1.435 20.08 1.565 ;
 RECT 19.95 0.505 20.08 0.635 ;
 RECT 19.475 1.415 19.605 1.545 ;
 RECT 19.475 0.505 19.605 0.635 ;
 RECT 18.915 1.415 19.045 1.545 ;
 RECT 18.915 0.505 19.045 0.635 ;
 RECT 12.58 0.555 12.71 0.685 ;
 RECT 10.585 2.01 10.715 2.14 ;
 RECT 10.725 1.21 10.855 1.34 ;
 RECT 10.585 0.605 10.715 0.735 ;
 RECT 11.145 2.025 11.275 2.155 ;
 RECT 11.145 0.605 11.275 0.735 ;
 RECT 9.245 0.91 9.375 1.04 ;
 RECT 12.58 1.6 12.71 1.73 ;
 RECT 12.1 0.395 12.23 0.525 ;
 RECT 9.465 1.305 9.595 1.435 ;
 RECT 7.03 2.335 7.16 2.465 ;
 RECT 6.99 0.24 7.12 0.37 ;
 RECT 7.775 1.25 7.905 1.38 ;
 RECT 2.785 1.245 2.915 1.375 ;
 RECT 6.16 1.57 6.29 1.7 ;
 RECT 5.83 0.89 5.96 1.02 ;
 RECT 5.52 1.28 5.65 1.41 ;
 RECT 18.61 1.595 18.74 1.725 ;
 RECT 18.165 0.785 18.295 0.915 ;
 RECT 4.295 0.12 4.425 0.25 ;
 RECT 21.455 1.44 21.585 1.57 ;
 RECT 0.2 0.36 0.33 0.49 ;
 RECT 4.565 1.58 4.695 1.71 ;
 RECT 4.875 0.995 5.005 1.125 ;
 RECT 4.1 1.28 4.23 1.41 ;
 RECT 1.68 0.925 1.81 1.055 ;
 RECT 1.68 0.925 1.81 1.055 ;
 RECT 1.245 1.215 1.375 1.345 ;
 RECT 1.96 1.615 2.09 1.745 ;
 RECT 10.025 0.57 10.155 0.7 ;
 RECT 10.025 1.64 10.155 1.77 ;
 RECT 9.4 0.56 9.53 0.69 ;
 RECT 8.885 0.57 9.015 0.7 ;
 RECT 8.885 1.48 9.015 1.61 ;
 RECT 9.455 2.375 9.585 2.505 ;
 RECT 7.93 2.63 8.06 2.76 ;
 RECT 3.48 1.935 3.61 2.065 ;
 RECT 3.68 0.6 3.81 0.73 ;
 RECT 1.075 2.035 1.205 2.165 ;
 RECT 8.505 1.705 8.635 1.835 ;
 RECT 8.505 0.6 8.635 0.73 ;
 RECT 7.945 0.6 8.075 0.73 ;
 RECT 7.37 0.6 7.5 0.73 ;
 RECT 7.37 1.48 7.5 1.61 ;
 RECT 6.81 0.6 6.94 0.73 ;
 RECT 1.85 1.975 1.98 2.105 ;
 RECT 1.85 0.595 1.98 0.725 ;
 RECT 1.075 0.16 1.205 0.29 ;
 RECT 0.605 0.595 0.735 0.725 ;
 RECT 0.605 1.975 0.735 2.105 ;
 RECT 15.555 0.225 15.685 0.355 ;
 RECT 13.82 1.655 13.95 1.785 ;
 RECT 15.31 0.635 15.44 0.765 ;
 RECT 14.83 0.635 14.96 0.765 ;
 RECT 14.83 2.075 14.96 2.205 ;
 RECT 14.015 2.05 14.145 2.18 ;
 RECT 12.265 0.915 12.395 1.045 ;
 RECT 2.445 0.28 2.575 0.41 ;
 RECT 16.095 0.89 16.225 1.02 ;
 LAYER M1 ;
 RECT 7.725 1.21 7.955 1.245 ;
 RECT 7.725 1.385 7.955 1.42 ;
 RECT 7.725 1.245 8.64 1.385 ;
 RECT 8.5 0.55 8.64 1.245 ;
 RECT 8.5 1.385 8.64 1.9 ;
 RECT 14.14 0.925 14.37 0.955 ;
 RECT 13.815 0.955 14.37 1.095 ;
 RECT 14.14 1.095 14.37 1.135 ;
 RECT 13.815 1.095 13.955 1.835 ;
 RECT 11.14 0.385 11.28 2.21 ;
 RECT 11.805 0.385 11.945 0.75 ;
 RECT 11.14 0.245 11.945 0.385 ;
 RECT 12.26 0.89 12.4 1.095 ;
 RECT 11.805 0.75 12.4 0.89 ;
 RECT 7.365 0.55 7.505 1.475 ;
 RECT 7.3 1.475 7.57 1.615 ;
 RECT 14.45 1.845 14.59 2.45 ;
 RECT 13.415 2.385 13.555 2.45 ;
 RECT 13.415 2.45 14.59 2.59 ;
 RECT 13.415 2.59 13.555 2.65 ;
 RECT 15.305 0.585 15.445 1.705 ;
 RECT 14.45 1.705 15.445 1.845 ;
 RECT 15.305 1.845 15.445 2.265 ;
 RECT 17.505 0.36 17.645 0.5 ;
 RECT 15.455 0.22 17.645 0.36 ;
 RECT 17.505 0.5 19.05 0.64 ;
 RECT 18.91 0.435 19.05 0.5 ;
 RECT 18.91 0.64 19.05 1.61 ;
 RECT 0.6 0.545 0.74 0.58 ;
 RECT 0.6 0.72 0.74 2.155 ;
 RECT 1.37 0.38 1.51 0.58 ;
 RECT 0.6 0.58 1.51 0.72 ;
 RECT 1.37 0.25 2.655 0.38 ;
 RECT 1.38 0.24 2.655 0.25 ;
 RECT 2.3 0.38 2.655 0.45 ;
 RECT 2.235 0.73 2.375 1.24 ;
 RECT 2.235 1.38 2.375 1.97 ;
 RECT 1.78 1.97 2.375 2.11 ;
 RECT 1.78 0.59 2.375 0.73 ;
 RECT 2.735 1.205 2.965 1.24 ;
 RECT 2.235 1.24 2.965 1.38 ;
 RECT 2.735 1.38 2.965 1.415 ;
 RECT 15.4 2.52 17.645 2.65 ;
 RECT 15.4 2.65 17.635 2.66 ;
 RECT 17.505 1.33 17.645 2.52 ;
 RECT 19.945 0.64 20.085 1.925 ;
 RECT 18.155 1.33 18.295 1.925 ;
 RECT 19.88 0.5 20.13 0.64 ;
 RECT 17.505 1.19 18.295 1.33 ;
 RECT 18.155 1.925 20.085 2.065 ;
 RECT 3.77 1.13 3.91 2.42 ;
 RECT 3.105 1.975 3.25 2.155 ;
 RECT 3.105 0.505 3.245 1.975 ;
 RECT 3.11 2.155 3.25 2.42 ;
 RECT 3.11 2.42 3.91 2.56 ;
 RECT 3.77 0.99 5.055 1.13 ;
 RECT 17.225 0.64 17.365 0.78 ;
 RECT 17.225 0.92 17.365 1.455 ;
 RECT 17.225 0.78 18.36 0.92 ;
 RECT 17.12 0.5 17.365 0.64 ;
 RECT 18.605 0.92 18.745 1.785 ;
 RECT 18.52 0.78 18.77 0.92 ;
 RECT 5.195 0.55 5.335 1.275 ;
 RECT 4.05 1.275 5.335 1.415 ;
 RECT 5.195 1.415 5.335 1.71 ;
 RECT 20.27 0.36 20.41 0.79 ;
 RECT 19.47 0.36 19.61 1.41 ;
 RECT 19.405 1.41 19.675 1.55 ;
 RECT 19.47 0.22 20.41 0.36 ;
 RECT 20.27 0.79 20.89 0.93 ;
 RECT 3.475 0.6 3.88 0.735 ;
 RECT 3.475 0.735 3.615 2.13 ;
 RECT 4.755 0.6 4.895 0.61 ;
 RECT 4.755 0.41 4.895 0.46 ;
 RECT 3.475 0.595 4.895 0.6 ;
 RECT 3.68 0.46 4.895 0.595 ;
 RECT 4.755 0.275 5.655 0.41 ;
 RECT 5.515 0.41 5.655 1.475 ;
 RECT 4.755 0.27 5.59 0.275 ;
 RECT 6.69 2.085 6.83 2.33 ;
 RECT 4.555 1.945 6.83 2.085 ;
 RECT 5.825 0.835 5.965 1.945 ;
 RECT 4.56 1.715 4.7 1.945 ;
 RECT 4.49 1.575 4.765 1.715 ;
 RECT 6.69 2.33 9.2 2.47 ;
 RECT 9.06 2.23 9.2 2.33 ;
 RECT 9.06 2.09 10.16 2.23 ;
 RECT 10.02 0.52 10.16 2.09 ;
 RECT 10.86 1.775 11 2.435 ;
 RECT 10.3 1.635 11 1.775 ;
 RECT 10.3 1.775 10.44 2.52 ;
 RECT 10.07 2.52 10.44 2.66 ;
 RECT 10.86 2.435 11.955 2.575 ;
 RECT 11.815 2.135 11.955 2.435 ;
 RECT 12.855 1.86 12.995 1.995 ;
 RECT 11.815 1.995 12.995 2.135 ;
 RECT 13.53 2.045 14.195 2.185 ;
 RECT 13.53 1.86 13.67 2.045 ;
 RECT 13.53 0.63 14.195 0.77 ;
 RECT 13.53 0.77 13.67 1.72 ;
 RECT 12.855 1.72 13.67 1.86 ;
 RECT 8.22 0.38 8.36 0.93 ;
 RECT 8.88 0.38 9.02 1.3 ;
 RECT 8.22 0.24 9.02 0.38 ;
 RECT 8.88 1.44 9.02 1.66 ;
 RECT 7.655 0.93 8.36 1.07 ;
 RECT 6.325 0.375 6.465 1.26 ;
 RECT 7.655 0.375 7.795 0.93 ;
 RECT 6.155 1.26 6.465 1.4 ;
 RECT 6.155 1.4 6.295 1.77 ;
 RECT 6.325 0.235 7.795 0.375 ;
 RECT 9.46 1.255 9.6 1.3 ;
 RECT 9.46 1.44 9.6 1.49 ;
 RECT 8.88 1.3 9.6 1.44 ;
 RECT 21.03 0.435 21.17 1.07 ;
 RECT 20.23 1.07 21.17 1.21 ;
 RECT 21.03 1.21 21.17 1.64 ;
 RECT 8.78 1.94 8.92 2.05 ;
 RECT 7.02 2.05 8.92 2.19 ;
 RECT 7.02 1.805 7.16 2.05 ;
 RECT 6.805 0.545 6.945 1.665 ;
 RECT 6.735 1.665 7.16 1.805 ;
 RECT 9.74 0.365 9.88 1.8 ;
 RECT 10.3 0.365 10.44 1.205 ;
 RECT 9.74 0.225 10.44 0.365 ;
 RECT 8.78 1.8 9.88 1.94 ;
 RECT 10.3 1.205 10.925 1.345 ;
 RECT 14.61 1.17 14.95 1.51 ;
 END
END RSDFFX1

MACRO RSDFFX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 23.68 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.965 1.13 1.39 1.47 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.63 0.92 1.865 1.06 ;
 RECT 1.645 1.445 2.095 1.495 ;
 RECT 1.65 1.495 2.095 1.805 ;
 RECT 1.645 1.06 1.785 1.445 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.63 2.23 2.08 2.55 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.185 1.09 12.455 1.5 ;
 RECT 12.185 1.5 12.325 1.855 ;
 RECT 12.185 0.525 12.325 1.09 ;
 END
 ANTENNADIFFAREA 0.584 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.235 1.595 13.375 1.855 ;
 RECT 12.955 1.295 13.375 1.595 ;
 RECT 13.235 0.48 13.375 1.295 ;
 END
 ANTENNADIFFAREA 0.6 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 23.68 2.96 ;
 RECT 7.875 2.615 8.11 2.8 ;
 RECT 9.34 2.37 9.61 2.51 ;
 RECT 2.565 1.97 2.965 2.11 ;
 RECT 5.92 2.51 6.15 2.65 ;
 RECT 4.225 2.51 4.495 2.65 ;
 RECT 15.47 2.025 15.61 2.8 ;
 RECT 1.07 1.985 1.21 2.8 ;
 RECT 12.71 2.275 12.85 2.8 ;
 RECT 0.185 1.64 0.345 2.8 ;
 RECT 11.705 2.275 11.845 2.8 ;
 RECT 13.715 2.275 13.855 2.8 ;
 RECT 10.58 1.94 10.72 2.8 ;
 RECT 9.405 2.51 9.545 2.8 ;
 RECT 2.825 2.11 2.965 2.8 ;
 RECT 5.965 2.65 6.105 2.8 ;
 RECT 4.29 2.65 4.43 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 23.68 0.08 ;
 RECT 9.33 0.555 9.6 0.695 ;
 RECT 5.93 0.555 6.18 0.695 ;
 RECT 18.43 0.22 18.68 0.36 ;
 RECT 15.47 0.08 15.61 0.815 ;
 RECT 12.755 0.08 12.895 0.575 ;
 RECT 7.94 0.08 8.08 0.78 ;
 RECT 1.07 0.08 1.21 0.355 ;
 RECT 21.195 0.08 21.335 0.65 ;
 RECT 0.185 0.08 0.345 0.84 ;
 RECT 11.625 0.08 11.765 0.575 ;
 RECT 4.29 0.08 4.43 0.32 ;
 RECT 10.58 0.08 10.72 0.785 ;
 RECT 13.71 0.08 13.85 0.575 ;
 RECT 9.395 0.08 9.535 0.555 ;
 RECT 5.995 0.08 6.135 0.555 ;
 RECT 18.475 0.08 18.615 0.22 ;
 RECT 2.82 0.08 2.96 0.59 ;
 RECT 2.565 0.59 2.96 0.73 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 22.05 1.4 22.39 1.765 ;
 RECT 18.475 2.225 22.205 2.385 ;
 RECT 18.43 1.47 18.66 1.61 ;
 RECT 21.15 1.395 21.29 2.225 ;
 RECT 22.065 1.765 22.205 2.225 ;
 RECT 18.475 1.61 18.615 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 16.6 0.76 16.98 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.22 0.84 9.56 1.12 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END CLK

 OBS
 LAYER PO ;
 RECT 9.135 0.33 9.235 0.86 ;
 RECT 9.135 1.09 9.235 2.235 ;
 RECT 9.135 0.86 9.445 1.09 ;
 RECT 14.425 1.835 14.525 2.425 ;
 RECT 14.415 1.605 14.645 1.835 ;
 RECT 7.065 1.445 7.165 2.285 ;
 RECT 6.98 2.285 7.21 2.515 ;
 RECT 4.945 0.38 5.045 0.945 ;
 RECT 4.945 1.175 5.045 2.36 ;
 RECT 4.825 0.945 5.055 1.175 ;
 RECT 21.45 0.27 21.55 0.745 ;
 RECT 21.45 0.975 21.55 1.855 ;
 RECT 21.305 0.745 21.55 0.975 ;
 RECT 4.635 1.76 4.735 2.34 ;
 RECT 4.515 1.53 4.745 1.76 ;
 RECT 20.845 0.275 20.945 1.025 ;
 RECT 20.845 1.255 20.945 1.86 ;
 RECT 20.845 1.025 21.125 1.255 ;
 RECT 4.05 0.38 4.15 1.23 ;
 RECT 4.05 1.46 4.15 2.34 ;
 RECT 4.05 1.23 4.28 1.46 ;
 RECT 0.855 0.345 0.955 1.23 ;
 RECT 0.855 1.33 0.955 2.385 ;
 RECT 0.855 1.23 1.425 1.33 ;
 RECT 1.195 1.165 1.425 1.23 ;
 RECT 1.195 1.33 1.425 1.395 ;
 RECT 1.325 0.345 1.425 1.165 ;
 RECT 1.325 1.395 1.425 2.385 ;
 RECT 19.185 0.865 19.91 0.965 ;
 RECT 19.185 0.735 19.415 0.865 ;
 RECT 19.81 0.275 19.91 0.865 ;
 RECT 5.47 1.34 5.7 1.45 ;
 RECT 5.47 0.38 5.57 1.24 ;
 RECT 5.47 1.45 5.57 2.345 ;
 RECT 6.565 0.38 6.665 1.24 ;
 RECT 6.565 1.34 6.665 2.475 ;
 RECT 5.47 1.24 6.665 1.34 ;
 RECT 8.22 0.37 8.32 2.68 ;
 RECT 10.09 2.475 10.32 2.68 ;
 RECT 8.22 2.68 10.32 2.78 ;
 RECT 5.775 0.84 6.02 0.87 ;
 RECT 5.775 0.97 6.02 1.06 ;
 RECT 5.775 0.38 5.875 0.84 ;
 RECT 6.25 0.38 6.35 0.87 ;
 RECT 5.775 0.87 6.35 0.97 ;
 RECT 9.675 0.33 9.775 1.27 ;
 RECT 9.675 1.49 9.775 2.235 ;
 RECT 9.415 1.27 9.775 1.49 ;
 RECT 7.67 0.37 7.77 1.21 ;
 RECT 7.67 1.42 7.77 2.16 ;
 RECT 7.67 1.21 7.955 1.42 ;
 RECT 1.63 0.335 1.73 0.875 ;
 RECT 1.63 0.875 1.86 1.105 ;
 RECT 6.24 1.75 6.34 2.48 ;
 RECT 6.11 1.53 6.34 1.63 ;
 RECT 6.11 1.73 6.34 1.75 ;
 RECT 5.77 1.73 5.87 2.34 ;
 RECT 5.77 1.63 6.34 1.73 ;
 RECT 14.42 0.385 14.52 1.325 ;
 RECT 14.955 2.605 16.305 2.695 ;
 RECT 16.075 2.475 16.305 2.605 ;
 RECT 14.955 1.425 15.055 2.605 ;
 RECT 14.42 1.325 15.055 1.425 ;
 RECT 14.96 2.695 16.305 2.705 ;
 RECT 1.91 1.565 2.2 1.795 ;
 RECT 2.1 1.795 2.2 2.385 ;
 RECT 13.02 0.105 13.12 0.87 ;
 RECT 12.875 0.87 13.12 0.88 ;
 RECT 12.875 0.88 13.59 0.98 ;
 RECT 13.49 0.205 13.59 0.88 ;
 RECT 14.91 0.205 15.01 0.925 ;
 RECT 13.02 1.085 13.12 1.23 ;
 RECT 13.02 1.23 13.59 1.33 ;
 RECT 13.02 1.33 13.12 2.755 ;
 RECT 13.49 1.33 13.59 2.77 ;
 RECT 12.875 0.98 13.12 1.085 ;
 RECT 16.15 0.205 16.38 0.4 ;
 RECT 13.49 0.105 16.38 0.205 ;
 RECT 14.785 0.925 15.015 1.135 ;
 RECT 12.44 0.98 12.54 1.22 ;
 RECT 10.675 1.22 12.54 1.32 ;
 RECT 12.44 1.32 12.54 2.75 ;
 RECT 10.87 0.365 10.97 1.16 ;
 RECT 10.675 1.16 10.97 1.22 ;
 RECT 10.87 1.39 10.97 2.47 ;
 RECT 10.675 1.32 10.97 1.39 ;
 RECT 11.97 0.095 12.07 0.88 ;
 RECT 12.44 0.105 12.54 0.88 ;
 RECT 11.97 1.32 12.07 2.77 ;
 RECT 11.97 0.88 12.54 0.98 ;
 RECT 4.545 0.1 7.24 0.2 ;
 RECT 7.14 0.42 7.24 0.95 ;
 RECT 6.94 0.2 7.24 0.42 ;
 RECT 4.545 0.2 4.645 0.97 ;
 RECT 18.18 0.145 18.28 0.945 ;
 RECT 18.18 1.045 18.28 1.76 ;
 RECT 15.255 0.385 15.355 1.215 ;
 RECT 15.255 1.215 15.53 1.27 ;
 RECT 15.255 1.425 15.355 2.425 ;
 RECT 15.255 1.37 15.53 1.425 ;
 RECT 15.73 1.045 15.83 1.27 ;
 RECT 15.255 1.27 15.83 1.37 ;
 RECT 15.73 1.37 15.83 2.425 ;
 RECT 20.37 1.145 20.47 2.09 ;
 RECT 19.335 1.86 19.435 2.09 ;
 RECT 19.205 1.545 19.435 1.76 ;
 RECT 16.69 0.84 16.92 0.945 ;
 RECT 16.69 1.045 16.92 1.07 ;
 RECT 15.73 0.385 15.83 0.945 ;
 RECT 15.73 0.945 18.28 1.045 ;
 RECT 19.335 2.09 20.47 2.19 ;
 RECT 18.18 1.76 19.435 1.86 ;
 RECT 18.76 0.965 18.86 1.145 ;
 RECT 20.37 0.275 20.47 0.865 ;
 RECT 18.76 1.145 20.19 1.245 ;
 RECT 20.09 0.965 20.19 1.145 ;
 RECT 19.9 1.245 20 1.86 ;
 RECT 18.76 0.735 18.99 0.965 ;
 RECT 20.09 0.865 20.47 0.965 ;
 RECT 1.63 1.385 1.73 2.34 ;
 RECT 2.1 0.365 2.2 1.285 ;
 RECT 1.63 1.285 2.2 1.385 ;
 RECT 1.63 2.34 1.86 2.55 ;
 RECT 14.115 0.385 14.215 2.405 ;
 RECT 14.015 2.405 14.245 2.635 ;
 RECT 2.885 0.35 2.985 1.205 ;
 RECT 2.885 1.415 2.985 2.395 ;
 RECT 2.735 1.205 2.985 1.415 ;
 RECT 2.405 0.43 2.505 2.385 ;
 RECT 2.395 0.22 2.625 0.43 ;
 LAYER CO ;
 RECT 9.265 0.91 9.395 1.04 ;
 RECT 13.715 0.395 13.845 0.525 ;
 RECT 13.72 2.34 13.85 2.47 ;
 RECT 11.63 0.395 11.76 0.525 ;
 RECT 11.71 2.34 11.84 2.47 ;
 RECT 19.235 0.785 19.365 0.915 ;
 RECT 21.355 0.795 21.485 0.925 ;
 RECT 20.945 1.075 21.075 1.205 ;
 RECT 21.68 0.505 21.81 0.635 ;
 RECT 21.68 1.44 21.81 1.57 ;
 RECT 21.2 0.47 21.33 0.6 ;
 RECT 21.155 1.455 21.285 1.585 ;
 RECT 20.595 1.435 20.725 1.565 ;
 RECT 20.595 0.505 20.725 0.635 ;
 RECT 20.12 1.415 20.25 1.545 ;
 RECT 20.12 0.505 20.25 0.635 ;
 RECT 19.56 1.415 19.69 1.545 ;
 RECT 19.56 0.505 19.69 0.635 ;
 RECT 13.24 0.555 13.37 0.685 ;
 RECT 10.585 2.01 10.715 2.14 ;
 RECT 10.725 1.21 10.855 1.34 ;
 RECT 10.585 0.605 10.715 0.735 ;
 RECT 11.145 2.025 11.275 2.155 ;
 RECT 11.145 0.605 11.275 0.735 ;
 RECT 9.465 1.31 9.595 1.44 ;
 RECT 7.03 2.335 7.16 2.465 ;
 RECT 6.99 0.24 7.12 0.37 ;
 RECT 6.16 1.57 6.29 1.7 ;
 RECT 5.83 0.89 5.96 1.02 ;
 RECT 5.52 1.28 5.65 1.41 ;
 RECT 4.565 1.58 4.695 1.71 ;
 RECT 4.875 0.995 5.005 1.125 ;
 RECT 4.1 1.28 4.23 1.41 ;
 RECT 1.68 0.925 1.81 1.055 ;
 RECT 1.68 0.925 1.81 1.055 ;
 RECT 1.245 1.215 1.375 1.345 ;
 RECT 1.96 1.615 2.09 1.745 ;
 RECT 10.025 0.57 10.155 0.7 ;
 RECT 10.025 1.845 10.155 1.975 ;
 RECT 9.4 0.56 9.53 0.69 ;
 RECT 8.885 0.57 9.015 0.7 ;
 RECT 8.885 1.48 9.015 1.61 ;
 RECT 9.41 2.375 9.54 2.505 ;
 RECT 7.93 2.63 8.06 2.76 ;
 RECT 3.48 1.935 3.61 2.065 ;
 RECT 3.68 0.6 3.81 0.73 ;
 RECT 6.81 1.67 6.94 1.8 ;
 RECT 4.295 2.515 4.425 2.645 ;
 RECT 5.97 2.515 6.1 2.645 ;
 RECT 5.2 1.52 5.33 1.65 ;
 RECT 1.075 2.035 1.205 2.165 ;
 RECT 8.505 1.705 8.635 1.835 ;
 RECT 8.505 0.6 8.635 0.73 ;
 RECT 7.945 0.6 8.075 0.73 ;
 RECT 7.37 0.6 7.5 0.73 ;
 RECT 7.37 1.48 7.5 1.61 ;
 RECT 6.81 0.6 6.94 0.73 ;
 RECT 6 0.555 6.13 0.685 ;
 RECT 5.2 0.6 5.33 0.73 ;
 RECT 3.11 1.975 3.24 2.105 ;
 RECT 3.11 0.595 3.24 0.725 ;
 RECT 2.635 0.595 2.765 0.725 ;
 RECT 2.635 1.975 2.765 2.105 ;
 RECT 1.85 1.955 1.98 2.085 ;
 RECT 1.85 0.595 1.98 0.725 ;
 RECT 1.075 0.15 1.205 0.28 ;
 RECT 0.605 0.595 0.735 0.725 ;
 RECT 0.605 1.975 0.735 2.105 ;
 RECT 16.2 0.225 16.33 0.355 ;
 RECT 18.48 1.475 18.61 1.605 ;
 RECT 17.875 1.255 18.005 1.385 ;
 RECT 17.83 0.505 17.96 0.635 ;
 RECT 16.125 2.525 16.255 2.655 ;
 RECT 14.065 2.455 14.195 2.585 ;
 RECT 14.465 1.655 14.595 1.785 ;
 RECT 15.955 0.615 16.085 0.745 ;
 RECT 15.475 0.615 15.605 0.745 ;
 RECT 15.475 2.075 15.605 2.205 ;
 RECT 14.66 2.05 14.79 2.18 ;
 RECT 14.66 0.615 14.79 0.745 ;
 RECT 15.955 2.065 16.085 2.195 ;
 RECT 12.19 1.675 12.32 1.805 ;
 RECT 10.14 2.525 10.27 2.655 ;
 RECT 12.925 0.915 13.055 1.045 ;
 RECT 13.24 1.675 13.37 1.805 ;
 RECT 12.76 0.395 12.89 0.525 ;
 RECT 12.19 0.585 12.32 0.715 ;
 RECT 12.715 2.34 12.845 2.47 ;
 RECT 15.35 1.255 15.48 1.385 ;
 RECT 14.835 0.965 14.965 1.095 ;
 RECT 2.445 0.26 2.575 0.39 ;
 RECT 7.775 1.25 7.905 1.38 ;
 RECT 2.785 1.245 2.915 1.375 ;
 RECT 16.74 0.89 16.87 1.02 ;
 RECT 19.255 1.595 19.385 1.725 ;
 RECT 18.81 0.785 18.94 0.915 ;
 RECT 4.295 0.12 4.425 0.25 ;
 RECT 22.1 1.44 22.23 1.57 ;
 RECT 0.2 0.36 0.33 0.49 ;
 RECT 0.2 0.62 0.33 0.75 ;
 RECT 0.2 1.71 0.33 1.84 ;
 RECT 0.2 1.97 0.33 2.1 ;
 RECT 0.2 2.23 0.33 2.36 ;
 RECT 18.48 0.225 18.61 0.355 ;
 RECT 1.68 2.38 1.81 2.51 ;
 LAYER M1 ;
 RECT 17.87 0.64 18.01 0.78 ;
 RECT 17.87 0.92 18.01 1.455 ;
 RECT 17.87 0.78 19.005 0.92 ;
 RECT 17.765 0.5 18.01 0.64 ;
 RECT 19.25 0.92 19.39 1.785 ;
 RECT 19.165 0.78 19.415 0.92 ;
 RECT 18.15 0.36 18.29 0.5 ;
 RECT 16.1 0.22 18.29 0.36 ;
 RECT 19.555 0.435 19.695 0.5 ;
 RECT 19.555 0.64 19.695 1.61 ;
 RECT 18.15 0.5 19.695 0.64 ;
 RECT 7.365 0.55 7.505 1.475 ;
 RECT 7.3 1.475 7.57 1.615 ;
 RECT 7.725 1.21 7.955 1.245 ;
 RECT 7.725 1.385 7.955 1.42 ;
 RECT 7.725 1.245 8.64 1.385 ;
 RECT 8.5 0.55 8.64 1.245 ;
 RECT 8.5 1.385 8.64 1.9 ;
 RECT 0.6 0.545 0.74 0.57 ;
 RECT 0.6 0.71 0.74 2.155 ;
 RECT 1.365 0.36 1.505 0.57 ;
 RECT 0.6 0.57 1.51 0.71 ;
 RECT 2.275 0.36 2.625 0.43 ;
 RECT 1.365 0.22 2.625 0.36 ;
 RECT 11.905 0.385 12.045 0.88 ;
 RECT 11.14 0.88 12.045 1.02 ;
 RECT 11.14 0.55 11.28 0.88 ;
 RECT 11.14 1.02 11.28 2.21 ;
 RECT 12.465 0.385 12.605 0.75 ;
 RECT 11.905 0.245 12.605 0.385 ;
 RECT 12.92 0.89 13.06 1.095 ;
 RECT 12.465 0.75 13.06 0.89 ;
 RECT 2.235 1.02 2.375 1.24 ;
 RECT 1.78 0.59 2.165 0.73 ;
 RECT 2.025 0.73 2.165 0.88 ;
 RECT 2.025 0.88 2.375 1.02 ;
 RECT 2.235 1.38 2.375 1.95 ;
 RECT 1.78 1.95 2.375 2.09 ;
 RECT 2.735 1.205 2.965 1.24 ;
 RECT 2.235 1.24 2.965 1.38 ;
 RECT 2.735 1.38 2.965 1.415 ;
 RECT 20.915 0.36 21.055 0.79 ;
 RECT 20.115 0.36 20.255 1.41 ;
 RECT 20.05 1.41 20.32 1.55 ;
 RECT 20.115 0.22 21.055 0.36 ;
 RECT 20.915 0.79 21.535 0.93 ;
 RECT 14.46 1.095 14.6 1.835 ;
 RECT 14.785 0.925 15.015 0.955 ;
 RECT 14.46 0.955 15.015 1.095 ;
 RECT 14.785 1.095 15.015 1.135 ;
 RECT 3.475 0.6 3.88 0.735 ;
 RECT 3.475 0.735 3.615 2.13 ;
 RECT 4.755 0.41 4.895 0.46 ;
 RECT 3.475 0.595 4.895 0.6 ;
 RECT 3.68 0.46 4.895 0.595 ;
 RECT 4.755 0.275 5.655 0.41 ;
 RECT 5.515 0.41 5.655 1.475 ;
 RECT 4.755 0.27 5.59 0.275 ;
 RECT 4.755 0.6 4.895 0.61 ;
 RECT 21.675 0.435 21.815 1.07 ;
 RECT 20.875 1.07 21.815 1.21 ;
 RECT 21.675 1.21 21.815 1.64 ;
 RECT 8.22 0.24 9.02 0.38 ;
 RECT 8.88 0.38 9.02 1.305 ;
 RECT 8.22 0.38 8.36 0.93 ;
 RECT 8.88 1.445 9.02 1.66 ;
 RECT 7.655 0.93 8.36 1.07 ;
 RECT 6.325 0.375 6.465 1.26 ;
 RECT 7.655 0.375 7.795 0.93 ;
 RECT 6.155 1.26 6.465 1.4 ;
 RECT 6.155 1.4 6.295 1.77 ;
 RECT 6.325 0.235 7.795 0.375 ;
 RECT 8.88 1.305 9.6 1.445 ;
 RECT 9.46 1.26 9.6 1.305 ;
 RECT 9.46 1.445 9.6 1.51 ;
 RECT 18.15 1.33 18.29 2.52 ;
 RECT 16.045 2.52 18.29 2.66 ;
 RECT 18.8 1.33 18.94 1.925 ;
 RECT 20.59 0.64 20.73 1.925 ;
 RECT 18.15 1.19 18.94 1.33 ;
 RECT 18.8 1.925 20.73 2.065 ;
 RECT 20.525 0.5 20.775 0.64 ;
 RECT 10.3 1.775 10.44 2.52 ;
 RECT 10.07 2.52 10.44 2.66 ;
 RECT 11.42 2.135 11.56 2.435 ;
 RECT 10.86 1.775 11 2.435 ;
 RECT 10.3 1.635 11 1.775 ;
 RECT 10.86 2.435 11.56 2.575 ;
 RECT 13.515 1.86 13.655 1.995 ;
 RECT 11.42 1.995 13.655 2.135 ;
 RECT 14.175 0.75 14.315 1.72 ;
 RECT 14.175 2.045 14.84 2.185 ;
 RECT 14.175 1.86 14.315 2.045 ;
 RECT 13.515 1.72 14.315 1.86 ;
 RECT 14.175 0.61 14.86 0.75 ;
 RECT 3.77 1.13 3.91 2.42 ;
 RECT 3.105 1.975 3.25 2.155 ;
 RECT 3.105 0.48 3.245 1.975 ;
 RECT 3.11 2.155 3.25 2.42 ;
 RECT 3.11 2.42 3.91 2.56 ;
 RECT 3.77 0.99 5.055 1.13 ;
 RECT 8.78 1.94 8.92 2.05 ;
 RECT 7.02 2.05 8.92 2.19 ;
 RECT 7.02 1.805 7.16 2.05 ;
 RECT 6.805 0.545 6.945 1.665 ;
 RECT 6.735 1.665 7.16 1.805 ;
 RECT 10.3 0.365 10.44 1.205 ;
 RECT 9.74 0.365 9.88 1.8 ;
 RECT 9.74 0.225 10.44 0.365 ;
 RECT 8.78 1.8 9.88 1.94 ;
 RECT 10.3 1.205 10.925 1.345 ;
 RECT 15.095 1.845 15.235 2.45 ;
 RECT 14.06 2.385 14.2 2.45 ;
 RECT 14.06 2.45 15.235 2.59 ;
 RECT 14.06 2.59 14.2 2.65 ;
 RECT 15.95 0.55 16.09 1.705 ;
 RECT 15.095 1.705 16.09 1.845 ;
 RECT 15.95 1.845 16.09 2.265 ;
 RECT 9.06 2.23 9.2 2.33 ;
 RECT 6.69 2.33 9.2 2.47 ;
 RECT 4.555 1.945 6.83 2.085 ;
 RECT 6.69 2.085 6.83 2.33 ;
 RECT 5.825 0.835 5.965 1.945 ;
 RECT 4.56 1.715 4.7 1.945 ;
 RECT 4.49 1.575 4.765 1.715 ;
 RECT 9.06 2.09 10.16 2.23 ;
 RECT 10.02 0.52 10.16 2.09 ;
 RECT 15.255 1.17 15.595 1.51 ;
 RECT 5.195 0.55 5.335 1.275 ;
 RECT 5.195 1.415 5.335 1.71 ;
 RECT 4.05 1.275 5.335 1.415 ;
 END
END RSDFFX2

MACRO PGX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 RECT 2.01 1.855 2.15 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 RECT 2.01 0.08 2.15 0.82 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.295 2.27 1.635 2.55 ;
 END
 ANTENNAGATEAREA 0.112 ;
 END INP

 PIN INN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.3 0.26 1.6 0.63 ;
 END
 ANTENNAGATEAREA 0.035 ;
 END INN

 PIN INQ2
 DIRECTION INOUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.985 0.795 1.265 1.185 ;
 RECT 0.985 1.185 1.125 2.615 ;
 RECT 0.985 0.335 1.125 0.795 ;
 END
 ANTENNADIFFAREA 0.455 ;
 END INQ2

 PIN INQ1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.365 0.76 0.645 1.185 ;
 RECT 0.505 1.185 0.645 2.615 ;
 RECT 0.505 0.335 0.645 0.76 ;
 END
 ANTENNADIFFAREA 0.441 ;
 END INQ1

 OBS
 LAYER PO ;
 RECT 1.3 0.195 1.53 0.54 ;
 RECT 0.76 0.195 0.86 0.805 ;
 RECT 0.76 0.095 1.53 0.195 ;
 RECT 0.76 2.685 1.395 2.785 ;
 RECT 1.295 2.5 1.395 2.685 ;
 RECT 0.76 1.305 0.86 2.685 ;
 RECT 1.295 2.27 1.525 2.5 ;
 LAYER CO ;
 RECT 1.35 0.36 1.48 0.49 ;
 RECT 1.345 2.32 1.475 2.45 ;
 RECT 2.015 0.37 2.145 0.5 ;
 RECT 2.015 1.905 2.145 2.035 ;
 RECT 2.015 0.64 2.145 0.77 ;
 RECT 2.015 2.175 2.145 2.305 ;
 RECT 0.99 0.385 1.12 0.515 ;
 RECT 0.51 0.385 0.64 0.515 ;
 RECT 0.51 1.89 0.64 2.02 ;
 RECT 0.51 1.62 0.64 1.75 ;
 RECT 0.99 1.635 1.12 1.765 ;
 RECT 0.99 1.895 1.12 2.025 ;
 RECT 0.99 2.165 1.12 2.295 ;
 RECT 0.99 2.435 1.12 2.565 ;
 RECT 0.51 2.16 0.64 2.29 ;
 RECT 0.51 2.435 0.64 2.565 ;
 END
END PGX1

MACRO PGX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.88 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.88 2.96 ;
 RECT 2.33 1.855 2.47 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.88 0.08 ;
 RECT 2.33 0.08 2.47 0.825 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.625 2.235 1.965 2.66 ;
 END
 ANTENNAGATEAREA 0.224 ;
 END INP

 PIN INN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.62 0.235 1.945 0.635 ;
 END
 ANTENNAGATEAREA 0.07 ;
 END INN

 PIN INQ2
 DIRECTION INOUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.635 1.15 0.965 1.415 ;
 RECT 0.825 1.415 0.965 2.615 ;
 RECT 0.825 0.525 0.965 1.15 ;
 END
 ANTENNADIFFAREA 0.572 ;
 END INQ2

 PIN INQ1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.305 0.825 1.635 1.17 ;
 RECT 1.305 1.17 1.445 2.615 ;
 RECT 0.315 0.245 1.445 0.385 ;
 RECT 1.305 0.385 1.445 0.825 ;
 RECT 0.315 0.385 0.455 2.615 ;
 END
 ANTENNADIFFAREA 1.058 ;
 END INQ1

 OBS
 LAYER PO ;
 RECT 0.59 0.285 1.85 0.385 ;
 RECT 0.59 0.385 0.69 0.995 ;
 RECT 1.08 0.385 1.18 0.995 ;
 RECT 1.62 0.385 1.85 0.515 ;
 RECT 1.625 2.66 1.725 2.685 ;
 RECT 0.59 2.685 1.725 2.785 ;
 RECT 0.59 1.305 0.69 2.685 ;
 RECT 1.08 1.305 1.18 2.685 ;
 RECT 1.625 2.43 1.855 2.66 ;
 LAYER CO ;
 RECT 1.67 0.335 1.8 0.465 ;
 RECT 1.675 2.48 1.805 2.61 ;
 RECT 1.67 0.335 1.8 0.465 ;
 RECT 1.675 2.48 1.805 2.61 ;
 RECT 2.335 1.905 2.465 2.035 ;
 RECT 2.335 0.375 2.465 0.505 ;
 RECT 0.32 0.575 0.45 0.705 ;
 RECT 0.32 2.435 0.45 2.565 ;
 RECT 0.32 1.89 0.45 2.02 ;
 RECT 0.32 1.62 0.45 1.75 ;
 RECT 0.32 2.16 0.45 2.29 ;
 RECT 2.335 0.645 2.465 0.775 ;
 RECT 2.335 2.175 2.465 2.305 ;
 RECT 1.31 0.575 1.44 0.705 ;
 RECT 0.83 0.575 0.96 0.705 ;
 RECT 0.83 1.89 0.96 2.02 ;
 RECT 0.83 1.62 0.96 1.75 ;
 RECT 1.31 1.635 1.44 1.765 ;
 RECT 1.31 1.895 1.44 2.025 ;
 RECT 1.31 2.165 1.44 2.295 ;
 RECT 1.31 2.435 1.44 2.565 ;
 RECT 0.83 2.16 0.96 2.29 ;
 RECT 0.83 2.435 0.96 2.565 ;
 END
END PGX2

MACRO PGX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 3.025 1.855 3.165 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 3.025 0.08 3.165 0.81 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.37 2.24 2.725 2.66 ;
 END
 ANTENNAGATEAREA 0.448 ;
 END INP

 PIN INN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.365 0.29 2.885 0.695 ;
 END
 ANTENNAGATEAREA 0.14 ;
 END INN

 PIN INQ1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.59 1.15 0.92 1.42 ;
 RECT 0.59 0.525 0.73 1.15 ;
 RECT 0.59 1.42 0.73 2.515 ;
 RECT 1.57 0.525 1.71 2.515 ;
 RECT 0.585 2.515 1.71 2.655 ;
 END
 ANTENNADIFFAREA 1.116 ;
 END INQ1

 PIN INQ2
 DIRECTION INOUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.895 1.115 2.28 1.415 ;
 RECT 2.05 1.415 2.19 2.575 ;
 RECT 0.12 0.245 2.19 0.385 ;
 RECT 2.05 0.385 2.19 1.115 ;
 RECT 1.06 0.385 1.2 2.3 ;
 RECT 0.12 0.385 0.26 2.575 ;
 END
 ANTENNADIFFAREA 1.468 ;
 END INQ2

 OBS
 LAYER PO ;
 RECT 0.375 0.385 0.475 0.995 ;
 RECT 0.375 0.285 2.6 0.385 ;
 RECT 0.845 0.385 0.945 0.995 ;
 RECT 1.335 0.385 1.435 0.995 ;
 RECT 1.825 0.385 1.925 0.995 ;
 RECT 2.37 0.385 2.6 0.515 ;
 RECT 0.375 1.265 0.475 2.675 ;
 RECT 0.845 1.265 0.945 2.675 ;
 RECT 1.335 1.265 1.435 2.675 ;
 RECT 1.825 1.265 1.925 2.675 ;
 RECT 2.37 2.465 2.6 2.675 ;
 RECT 0.375 2.675 2.6 2.775 ;
 LAYER CO ;
 RECT 3.03 0.63 3.16 0.76 ;
 RECT 3.03 2.175 3.16 2.305 ;
 RECT 2.055 0.575 2.185 0.705 ;
 RECT 1.575 0.575 1.705 0.705 ;
 RECT 1.575 1.85 1.705 1.98 ;
 RECT 1.575 1.58 1.705 1.71 ;
 RECT 2.055 1.595 2.185 1.725 ;
 RECT 2.055 1.855 2.185 1.985 ;
 RECT 2.055 2.125 2.185 2.255 ;
 RECT 2.055 2.395 2.185 2.525 ;
 RECT 1.575 2.12 1.705 2.25 ;
 RECT 1.575 2.395 1.705 2.525 ;
 RECT 2.42 0.335 2.55 0.465 ;
 RECT 2.42 2.515 2.55 2.645 ;
 RECT 3.03 0.36 3.16 0.49 ;
 RECT 3.03 1.905 3.16 2.035 ;
 RECT 0.125 0.575 0.255 0.705 ;
 RECT 0.595 0.575 0.725 0.705 ;
 RECT 0.125 2.12 0.255 2.25 ;
 RECT 0.125 2.395 0.255 2.525 ;
 RECT 0.125 1.85 0.255 1.98 ;
 RECT 0.125 1.58 0.255 1.71 ;
 RECT 0.595 2.12 0.725 2.25 ;
 RECT 0.595 2.395 0.725 2.525 ;
 RECT 0.595 1.85 0.725 1.98 ;
 RECT 0.595 1.58 0.725 1.71 ;
 RECT 1.065 0.575 1.195 0.705 ;
 RECT 1.065 1.85 1.195 1.98 ;
 RECT 1.065 1.58 1.195 1.71 ;
 RECT 1.065 2.12 1.195 2.25 ;
 END
END PGX4

MACRO RDFFNX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 19.84 BY 2.88 ;
 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.085 1.145 6.395 1.415 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.32 1.5 8.46 2.295 ;
 RECT 8.32 1.09 8.74 1.5 ;
 RECT 8.32 0.525 8.46 1.09 ;
 END
 ANTENNADIFFAREA 0.504 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.37 1.295 9.51 1.79 ;
 RECT 9.37 0.97 9.755 1.295 ;
 RECT 9.37 0.48 9.51 0.97 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 19.84 2.96 ;
 RECT 4.67 2.615 4.905 2.8 ;
 RECT 6.135 2.37 6.405 2.51 ;
 RECT 2.715 2.51 2.945 2.65 ;
 RECT 1.02 2.51 1.29 2.65 ;
 RECT 8.89 2.275 9.03 2.8 ;
 RECT 7.375 1.94 7.515 2.8 ;
 RECT 0.205 1.64 0.365 2.8 ;
 RECT 9.93 2 10.07 2.8 ;
 RECT 11.62 2.025 11.76 2.8 ;
 RECT 6.2 2.51 6.34 2.8 ;
 RECT 2.76 2.65 2.9 2.8 ;
 RECT 1.085 2.65 1.225 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 19.84 0.08 ;
 RECT 2.725 0.555 2.975 0.695 ;
 RECT 6.125 0.565 6.395 0.705 ;
 RECT 14.58 0.22 14.83 0.36 ;
 RECT 8.89 0.08 9.03 0.575 ;
 RECT 0.205 0.08 0.365 0.84 ;
 RECT 9.98 0.08 10.12 0.865 ;
 RECT 11.62 0.08 11.76 0.815 ;
 RECT 7.375 0.08 7.515 0.785 ;
 RECT 4.735 0.08 4.875 0.78 ;
 RECT 17.345 0.08 17.485 0.65 ;
 RECT 1.085 0.08 1.225 0.32 ;
 RECT 2.79 0.08 2.93 0.555 ;
 RECT 6.19 0.08 6.33 0.565 ;
 RECT 14.625 0.08 14.765 0.22 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 18.2 1.4 18.54 1.765 ;
 RECT 14.625 2.225 18.355 2.385 ;
 RECT 14.58 1.47 14.81 1.61 ;
 RECT 17.3 1.395 17.44 2.225 ;
 RECT 18.215 1.765 18.355 2.225 ;
 RECT 14.625 1.61 14.765 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.75 0.81 13.13 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.45 0.825 1.85 1.135 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 8.575 1.32 8.675 2.75 ;
 RECT 7.47 1.22 8.675 1.32 ;
 RECT 11.405 1.215 11.68 1.27 ;
 RECT 11.405 1.37 11.68 1.425 ;
 RECT 11.405 1.27 11.98 1.37 ;
 RECT 11.88 1.045 11.98 1.27 ;
 RECT 11.88 1.37 11.98 2.425 ;
 RECT 14.33 1.045 14.43 1.76 ;
 RECT 11.405 0.385 11.505 1.215 ;
 RECT 11.405 1.425 11.505 2.425 ;
 RECT 12.84 0.84 13.07 0.945 ;
 RECT 12.84 1.045 13.07 1.07 ;
 RECT 11.88 0.385 11.98 0.945 ;
 RECT 11.88 0.945 14.43 1.045 ;
 RECT 14.33 0.145 14.43 0.945 ;
 RECT 15.485 1.86 15.585 2.09 ;
 RECT 15.355 1.545 15.585 1.76 ;
 RECT 16.52 1.145 16.62 2.09 ;
 RECT 14.33 1.76 15.585 1.86 ;
 RECT 15.485 2.09 16.62 2.19 ;
 RECT 5.015 0.37 5.115 2.68 ;
 RECT 6.885 2.475 7.115 2.68 ;
 RECT 5.015 2.68 7.115 2.78 ;
 RECT 6.47 0.33 6.57 1.175 ;
 RECT 6.47 1.395 6.57 2.235 ;
 RECT 6.21 1.175 6.57 1.395 ;
 RECT 10.265 0.385 10.365 2.405 ;
 RECT 10.165 2.405 10.395 2.635 ;
 RECT 3.86 1.445 3.96 2.285 ;
 RECT 3.775 2.285 4.005 2.515 ;
 RECT 10.575 1.835 10.675 2.425 ;
 RECT 10.565 1.605 10.795 1.835 ;
 RECT 2.265 1.34 2.495 1.45 ;
 RECT 2.265 0.38 2.365 1.24 ;
 RECT 2.265 1.45 2.365 2.345 ;
 RECT 3.36 0.38 3.46 1.24 ;
 RECT 2.265 1.24 3.46 1.34 ;
 RECT 3.36 1.34 3.46 2.58 ;
 RECT 1.34 0.1 4.035 0.2 ;
 RECT 3.735 0.2 4.035 0.42 ;
 RECT 1.34 0.2 1.44 0.97 ;
 RECT 3.935 0.42 4.035 0.95 ;
 RECT 5.93 0.33 6.03 2.135 ;
 RECT 5.81 2.135 6.04 2.365 ;
 RECT 1.74 0.38 1.84 0.945 ;
 RECT 1.74 1.175 1.84 2.36 ;
 RECT 1.62 0.945 1.85 1.175 ;
 RECT 2.57 0.87 3.145 0.97 ;
 RECT 3.045 0.38 3.145 0.87 ;
 RECT 2.57 0.84 2.815 0.87 ;
 RECT 2.57 0.97 2.815 1.06 ;
 RECT 2.57 0.38 2.67 0.84 ;
 RECT 1.43 1.76 1.53 2.34 ;
 RECT 1.31 1.53 1.54 1.76 ;
 RECT 0.88 0.38 0.98 1.23 ;
 RECT 0.88 1.46 0.98 2.34 ;
 RECT 0.88 1.23 1.115 1.46 ;
 RECT 4.465 0.37 4.565 1.21 ;
 RECT 4.465 1.21 4.75 1.42 ;
 RECT 4.465 1.42 4.565 2.16 ;
 RECT 3.035 1.75 3.135 2.585 ;
 RECT 2.905 1.53 3.135 1.63 ;
 RECT 2.905 1.73 3.135 1.75 ;
 RECT 2.565 1.73 2.665 2.34 ;
 RECT 2.565 1.63 3.135 1.73 ;
 RECT 16.995 0.275 17.095 1.025 ;
 RECT 16.995 1.255 17.095 1.86 ;
 RECT 16.995 1.025 17.275 1.255 ;
 RECT 15.335 0.865 16.06 0.965 ;
 RECT 15.335 0.735 15.565 0.865 ;
 RECT 15.96 0.275 16.06 0.865 ;
 RECT 9.155 0.105 12.53 0.205 ;
 RECT 9.155 0.205 9.255 0.87 ;
 RECT 11.06 0.205 11.16 0.925 ;
 RECT 12.3 0.205 12.53 0.4 ;
 RECT 9.155 1.085 9.255 2.755 ;
 RECT 9.01 0.87 9.255 1.085 ;
 RECT 10.935 0.925 11.165 1.135 ;
 RECT 14.91 0.965 15.01 1.145 ;
 RECT 16.52 0.275 16.62 0.865 ;
 RECT 16.24 0.965 16.34 1.145 ;
 RECT 14.91 1.145 16.34 1.245 ;
 RECT 16.05 1.245 16.15 1.86 ;
 RECT 14.91 0.735 15.14 0.965 ;
 RECT 16.24 0.865 16.62 0.965 ;
 RECT 11.105 2.605 12.455 2.695 ;
 RECT 11.11 2.695 12.455 2.705 ;
 RECT 11.105 1.425 11.205 2.605 ;
 RECT 10.57 0.385 10.67 1.325 ;
 RECT 10.57 1.325 11.205 1.425 ;
 RECT 12.225 2.475 12.455 2.605 ;
 RECT 17.6 0.27 17.7 0.745 ;
 RECT 17.6 0.975 17.7 1.855 ;
 RECT 17.455 0.745 17.7 0.975 ;
 RECT 7.665 0.365 7.765 1.16 ;
 RECT 7.47 1.16 7.765 1.22 ;
 RECT 7.665 1.39 7.765 2.47 ;
 RECT 7.47 1.32 7.765 1.39 ;
 RECT 8.575 0.105 8.675 1.22 ;
 LAYER CO ;
 RECT 12.105 2.065 12.235 2.195 ;
 RECT 8.325 1.715 8.455 1.845 ;
 RECT 3.825 2.335 3.955 2.465 ;
 RECT 6.935 2.525 7.065 2.655 ;
 RECT 2.955 1.57 3.085 1.7 ;
 RECT 9.06 0.915 9.19 1.045 ;
 RECT 2.315 1.28 2.445 1.41 ;
 RECT 1.36 1.58 1.49 1.71 ;
 RECT 1.67 0.995 1.8 1.125 ;
 RECT 0.935 1.28 1.065 1.41 ;
 RECT 6.82 0.57 6.95 0.7 ;
 RECT 6.82 1.87 6.95 2 ;
 RECT 6.195 0.57 6.325 0.7 ;
 RECT 5.68 0.57 5.81 0.7 ;
 RECT 5.68 1.48 5.81 1.61 ;
 RECT 6.205 2.375 6.335 2.505 ;
 RECT 4.725 2.63 4.855 2.76 ;
 RECT 0.62 1.935 0.75 2.065 ;
 RECT 0.62 0.6 0.75 0.73 ;
 RECT 3.605 1.67 3.735 1.8 ;
 RECT 1.09 2.515 1.22 2.645 ;
 RECT 2.765 2.515 2.895 2.645 ;
 RECT 1.995 1.52 2.125 1.65 ;
 RECT 5.3 1.705 5.43 1.835 ;
 RECT 5.3 0.6 5.43 0.73 ;
 RECT 4.74 0.6 4.87 0.73 ;
 RECT 4.165 0.6 4.295 0.73 ;
 RECT 4.165 1.48 4.295 1.61 ;
 RECT 3.605 0.6 3.735 0.73 ;
 RECT 2.795 0.555 2.925 0.685 ;
 RECT 1.995 0.6 2.125 0.73 ;
 RECT 12.35 0.225 12.48 0.355 ;
 RECT 14.63 1.475 14.76 1.605 ;
 RECT 14.025 1.255 14.155 1.385 ;
 RECT 13.98 0.505 14.11 0.635 ;
 RECT 12.275 2.525 12.405 2.655 ;
 RECT 10.215 2.455 10.345 2.585 ;
 RECT 10.615 1.655 10.745 1.785 ;
 RECT 12.105 0.635 12.235 0.765 ;
 RECT 11.625 0.635 11.755 0.765 ;
 RECT 11.625 2.075 11.755 2.205 ;
 RECT 15.385 0.785 15.515 0.915 ;
 RECT 17.83 0.505 17.96 0.635 ;
 RECT 17.83 1.44 17.96 1.57 ;
 RECT 16.745 1.435 16.875 1.565 ;
 RECT 16.745 0.505 16.875 0.635 ;
 RECT 8.895 0.395 9.025 0.525 ;
 RECT 8.325 0.585 8.455 0.715 ;
 RECT 11.5 1.255 11.63 1.385 ;
 RECT 10.985 0.965 11.115 1.095 ;
 RECT 6.26 1.215 6.39 1.345 ;
 RECT 3.785 0.24 3.915 0.37 ;
 RECT 2.625 0.89 2.755 1.02 ;
 RECT 4.57 1.25 4.7 1.38 ;
 RECT 17.505 0.795 17.635 0.925 ;
 RECT 17.095 1.075 17.225 1.205 ;
 RECT 17.35 0.47 17.48 0.6 ;
 RECT 17.305 1.455 17.435 1.585 ;
 RECT 9.375 1.6 9.505 1.73 ;
 RECT 8.325 2.105 8.455 2.235 ;
 RECT 8.895 2.34 9.025 2.47 ;
 RECT 5.86 2.185 5.99 2.315 ;
 RECT 12.89 0.89 13.02 1.02 ;
 RECT 15.405 1.595 15.535 1.725 ;
 RECT 14.96 0.785 15.09 0.915 ;
 RECT 1.09 0.12 1.22 0.25 ;
 RECT 18.25 1.44 18.38 1.57 ;
 RECT 0.22 0.36 0.35 0.49 ;
 RECT 0.22 0.62 0.35 0.75 ;
 RECT 0.22 1.71 0.35 1.84 ;
 RECT 0.22 1.97 0.35 2.1 ;
 RECT 0.22 2.23 0.35 2.36 ;
 RECT 14.63 0.225 14.76 0.355 ;
 RECT 16.27 1.415 16.4 1.545 ;
 RECT 16.27 0.505 16.4 0.635 ;
 RECT 15.71 1.415 15.84 1.545 ;
 RECT 15.71 0.505 15.84 0.635 ;
 RECT 9.375 0.555 9.505 0.685 ;
 RECT 7.38 2.01 7.51 2.14 ;
 RECT 7.52 1.21 7.65 1.34 ;
 RECT 7.38 0.605 7.51 0.735 ;
 RECT 7.94 2.025 8.07 2.155 ;
 RECT 7.94 0.605 8.07 0.735 ;
 RECT 10.81 2.05 10.94 2.18 ;
 RECT 10.81 0.635 10.94 0.765 ;
 RECT 9.985 0.635 10.115 0.765 ;
 RECT 9.935 2.06 10.065 2.19 ;
 LAYER M1 ;
 RECT 0.93 1.21 1.07 1.275 ;
 RECT 0.93 1.415 1.07 1.48 ;
 RECT 1.99 0.55 2.13 1.275 ;
 RECT 1.99 1.415 2.13 1.71 ;
 RECT 0.93 1.275 2.13 1.415 ;
 RECT 11.405 1.17 11.745 1.51 ;
 RECT 15.4 0.92 15.54 1.785 ;
 RECT 15.315 0.78 15.565 0.92 ;
 RECT 10.61 1.095 10.75 1.835 ;
 RECT 10.935 0.925 11.165 0.955 ;
 RECT 10.61 0.955 11.165 1.095 ;
 RECT 10.935 1.095 11.165 1.135 ;
 RECT 11.245 1.845 11.385 2.45 ;
 RECT 10.21 2.385 10.35 2.45 ;
 RECT 10.21 2.45 11.385 2.59 ;
 RECT 10.21 2.59 10.35 2.65 ;
 RECT 12.1 0.585 12.24 1.705 ;
 RECT 12.1 1.845 12.24 2.265 ;
 RECT 11.245 1.705 12.24 1.845 ;
 RECT 4.16 0.55 4.3 1.475 ;
 RECT 4.095 1.475 4.365 1.615 ;
 RECT 14.3 0.36 14.44 0.5 ;
 RECT 12.25 0.22 14.44 0.36 ;
 RECT 15.705 0.435 15.845 0.5 ;
 RECT 15.705 0.64 15.845 1.61 ;
 RECT 14.3 0.5 15.845 0.64 ;
 RECT 14.02 0.64 14.16 0.78 ;
 RECT 14.02 0.92 14.16 1.455 ;
 RECT 13.915 0.5 14.16 0.64 ;
 RECT 14.02 0.78 15.155 0.92 ;
 RECT 17.825 0.435 17.965 1.07 ;
 RECT 17.825 1.21 17.965 1.64 ;
 RECT 17.025 1.07 17.965 1.21 ;
 RECT 0.615 0.6 0.755 2.13 ;
 RECT 1.55 0.41 1.69 0.46 ;
 RECT 0.615 0.46 1.69 0.6 ;
 RECT 2.31 0.41 2.45 1.475 ;
 RECT 1.55 0.27 2.45 0.41 ;
 RECT 7.935 0.385 8.075 2.21 ;
 RECT 8.6 0.385 8.74 0.75 ;
 RECT 7.935 0.245 8.74 0.385 ;
 RECT 9.055 0.89 9.195 1.095 ;
 RECT 8.6 0.75 9.195 0.89 ;
 RECT 7.655 1.775 7.795 2.435 ;
 RECT 7.095 1.635 7.795 1.775 ;
 RECT 7.095 1.775 7.235 2.52 ;
 RECT 6.865 2.52 7.235 2.66 ;
 RECT 9.65 1.86 9.79 1.995 ;
 RECT 8.61 1.995 9.79 2.135 ;
 RECT 8.61 2.135 8.75 2.435 ;
 RECT 7.655 2.435 8.75 2.575 ;
 RECT 10.325 2.045 10.99 2.185 ;
 RECT 10.325 1.86 10.465 2.045 ;
 RECT 10.325 0.63 10.99 0.77 ;
 RECT 10.325 0.77 10.465 1.72 ;
 RECT 9.65 1.72 10.465 1.86 ;
 RECT 3.485 2.33 5.995 2.47 ;
 RECT 5.855 2.23 5.995 2.33 ;
 RECT 3.485 2.085 3.625 2.33 ;
 RECT 1.355 1.945 3.625 2.085 ;
 RECT 2.62 0.835 2.76 1.945 ;
 RECT 1.355 1.715 1.495 1.945 ;
 RECT 1.285 1.575 1.56 1.715 ;
 RECT 5.855 2.09 6.955 2.23 ;
 RECT 6.815 0.52 6.955 2.09 ;
 RECT 3.12 0.375 3.26 1.26 ;
 RECT 4.45 0.375 4.59 0.93 ;
 RECT 2.95 1.26 3.26 1.4 ;
 RECT 2.95 1.4 3.09 1.77 ;
 RECT 3.12 0.235 4.59 0.375 ;
 RECT 5.015 0.24 5.815 0.38 ;
 RECT 5.675 0.38 5.815 1.66 ;
 RECT 5.015 0.38 5.155 0.93 ;
 RECT 4.45 0.93 5.155 1.07 ;
 RECT 17.065 0.36 17.205 0.79 ;
 RECT 16.265 0.36 16.405 1.41 ;
 RECT 16.2 1.41 16.47 1.55 ;
 RECT 16.265 0.22 17.205 0.36 ;
 RECT 17.065 0.79 17.685 0.93 ;
 RECT 5.575 1.94 5.715 2.05 ;
 RECT 3.815 2.05 5.715 2.19 ;
 RECT 3.815 1.805 3.955 2.05 ;
 RECT 3.6 0.545 3.74 1.665 ;
 RECT 3.53 1.665 3.955 1.805 ;
 RECT 7.095 0.365 7.235 1.205 ;
 RECT 6.535 0.365 6.675 1.8 ;
 RECT 6.535 0.225 7.235 0.365 ;
 RECT 5.575 1.8 6.675 1.94 ;
 RECT 7.095 1.205 7.72 1.345 ;
 RECT 5.295 0.55 5.435 1.245 ;
 RECT 5.295 1.385 5.435 1.9 ;
 RECT 4.52 1.245 5.435 1.385 ;
 RECT 4.52 1.21 4.75 1.245 ;
 RECT 4.52 1.385 4.75 1.42 ;
 RECT 14.3 1.33 14.44 2.52 ;
 RECT 12.195 2.52 14.44 2.66 ;
 RECT 14.95 1.33 15.09 1.925 ;
 RECT 16.74 0.64 16.88 1.925 ;
 RECT 14.3 1.19 15.09 1.33 ;
 RECT 14.95 1.925 16.88 2.065 ;
 RECT 16.675 0.5 16.925 0.64 ;
 END
END RDFFNX1

MACRO RDFFNSRASX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.84 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.895 0.59 21.265 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.125 1.435 26.465 1.8 ;
 RECT 24.445 1.99 26.31 2.13 ;
 RECT 22.215 2.22 24.585 2.36 ;
 RECT 26.17 1.8 26.31 1.99 ;
 RECT 24.445 1.435 24.585 1.99 ;
 RECT 22.215 1.39 22.355 2.22 ;
 RECT 23.6 1.37 23.74 2.22 ;
 RECT 24.445 2.13 24.585 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.84 2.12 1.16 2.585 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.825 0.08 2.105 0.295 ;
 RECT 24.565 0.08 24.805 0.26 ;
 RECT 5.755 0.31 6.045 0.45 ;
 RECT 9.44 0.615 9.71 0.755 ;
 RECT 13.365 0.275 14.39 0.415 ;
 RECT 17.725 0.335 17.99 0.495 ;
 RECT 14.25 0.75 15.195 0.89 ;
 RECT 0 -0.08 27.84 0.08 ;
 RECT 0.335 0.08 0.475 0.775 ;
 RECT 1.305 0.08 1.445 0.97 ;
 RECT 4.65 0.08 4.885 0.46 ;
 RECT 19.37 0.08 19.51 0.82 ;
 RECT 22.215 0.08 22.355 0.36 ;
 RECT 23.43 0.08 23.57 0.35 ;
 RECT 5.835 0.08 5.975 0.31 ;
 RECT 9.505 0.08 9.645 0.615 ;
 RECT 13.365 0.415 13.505 0.945 ;
 RECT 13.365 0.08 13.505 0.275 ;
 RECT 17.78 0.08 17.92 0.335 ;
 RECT 15.055 0.89 15.195 1.11 ;
 RECT 14.25 0.415 14.39 0.75 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.18 1.205 17.43 1.445 ;
 RECT 17.29 0.915 17.43 1.205 ;
 RECT 18.295 1.84 18.435 1.885 ;
 RECT 18.295 0.915 18.435 1.7 ;
 RECT 17.29 1.84 17.43 1.885 ;
 RECT 17.29 1.7 18.435 1.84 ;
 RECT 17.29 1.445 17.43 1.7 ;
 END
 ANTENNADIFFAREA 0.7 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 17.635 2.6 17.9 2.8 ;
 RECT 19.225 2.6 19.49 2.8 ;
 RECT 9.25 2.215 9.525 2.355 ;
 RECT 0 2.8 27.84 2.96 ;
 RECT 0.335 1.74 0.475 2.8 ;
 RECT 1.98 2.34 2.23 2.8 ;
 RECT 1.305 1.98 1.445 2.8 ;
 RECT 5.835 1.98 5.975 2.8 ;
 RECT 6.865 2 7.005 2.8 ;
 RECT 12.275 2.335 12.545 2.8 ;
 RECT 5.355 2.615 5.495 2.8 ;
 RECT 5.355 2.405 5.685 2.615 ;
 RECT 5.355 2.07 5.495 2.405 ;
 RECT 9.315 2.355 9.455 2.8 ;
 RECT 9.315 2.195 9.455 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 1.475 1.685 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.69 1.095 18.95 1.335 ;
 RECT 18.81 0.51 18.95 1.095 ;
 RECT 19.87 1.905 20.01 1.91 ;
 RECT 18.81 1.765 20.01 1.905 ;
 RECT 19.87 0.56 20.01 1.765 ;
 RECT 18.81 1.905 18.95 1.915 ;
 RECT 18.81 1.335 18.95 1.765 ;
 END
 ANTENNADIFFAREA 0.568 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.73 2.255 10.04 2.465 ;
 RECT 9.8 2.465 10.04 2.47 ;
 RECT 9.8 2.12 10.04 2.255 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.24 1.795 7.48 2.04 ;
 RECT 6.655 1.795 6.885 1.83 ;
 RECT 6.655 1.655 7.48 1.795 ;
 RECT 6.655 1.62 6.885 1.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 OBS
 LAYER PO ;
 RECT 2.405 0.195 4.56 0.285 ;
 RECT 11.195 0.195 11.295 1.29 ;
 RECT 12.09 1.39 12.285 1.405 ;
 RECT 3.225 1.565 3.325 2.675 ;
 RECT 2.34 1.62 2.44 2.675 ;
 RECT 1.905 1.44 2.15 1.52 ;
 RECT 1.905 1.62 2.15 1.69 ;
 RECT 4.46 0.285 4.56 1.24 ;
 RECT 11.195 1.29 12.285 1.39 ;
 RECT 2.34 2.675 3.325 2.775 ;
 RECT 12.09 1.405 12.32 1.615 ;
 RECT 22.475 1.245 22.575 2.02 ;
 RECT 22.345 1.035 22.575 1.245 ;
 RECT 12.585 0.105 15.41 0.205 ;
 RECT 12.585 0.205 12.685 1.91 ;
 RECT 15.31 0.205 15.41 1.265 ;
 RECT 11.765 1.71 11.865 1.91 ;
 RECT 10.68 1.61 11.865 1.71 ;
 RECT 10.68 0.475 10.78 1.61 ;
 RECT 11.23 1.71 11.33 2.425 ;
 RECT 7.345 0.475 7.445 0.895 ;
 RECT 11.765 1.91 12.685 2.01 ;
 RECT 7.345 0.375 10.78 0.475 ;
 RECT 7.22 0.895 7.45 1.105 ;
 RECT 12.895 0.455 14.825 0.535 ;
 RECT 14.595 0.535 14.825 0.6 ;
 RECT 14.595 0.39 14.825 0.435 ;
 RECT 12.975 0.435 14.825 0.455 ;
 RECT 12.895 0.535 13.125 0.665 ;
 RECT 13.75 0.535 13.98 0.835 ;
 RECT 13.75 0.835 13.85 2.39 ;
 RECT 22.78 0.215 22.88 0.995 ;
 RECT 22.78 0.995 23.02 1.205 ;
 RECT 22.78 1.205 22.88 2 ;
 RECT 25.175 0.375 25.275 0.99 ;
 RECT 25.175 0.99 25.425 1.2 ;
 RECT 25.175 1.2 25.275 2.27 ;
 RECT 25.175 2.27 25.46 2.48 ;
 RECT 10.16 0.655 10.26 2.305 ;
 RECT 10.465 2.3 10.695 2.305 ;
 RECT 10.465 2.405 10.695 2.51 ;
 RECT 10.16 2.305 10.695 2.405 ;
 RECT 22 0.21 22.1 0.755 ;
 RECT 22 0.855 22.1 2.2 ;
 RECT 24.865 1.125 24.965 2.2 ;
 RECT 21.035 0.755 22.57 0.84 ;
 RECT 21.035 0.84 22.565 0.855 ;
 RECT 22.47 0.215 22.57 0.755 ;
 RECT 21.035 0.595 21.265 0.755 ;
 RECT 22 2.2 24.965 2.3 ;
 RECT 23.69 0.38 23.79 0.96 ;
 RECT 23.69 1.06 23.79 1.14 ;
 RECT 23.27 0.935 23.5 0.96 ;
 RECT 23.27 0.96 23.79 1.06 ;
 RECT 23.27 1.06 23.5 1.145 ;
 RECT 23.69 1.14 23.96 1.24 ;
 RECT 23.86 1.24 23.96 1.84 ;
 RECT 24.055 0.22 24.285 0.28 ;
 RECT 24.055 0.38 24.285 0.43 ;
 RECT 23.69 0.28 24.285 0.38 ;
 RECT 7.945 1.575 8.045 2.485 ;
 RECT 8.455 1.575 8.685 1.685 ;
 RECT 7.945 1.475 8.685 1.575 ;
 RECT 25.875 0.195 25.975 2.665 ;
 RECT 24.865 0.095 25.975 0.195 ;
 RECT 21.24 1.245 21.34 2.665 ;
 RECT 24.865 0.195 24.965 0.945 ;
 RECT 21.24 1.2 21.525 1.245 ;
 RECT 21.295 1.035 21.525 1.1 ;
 RECT 21.24 2.665 25.975 2.765 ;
 RECT 21.24 1.1 21.57 1.2 ;
 RECT 12.17 0.795 12.335 0.925 ;
 RECT 11.49 0.885 11.72 0.925 ;
 RECT 11.49 1.025 11.72 1.095 ;
 RECT 11.49 0.925 12.335 1.025 ;
 RECT 12.17 0.585 12.4 0.795 ;
 RECT 3.27 0.705 3.37 1.165 ;
 RECT 2.83 1.27 2.93 1.445 ;
 RECT 3.27 0.47 3.555 0.705 ;
 RECT 2.83 1.17 3.37 1.265 ;
 RECT 2.83 1.265 3.205 1.27 ;
 RECT 3.06 1.165 3.37 1.17 ;
 RECT 2.685 1.445 2.93 1.69 ;
 RECT 4.16 0.715 4.26 1.61 ;
 RECT 4.195 1.71 4.295 2.48 ;
 RECT 4.16 1.61 4.295 1.71 ;
 RECT 4.04 0.485 4.28 0.715 ;
 RECT 9.765 0.655 9.865 1.205 ;
 RECT 9.16 1.305 9.39 1.475 ;
 RECT 9.16 1.205 9.865 1.305 ;
 RECT 1.565 0.49 1.665 1.495 ;
 RECT 1.37 1.495 1.665 1.745 ;
 RECT 1.565 1.745 1.665 2.37 ;
 RECT 3.72 1.33 3.86 1.475 ;
 RECT 3.72 1.71 3.82 2.475 ;
 RECT 3.76 0.65 3.86 1.33 ;
 RECT 3.72 1.475 3.95 1.71 ;
 RECT 0.92 2.365 1.19 2.575 ;
 RECT 1.09 0.425 1.19 2.365 ;
 RECT 8.87 0.655 8.97 1.18 ;
 RECT 8.87 1.28 8.97 1.655 ;
 RECT 7.955 0.66 8.055 1.18 ;
 RECT 8.87 1.655 9.83 1.755 ;
 RECT 9.73 1.755 9.83 2.255 ;
 RECT 8.87 1.755 8.97 2.51 ;
 RECT 7.955 1.18 8.97 1.28 ;
 RECT 9.73 2.255 9.96 2.465 ;
 RECT 5.39 0.54 5.715 0.71 ;
 RECT 5.615 0.71 5.715 2.405 ;
 RECT 5.455 2.405 5.715 2.61 ;
 RECT 5.455 2.61 5.685 2.615 ;
 RECT 5.39 0.5 5.62 0.54 ;
 RECT 16.19 0.77 16.29 2.155 ;
 RECT 16.19 0.55 16.29 0.56 ;
 RECT 16.19 0.56 16.445 0.77 ;
 RECT 16.825 0.43 16.925 1.245 ;
 RECT 17.555 0.39 17.655 1.4 ;
 RECT 17.555 1.5 17.655 2.37 ;
 RECT 18.045 0.51 18.145 1.4 ;
 RECT 18.045 1.5 18.145 2.37 ;
 RECT 16.76 0.22 16.99 0.29 ;
 RECT 16.76 0.39 16.99 0.43 ;
 RECT 16.76 0.29 17.655 0.39 ;
 RECT 17.555 1.4 18.145 1.5 ;
 RECT 16.775 1.245 17.005 1.455 ;
 RECT 4.98 2.445 5.24 2.655 ;
 RECT 5.14 1.79 5.24 2.445 ;
 RECT 15.25 1.445 15.35 2.035 ;
 RECT 15.235 2.035 15.465 2.245 ;
 RECT 15.72 0.55 15.82 2.69 ;
 RECT 6.65 1.58 6.75 1.62 ;
 RECT 6.39 1.01 6.49 1.48 ;
 RECT 6.65 1.83 6.75 2.69 ;
 RECT 6.65 1.62 6.885 1.83 ;
 RECT 6.39 1.48 6.75 1.58 ;
 RECT 6.65 2.69 15.82 2.79 ;
 RECT 6.09 0.98 6.19 1.615 ;
 RECT 5.95 1.615 6.19 1.825 ;
 RECT 6.09 1.825 6.19 2.51 ;
 RECT 19.07 1.25 19.32 1.33 ;
 RECT 19.07 1.33 19.75 1.43 ;
 RECT 19.07 1.43 19.32 1.46 ;
 RECT 19.65 0.365 19.75 1.33 ;
 RECT 19.07 0.385 19.17 1.25 ;
 RECT 19.07 1.46 19.17 2.575 ;
 RECT 19.65 1.43 19.75 2.575 ;
 RECT 20.255 0.22 20.485 0.265 ;
 RECT 20.255 0.365 20.485 0.43 ;
 RECT 19.65 0.265 20.485 0.365 ;
 RECT 14.22 0.73 14.32 1.39 ;
 RECT 14.085 1.39 14.32 1.6 ;
 RECT 14.22 1.6 14.32 2.39 ;
 RECT 2.405 0.285 2.505 1.52 ;
 RECT 1.905 1.52 2.505 1.62 ;
 RECT 2.405 0.185 11.295 0.195 ;
 RECT 4.46 0.095 11.295 0.185 ;
 LAYER CO ;
 RECT 6.87 2.11 7 2.24 ;
 RECT 19.375 0.62 19.505 0.75 ;
 RECT 5.36 2.135 5.49 2.265 ;
 RECT 2.975 2.105 3.105 2.235 ;
 RECT 3.94 2.11 4.07 2.24 ;
 RECT 1.895 0.145 2.025 0.275 ;
 RECT 10.945 1.9 11.075 2.03 ;
 RECT 0.34 2.345 0.47 2.475 ;
 RECT 2.05 2.345 2.18 2.475 ;
 RECT 23 0.435 23.13 0.565 ;
 RECT 17.295 1.705 17.425 1.835 ;
 RECT 6.65 1.23 6.78 1.36 ;
 RECT 15.47 1.705 15.6 1.835 ;
 RECT 5.84 2.075 5.97 2.205 ;
 RECT 3.49 0.88 3.62 1.01 ;
 RECT 13.5 1.835 13.63 1.965 ;
 RECT 0.97 2.405 1.1 2.535 ;
 RECT 9.78 2.295 9.91 2.425 ;
 RECT 5.505 2.445 5.635 2.575 ;
 RECT 5.44 0.54 5.57 0.67 ;
 RECT 19.14 1.29 19.27 1.42 ;
 RECT 16.825 1.285 16.955 1.415 ;
 RECT 14.645 0.43 14.775 0.56 ;
 RECT 16.265 0.6 16.395 0.73 ;
 RECT 16.81 0.26 16.94 0.39 ;
 RECT 5.03 2.485 5.16 2.615 ;
 RECT 15.285 2.075 15.415 2.205 ;
 RECT 6.705 1.66 6.835 1.79 ;
 RECT 6 1.655 6.13 1.785 ;
 RECT 20.305 0.26 20.435 0.39 ;
 RECT 25.245 1.03 25.375 1.16 ;
 RECT 12.945 0.495 13.075 0.625 ;
 RECT 14.135 1.43 14.265 1.56 ;
 RECT 12.22 0.625 12.35 0.755 ;
 RECT 12.14 1.445 12.27 1.575 ;
 RECT 22.395 1.075 22.525 1.205 ;
 RECT 7.27 0.935 7.4 1.065 ;
 RECT 23.32 0.975 23.45 1.105 ;
 RECT 13.8 0.665 13.93 0.795 ;
 RECT 22.84 1.035 22.97 1.165 ;
 RECT 25.28 2.31 25.41 2.44 ;
 RECT 10.515 2.34 10.645 2.47 ;
 RECT 21.085 0.635 21.215 0.765 ;
 RECT 24.105 0.26 24.235 0.39 ;
 RECT 8.505 1.515 8.635 1.645 ;
 RECT 21.345 1.075 21.475 1.205 ;
 RECT 11.54 0.925 11.67 1.055 ;
 RECT 3.02 0.88 3.15 1.01 ;
 RECT 11.45 1.87 11.58 2 ;
 RECT 4.89 2.11 5.02 2.24 ;
 RECT 4.705 0.32 4.835 0.45 ;
 RECT 22.22 0.135 22.35 0.265 ;
 RECT 1.965 1.495 2.095 1.625 ;
 RECT 1.915 0.745 2.045 0.875 ;
 RECT 1.785 1.995 1.915 2.125 ;
 RECT 8.62 1.995 8.75 2.125 ;
 RECT 0.34 0.59 0.47 0.72 ;
 RECT 8.175 2.07 8.305 2.2 ;
 RECT 10.945 0.595 11.075 0.725 ;
 RECT 2.74 1.49 2.87 1.62 ;
 RECT 9.21 1.28 9.34 1.41 ;
 RECT 18.815 1.725 18.945 1.855 ;
 RECT 0.34 2.085 0.47 2.215 ;
 RECT 6.38 2.045 6.51 2.175 ;
 RECT 1.43 1.55 1.56 1.68 ;
 RECT 13.37 0.765 13.5 0.895 ;
 RECT 1.31 0.74 1.44 0.87 ;
 RECT 24.615 0.12 24.745 0.25 ;
 RECT 4.095 0.53 4.225 0.66 ;
 RECT 18.815 0.62 18.945 0.75 ;
 RECT 12.345 2.38 12.475 2.51 ;
 RECT 8.62 0.905 8.75 1.035 ;
 RECT 21.75 1.425 21.88 1.555 ;
 RECT 0.34 0.33 0.47 0.46 ;
 RECT 16.535 0.92 16.665 1.05 ;
 RECT 22.22 1.475 22.35 1.605 ;
 RECT 10.42 0.875 10.55 1.005 ;
 RECT 2.625 0.79 2.755 0.92 ;
 RECT 14.44 1.835 14.57 1.965 ;
 RECT 3.47 2.07 3.6 2.2 ;
 RECT 26.175 1.475 26.305 1.605 ;
 RECT 18.3 1.705 18.43 1.835 ;
 RECT 19.875 1.71 20.005 1.84 ;
 RECT 17.295 0.975 17.425 1.105 ;
 RECT 0.84 0.74 0.97 0.87 ;
 RECT 2.56 1.825 2.69 1.955 ;
 RECT 10.42 1.945 10.55 2.075 ;
 RECT 1.31 2.05 1.44 2.18 ;
 RECT 21.5 0.505 21.63 0.635 ;
 RECT 7.695 2.015 7.825 2.145 ;
 RECT 23.435 0.12 23.565 0.25 ;
 RECT 23 1.485 23.13 1.615 ;
 RECT 25.395 1.465 25.525 1.595 ;
 RECT 15.94 1.705 16.07 1.835 ;
 RECT 25.395 0.595 25.525 0.725 ;
 RECT 3.77 1.525 3.9 1.655 ;
 RECT 9.32 2.225 9.45 2.355 ;
 RECT 18.3 0.975 18.43 1.105 ;
 RECT 19.29 2.64 19.42 2.77 ;
 RECT 0.84 1.67 0.97 1.8 ;
 RECT 17.785 0.36 17.915 0.49 ;
 RECT 19.875 0.63 20.005 0.76 ;
 RECT 23.94 0.595 24.07 0.725 ;
 RECT 3.375 0.525 3.505 0.655 ;
 RECT 4.42 1.825 4.55 1.955 ;
 RECT 24.45 1.49 24.58 1.62 ;
 RECT 16.415 1.705 16.545 1.835 ;
 RECT 17.7 2.64 17.83 2.77 ;
 RECT 24.08 1.405 24.21 1.535 ;
 RECT 7.7 0.905 7.83 1.035 ;
 RECT 5.84 0.315 5.97 0.445 ;
 RECT 8.175 0.905 8.305 1.035 ;
 RECT 11.45 0.595 11.58 0.725 ;
 RECT 9.51 0.62 9.64 0.75 ;
 RECT 23.605 1.445 23.735 1.575 ;
 RECT 0.34 1.825 0.47 1.955 ;
 RECT 14.475 1.035 14.605 1.165 ;
 RECT 15.06 0.91 15.19 1.04 ;
 LAYER M1 ;
 RECT 21.295 1.225 21.525 1.245 ;
 RECT 21.295 1.195 21.885 1.225 ;
 RECT 21.435 1.015 21.745 1.035 ;
 RECT 21.295 1.035 21.745 1.055 ;
 RECT 21.57 0.64 21.71 1.015 ;
 RECT 21.745 1.225 21.885 1.75 ;
 RECT 21.45 0.5 21.71 0.64 ;
 RECT 22.345 1.035 22.575 1.055 ;
 RECT 22.345 1.195 22.575 1.245 ;
 RECT 21.295 1.055 22.575 1.195 ;
 RECT 23.315 1.145 23.455 1.345 ;
 RECT 22.995 1.485 23.135 1.76 ;
 RECT 23.315 0.73 23.455 0.935 ;
 RECT 22.995 0.355 23.135 0.59 ;
 RECT 22.995 1.345 23.455 1.485 ;
 RECT 23.27 0.935 23.5 1.145 ;
 RECT 22.995 0.59 23.455 0.73 ;
 RECT 20.255 0.36 20.485 0.43 ;
 RECT 21.85 0.36 21.99 0.565 ;
 RECT 20.255 0.22 21.99 0.36 ;
 RECT 22.59 0.705 22.73 0.75 ;
 RECT 22.715 0.995 23.02 1.205 ;
 RECT 22.715 0.89 22.855 0.995 ;
 RECT 22.59 0.75 22.855 0.89 ;
 RECT 21.85 0.565 22.73 0.705 ;
 RECT 15.49 0.775 15.63 1.405 ;
 RECT 16.215 0.56 16.445 0.635 ;
 RECT 14.47 1.405 15.63 1.545 ;
 RECT 14.47 1.545 14.61 1.83 ;
 RECT 13.425 1.83 14.675 1.97 ;
 RECT 14.47 1.17 14.61 1.405 ;
 RECT 14.4 1.03 14.68 1.17 ;
 RECT 18.41 0.36 18.55 0.635 ;
 RECT 15.49 0.635 18.55 0.775 ;
 RECT 19.09 0.36 19.23 1.25 ;
 RECT 19.09 1.25 19.32 1.46 ;
 RECT 18.41 0.22 19.23 0.36 ;
 RECT 14.595 0.28 16.99 0.42 ;
 RECT 14.595 0.42 14.825 0.6 ;
 RECT 16.76 0.22 16.99 0.28 ;
 RECT 16.76 0.42 16.99 0.43 ;
 RECT 11.445 0.525 11.585 0.885 ;
 RECT 11.445 1.095 11.585 2.065 ;
 RECT 11.445 0.885 11.72 1.095 ;
 RECT 8.17 1.04 8.31 2.34 ;
 RECT 8.17 0.895 8.31 0.9 ;
 RECT 8.965 2.055 9.105 2.34 ;
 RECT 8.1 0.9 8.375 1.04 ;
 RECT 8.17 2.34 9.105 2.48 ;
 RECT 9.49 1.66 9.63 1.915 ;
 RECT 8.965 1.915 9.63 2.055 ;
 RECT 9.49 1.52 11.08 1.66 ;
 RECT 10.94 0.525 11.08 1.52 ;
 RECT 10.94 1.66 11.08 2.11 ;
 RECT 10.415 0.765 10.555 1.52 ;
 RECT 10.415 1.66 10.555 2.145 ;
 RECT 13.75 0.57 13.98 0.95 ;
 RECT 12.17 0.585 13.125 0.63 ;
 RECT 12.895 0.63 13.125 0.665 ;
 RECT 12.895 0.455 13.125 0.49 ;
 RECT 12.195 0.49 13.125 0.585 ;
 RECT 12.17 0.63 12.4 0.795 ;
 RECT 3.765 0.895 7.45 1.035 ;
 RECT 7.22 1.035 7.45 1.105 ;
 RECT 3.765 0.66 3.905 0.895 ;
 RECT 3.305 0.52 3.905 0.66 ;
 RECT 1.865 0.88 2.005 1.475 ;
 RECT 1.825 1.63 1.965 1.99 ;
 RECT 1.825 1.475 2.17 1.63 ;
 RECT 1.715 1.99 1.965 2.13 ;
 RECT 1.865 0.74 2.185 0.88 ;
 RECT 3.31 1.82 4.89 1.96 ;
 RECT 4.75 1.79 4.89 1.82 ;
 RECT 3.395 1.96 3.675 2.215 ;
 RECT 3.485 0.805 3.625 1.22 ;
 RECT 3.31 1.22 3.625 1.36 ;
 RECT 3.31 1.36 3.45 1.82 ;
 RECT 5.95 1.615 6.18 1.65 ;
 RECT 5.95 1.79 6.18 1.825 ;
 RECT 4.75 1.65 6.185 1.79 ;
 RECT 13.74 1.23 13.88 1.42 ;
 RECT 11.89 1.09 13.88 1.23 ;
 RECT 11.89 0.385 12.03 1.09 ;
 RECT 9.88 0.385 10.02 0.9 ;
 RECT 9.88 0.255 12.03 0.385 ;
 RECT 9.88 0.245 12.025 0.255 ;
 RECT 8.965 0.9 10.02 1.04 ;
 RECT 8.965 0.745 9.105 0.9 ;
 RECT 4.045 0.605 9.105 0.745 ;
 RECT 5.39 0.5 5.62 0.605 ;
 RECT 4.045 0.485 4.36 0.605 ;
 RECT 14.085 1.39 14.315 1.42 ;
 RECT 13.74 1.42 14.315 1.56 ;
 RECT 14.085 1.56 14.315 1.6 ;
 RECT 0.615 0.875 0.755 1.195 ;
 RECT 0.615 1.335 0.755 1.665 ;
 RECT 0.615 1.665 1.02 1.805 ;
 RECT 0.615 0.735 1.04 0.875 ;
 RECT 1.585 0.6 1.725 1.195 ;
 RECT 0.615 1.195 1.725 1.335 ;
 RECT 3.015 0.36 3.155 2.035 ;
 RECT 2.33 0.22 3.155 0.36 ;
 RECT 2.33 0.36 2.47 0.46 ;
 RECT 2.97 2.17 3.11 2.305 ;
 RECT 2.97 2.035 3.155 2.17 ;
 RECT 1.585 0.46 2.47 0.6 ;
 RECT 2.62 1.67 2.76 1.82 ;
 RECT 2.62 1.96 2.76 2.445 ;
 RECT 4.98 2.585 5.21 2.655 ;
 RECT 2.62 2.585 2.76 2.65 ;
 RECT 2.62 0.5 2.76 1.44 ;
 RECT 2.62 1.44 2.875 1.67 ;
 RECT 2.49 1.82 2.76 1.96 ;
 RECT 2.62 2.445 5.21 2.585 ;
 RECT 12.86 1.895 13 2.39 ;
 RECT 17.005 2.205 17.145 2.39 ;
 RECT 12.86 2.39 17.145 2.53 ;
 RECT 11.735 1.755 13 1.895 ;
 RECT 11.735 1.895 11.875 2.34 ;
 RECT 10.465 2.3 10.695 2.34 ;
 RECT 10.465 2.48 10.695 2.51 ;
 RECT 10.465 2.34 11.875 2.48 ;
 RECT 20.89 2.205 21.03 2.52 ;
 RECT 17.005 2.065 21.03 2.205 ;
 RECT 25.23 2.48 25.37 2.52 ;
 RECT 20.89 2.52 25.37 2.66 ;
 RECT 25.23 2.27 25.46 2.48 ;
 RECT 16.3 1.7 16.595 1.84 ;
 RECT 16.3 1.84 16.44 2.075 ;
 RECT 15.605 1.84 15.745 2.075 ;
 RECT 15.41 1.7 15.745 1.84 ;
 RECT 15.605 2.075 16.44 2.215 ;
 RECT 16.495 1.055 16.635 1.245 ;
 RECT 15.935 1.385 16.075 1.625 ;
 RECT 16.775 1.385 17.005 1.455 ;
 RECT 15.935 1.245 17.005 1.385 ;
 RECT 16.465 0.915 16.765 1.055 ;
 RECT 15.905 1.625 16.16 1.92 ;
 RECT 13.14 1.56 13.28 2.11 ;
 RECT 13.14 2.11 15.465 2.245 ;
 RECT 13.14 2.245 15.46 2.25 ;
 RECT 15.235 2.035 15.465 2.11 ;
 RECT 12.09 1.405 12.32 1.42 ;
 RECT 12.09 1.56 12.32 1.615 ;
 RECT 12.09 1.42 13.28 1.56 ;
 RECT 9.205 1.21 9.345 1.635 ;
 RECT 8.615 1.04 8.755 1.475 ;
 RECT 8.455 1.475 8.755 1.635 ;
 RECT 8.615 1.685 9.345 1.775 ;
 RECT 8.615 1.775 8.755 2.18 ;
 RECT 8.455 1.635 9.345 1.685 ;
 RECT 8.545 0.9 8.82 1.04 ;
 RECT 3.87 2.105 5.09 2.245 ;
 RECT 4.43 1.225 7.08 1.25 ;
 RECT 6.375 1.365 6.515 2.25 ;
 RECT 4.43 1.365 4.57 1.5 ;
 RECT 3.6 1.64 4.105 1.675 ;
 RECT 3.6 1.5 4.57 1.64 ;
 RECT 7.69 1.04 7.83 1.25 ;
 RECT 7.69 1.39 7.83 2.215 ;
 RECT 7.69 0.885 7.83 0.9 ;
 RECT 4.43 1.25 7.83 1.365 ;
 RECT 6.94 1.365 7.83 1.39 ;
 RECT 7.625 0.9 7.9 1.04 ;
 RECT 23.935 0.73 24.075 1.04 ;
 RECT 24.075 1.18 24.215 1.605 ;
 RECT 23.87 0.59 24.145 0.73 ;
 RECT 25.195 0.99 25.425 1.04 ;
 RECT 23.935 1.04 25.425 1.18 ;
 RECT 25.195 1.18 25.425 1.2 ;
 RECT 24.055 0.29 24.425 0.43 ;
 RECT 24.285 0.43 24.425 0.71 ;
 RECT 24.055 0.22 24.285 0.29 ;
 RECT 25.705 0.85 25.845 1.385 ;
 RECT 25.39 1.525 25.53 1.73 ;
 RECT 24.285 0.71 25.845 0.85 ;
 RECT 25.39 0.51 25.53 0.71 ;
 RECT 25.39 1.385 25.845 1.525 ;
 END
END RDFFNSRASX1

MACRO ISOLANDX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.395 1.445 0.79 1.725 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END ISO

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.335 1.185 1.755 1.565 ;
 RECT 1.335 1.125 1.555 1.185 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.01 1.28 2.4 1.6 ;
 RECT 2.01 1.6 2.15 2.505 ;
 RECT 2.2 0.365 2.34 1.28 ;
 END
 ANTENNADIFFAREA 0.503 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 RECT 0.51 2.14 0.725 2.28 ;
 RECT 0.79 2.48 1.275 2.8 ;
 RECT 0.51 2.28 0.65 2.8 ;
 RECT 1.525 1.825 1.665 2.8 ;
 RECT 0.585 1.87 0.725 2.14 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 RECT 0.52 0.75 0.785 0.89 ;
 RECT 0.905 0.08 1.395 0.42 ;
 RECT 1.73 0.08 1.87 0.57 ;
 RECT 0.585 0.08 0.725 0.75 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.84 0.52 0.94 1.06 ;
 RECT 0.84 1.29 0.94 2.38 ;
 RECT 0.71 1.06 0.94 1.29 ;
 RECT 0.37 0.515 0.47 1.47 ;
 RECT 0.37 1.7 0.47 2.41 ;
 RECT 0.365 1.47 0.595 1.7 ;
 RECT 1.14 1.125 1.555 1.265 ;
 RECT 1.14 0.52 1.24 1.125 ;
 RECT 1.31 1.265 1.555 1.355 ;
 RECT 1.31 1.355 1.41 2.405 ;
 RECT 1.78 0.985 2.085 1.09 ;
 RECT 1.78 1.09 1.88 2.775 ;
 RECT 1.83 0.86 2.085 0.985 ;
 RECT 1.985 0.1 2.085 0.86 ;
 LAYER CO ;
 RECT 1.215 0.255 1.345 0.385 ;
 RECT 0.955 0.255 1.085 0.385 ;
 RECT 1.1 2.53 1.23 2.66 ;
 RECT 0.84 2.53 0.97 2.66 ;
 RECT 1.88 0.91 2.01 1.04 ;
 RECT 1.375 1.175 1.505 1.305 ;
 RECT 0.76 1.11 0.89 1.24 ;
 RECT 2.205 0.42 2.335 0.55 ;
 RECT 2.015 1.6 2.145 1.73 ;
 RECT 2.015 1.93 2.145 2.06 ;
 RECT 2.015 2.305 2.145 2.435 ;
 RECT 1.735 0.39 1.865 0.52 ;
 RECT 1.53 2.305 1.66 2.435 ;
 RECT 0.415 1.52 0.545 1.65 ;
 RECT 1.36 0.755 1.49 0.885 ;
 RECT 1.53 1.965 1.66 2.095 ;
 RECT 1.06 1.93 1.19 2.06 ;
 RECT 0.59 0.755 0.72 0.885 ;
 RECT 0.59 1.93 0.72 2.06 ;
 RECT 0.12 0.755 0.25 0.885 ;
 RECT 0.12 1.93 0.25 2.06 ;
 LAYER M1 ;
 RECT 0.115 0.645 0.255 1.105 ;
 RECT 0.115 1.245 0.255 2.11 ;
 RECT 0.755 1.04 0.895 1.105 ;
 RECT 0.755 1.245 0.895 1.3 ;
 RECT 0.115 1.105 0.895 1.245 ;
 RECT 1.055 0.89 1.195 2.11 ;
 RECT 1.81 0.89 2.06 1.045 ;
 RECT 1.055 0.75 2.06 0.89 ;
 END
END ISOLANDX1

MACRO BSLEX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 RECT 2.11 1.925 2.25 2.8 ;
 RECT 0.285 1.54 0.425 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 RECT 2.095 0.08 2.235 0.825 ;
 RECT 0.285 0.08 0.425 0.66 ;
 END
 END VSS

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 0.835 0.615 1.11 ;
 END
 ANTENNAGATEAREA 0.073 ;
 END ENB

 PIN INOUT2
 DIRECTION INOUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.13 1.085 1.43 1.455 ;
 RECT 1.13 1.455 1.27 2.61 ;
 RECT 1.13 0.44 1.27 1.085 ;
 END
 ANTENNADIFFAREA 0.429 ;
 END INOUT2

 PIN INOUT1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.6 1.72 1.74 2.61 ;
 RECT 1.6 1.48 2.04 1.72 ;
 RECT 1.6 0.415 1.74 1.48 ;
 END
 ANTENNADIFFAREA 0.429 ;
 END INOUT1

 OBS
 LAYER PO ;
 RECT 0.385 0.85 0.64 0.895 ;
 RECT 0.385 0.995 0.64 1.08 ;
 RECT 0.385 0.895 1.485 0.995 ;
 RECT 1.385 0.175 1.485 0.895 ;
 RECT 0.54 0.34 0.64 0.85 ;
 RECT 0.54 1.08 0.64 1.965 ;
 RECT 0.665 2.68 1.485 2.78 ;
 RECT 1.385 1.3 1.485 2.68 ;
 RECT 0.665 2.455 0.895 2.68 ;
 LAYER CO ;
 RECT 0.435 0.9 0.565 1.03 ;
 RECT 0.715 2.505 0.845 2.635 ;
 RECT 1.605 0.49 1.735 0.62 ;
 RECT 2.115 1.975 2.245 2.105 ;
 RECT 2.1 0.38 2.23 0.51 ;
 RECT 1.605 2.43 1.735 2.56 ;
 RECT 0.76 1.575 0.89 1.705 ;
 RECT 0.76 0.525 0.89 0.655 ;
 RECT 0.29 0.48 0.42 0.61 ;
 RECT 0.29 1.59 0.42 1.72 ;
 RECT 2.1 0.645 2.23 0.775 ;
 RECT 2.115 2.245 2.245 2.375 ;
 RECT 1.135 0.49 1.265 0.62 ;
 RECT 1.135 1.885 1.265 2.015 ;
 RECT 1.135 1.615 1.265 1.745 ;
 RECT 1.605 1.635 1.735 1.765 ;
 RECT 1.605 1.895 1.735 2.025 ;
 RECT 1.605 2.165 1.735 2.295 ;
 RECT 1.135 2.155 1.265 2.285 ;
 RECT 1.135 2.43 1.265 2.56 ;
 LAYER M1 ;
 RECT 0.76 1.575 0.89 1.705 ;
 RECT 0.76 0.525 0.89 0.655 ;
 RECT 0.755 0.475 0.895 2.585 ;
 RECT 0.715 2.505 0.845 2.635 ;
 RECT 0.665 2.455 0.895 2.655 ;
 END
END BSLEX1

MACRO BSLEX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 2.755 1.98 2.895 2.8 ;
 RECT 0.225 1.555 0.365 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 0.225 0.08 0.365 0.85 ;
 RECT 2.755 0.08 2.895 0.83 ;
 END
 END VSS

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 1.12 0.555 1.4 ;
 END
 ANTENNAGATEAREA 0.146 ;
 END ENB

 PIN INOUT1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.24 1.48 2.68 1.72 ;
 RECT 1.25 0.22 2.38 0.36 ;
 RECT 1.08 0.54 1.46 0.68 ;
 RECT 1.08 1.24 1.39 1.38 ;
 RECT 2.24 1.72 2.38 2.615 ;
 RECT 2.24 0.36 2.38 1.48 ;
 RECT 1.25 0.36 1.39 0.54 ;
 RECT 1.25 1.38 1.39 2.615 ;
 RECT 1.08 0.68 1.22 1.24 ;
 END
 ANTENNADIFFAREA 1.029 ;
 END INOUT1

 PIN INOUT2
 DIRECTION INOUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.76 1.08 1.9 2.615 ;
 RECT 1.48 0.84 1.9 1.08 ;
 RECT 1.76 0.51 1.9 0.84 ;
 END
 ANTENNADIFFAREA 0.556 ;
 END INOUT2

 OBS
 LAYER PO ;
 RECT 0.48 0.425 0.58 0.94 ;
 RECT 0.48 0.94 2.115 1.04 ;
 RECT 0.48 1.04 0.58 1.12 ;
 RECT 1.525 0.27 1.625 0.94 ;
 RECT 2.015 0.27 2.115 0.94 ;
 RECT 0.48 1.35 0.58 2.265 ;
 RECT 0.35 1.12 0.58 1.35 ;
 RECT 1.525 1.305 1.625 2.685 ;
 RECT 2.015 1.305 2.115 2.685 ;
 RECT 0.76 2.685 2.115 2.785 ;
 RECT 0.76 2.455 0.99 2.685 ;
 LAYER CO ;
 RECT 0.7 0.67 0.83 0.8 ;
 RECT 0.23 1.605 0.36 1.735 ;
 RECT 0.23 1.875 0.36 2.005 ;
 RECT 0.7 1.605 0.83 1.735 ;
 RECT 0.7 1.875 0.83 2.005 ;
 RECT 1.255 0.545 1.385 0.675 ;
 RECT 1.255 2.435 1.385 2.565 ;
 RECT 1.255 1.89 1.385 2.02 ;
 RECT 1.255 1.62 1.385 1.75 ;
 RECT 1.255 2.16 1.385 2.29 ;
 RECT 2.76 0.65 2.89 0.78 ;
 RECT 2.76 2.3 2.89 2.43 ;
 RECT 1.765 1.89 1.895 2.02 ;
 RECT 1.765 1.62 1.895 1.75 ;
 RECT 2.245 1.635 2.375 1.765 ;
 RECT 2.245 1.895 2.375 2.025 ;
 RECT 2.245 2.165 2.375 2.295 ;
 RECT 2.245 2.435 2.375 2.565 ;
 RECT 1.765 2.16 1.895 2.29 ;
 RECT 1.765 2.435 1.895 2.565 ;
 RECT 0.4 1.17 0.53 1.3 ;
 RECT 0.81 2.505 0.94 2.635 ;
 RECT 0.4 1.17 0.53 1.3 ;
 RECT 0.81 2.505 0.94 2.635 ;
 RECT 2.76 0.38 2.89 0.51 ;
 RECT 2.76 2.03 2.89 2.16 ;
 RECT 2.245 0.545 2.375 0.675 ;
 RECT 1.765 0.585 1.895 0.715 ;
 RECT 0.23 0.67 0.36 0.8 ;
 LAYER M1 ;
 RECT 0.7 0.67 0.83 0.8 ;
 RECT 0.7 1.605 0.83 1.735 ;
 RECT 0.7 1.875 0.83 2.005 ;
 RECT 0.695 0.62 0.835 2.66 ;
 RECT 0.695 2.455 0.99 2.66 ;
 RECT 0.81 2.505 0.94 2.635 ;
 END
END BSLEX2

MACRO BSLEX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 3.93 2.01 4.07 2.8 ;
 RECT 0.36 1.765 0.5 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 3.93 0.08 4.07 0.835 ;
 RECT 0.36 0.08 0.5 0.595 ;
 END
 END VSS

 PIN INOUT2
 DIRECTION INOUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.415 1.48 3.96 1.72 ;
 RECT 1.485 0.245 3.555 0.385 ;
 RECT 3.415 1.72 3.555 2.58 ;
 RECT 2.425 0.385 2.565 2.305 ;
 RECT 1.485 0.385 1.625 2.58 ;
 RECT 3.415 0.385 3.555 1.48 ;
 END
 ANTENNADIFFAREA 1.428 ;
 END INOUT2

 PIN INOUT1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.8 1.16 2.095 1.4 ;
 RECT 1.955 0.525 2.095 1.16 ;
 RECT 1.955 1.4 2.095 2.52 ;
 RECT 2.935 0.525 3.075 2.52 ;
 RECT 1.95 2.52 3.075 2.66 ;
 END
 ANTENNADIFFAREA 1.084 ;
 END INOUT1

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 0.84 0.69 1.175 ;
 END
 ANTENNAGATEAREA 0.292 ;
 END ENB

 OBS
 LAYER PO ;
 RECT 1.74 1.37 1.84 2.65 ;
 RECT 2.21 1.27 2.31 2.65 ;
 RECT 2.7 1.27 2.8 2.65 ;
 RECT 3.19 1.27 3.29 2.65 ;
 RECT 1.74 2.65 3.29 2.75 ;
 RECT 1.11 1.37 1.34 1.48 ;
 RECT 1.11 1.27 1.84 1.37 ;
 RECT 0.46 0.965 0.715 0.985 ;
 RECT 0.46 0.985 3.29 1.085 ;
 RECT 0.46 1.085 0.715 1.175 ;
 RECT 1.74 0.285 1.84 0.985 ;
 RECT 2.21 0.285 2.31 0.985 ;
 RECT 2.7 0.285 2.8 0.985 ;
 RECT 3.19 0.285 3.29 0.985 ;
 RECT 0.615 0.14 0.715 0.965 ;
 RECT 0.615 1.175 0.715 2.75 ;
 LAYER CO ;
 RECT 3.42 2.4 3.55 2.53 ;
 RECT 2.94 2.125 3.07 2.255 ;
 RECT 2.94 2.4 3.07 2.53 ;
 RECT 3.935 2.06 4.065 2.19 ;
 RECT 3.935 0.375 4.065 0.505 ;
 RECT 0.365 2.4 0.495 2.53 ;
 RECT 0.835 2.4 0.965 2.53 ;
 RECT 0.365 2.125 0.495 2.255 ;
 RECT 0.835 2.125 0.965 2.255 ;
 RECT 0.365 1.855 0.495 1.985 ;
 RECT 0.835 1.855 0.965 1.985 ;
 RECT 0.835 1.585 0.965 1.715 ;
 RECT 0.835 0.39 0.965 0.52 ;
 RECT 0.835 0.68 0.965 0.81 ;
 RECT 0.365 0.39 0.495 0.52 ;
 RECT 3.42 0.585 3.55 0.715 ;
 RECT 2.94 0.585 3.07 0.715 ;
 RECT 1.16 1.31 1.29 1.44 ;
 RECT 0.51 1.005 0.64 1.135 ;
 RECT 2.43 0.585 2.56 0.715 ;
 RECT 1.96 0.585 2.09 0.715 ;
 RECT 1.49 0.585 1.62 0.715 ;
 RECT 1.49 2.125 1.62 2.255 ;
 RECT 1.49 2.4 1.62 2.53 ;
 RECT 1.49 1.855 1.62 1.985 ;
 RECT 1.49 1.585 1.62 1.715 ;
 RECT 1.96 2.125 2.09 2.255 ;
 RECT 1.96 2.4 2.09 2.53 ;
 RECT 1.96 1.855 2.09 1.985 ;
 RECT 1.96 1.585 2.09 1.715 ;
 RECT 2.43 1.855 2.56 1.985 ;
 RECT 2.43 1.585 2.56 1.715 ;
 RECT 2.43 2.125 2.56 2.255 ;
 RECT 3.935 0.645 4.065 0.775 ;
 RECT 3.935 2.33 4.065 2.46 ;
 RECT 2.94 1.855 3.07 1.985 ;
 RECT 2.94 1.585 3.07 1.715 ;
 RECT 3.42 1.6 3.55 1.73 ;
 RECT 3.42 1.86 3.55 1.99 ;
 RECT 3.42 2.13 3.55 2.26 ;
 LAYER M1 ;
 RECT 0.835 2.4 0.965 2.53 ;
 RECT 0.835 2.125 0.965 2.255 ;
 RECT 0.835 1.855 0.965 1.985 ;
 RECT 0.835 1.585 0.965 1.715 ;
 RECT 0.835 0.39 0.965 0.52 ;
 RECT 0.835 0.68 0.965 0.81 ;
 RECT 0.83 0.34 0.97 2.58 ;
 RECT 0.845 1.27 1.315 1.41 ;
 RECT 1.11 1.27 1.34 1.48 ;
 END
END BSLEX4

MACRO RSDFFNX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 23.04 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 1.295 1.39 1.635 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.65 1.64 2.095 1.97 ;
 RECT 1.63 1.085 1.93 1.225 ;
 RECT 1.79 1.225 1.93 1.64 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.925 0.32 2.295 0.615 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.27 1.125 9.6 1.415 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.525 1.5 11.665 2.295 ;
 RECT 11.525 1.09 11.945 1.5 ;
 RECT 11.525 0.525 11.665 1.09 ;
 END
 ANTENNADIFFAREA 0.504 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.575 1.43 12.715 1.79 ;
 RECT 12.575 1.135 12.945 1.43 ;
 RECT 12.575 0.48 12.715 1.135 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 23.04 2.96 ;
 RECT 7.875 2.615 8.11 2.8 ;
 RECT 9.34 2.37 9.61 2.51 ;
 RECT 4.225 2.51 4.495 2.65 ;
 RECT 5.92 2.51 6.15 2.65 ;
 RECT 2.565 2.135 2.965 2.275 ;
 RECT 1.07 2.115 1.21 2.8 ;
 RECT 12.095 2.275 12.235 2.8 ;
 RECT 0.185 1.64 0.345 2.8 ;
 RECT 10.58 1.94 10.72 2.8 ;
 RECT 14.825 2.025 14.965 2.8 ;
 RECT 13.135 2 13.275 2.8 ;
 RECT 9.405 2.51 9.545 2.8 ;
 RECT 4.29 2.65 4.43 2.8 ;
 RECT 5.965 2.65 6.105 2.8 ;
 RECT 2.825 2.275 2.965 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 23.04 0.08 ;
 RECT 9.33 0.555 9.6 0.695 ;
 RECT 5.93 0.555 6.18 0.695 ;
 RECT 17.785 0.22 18.035 0.36 ;
 RECT 20.55 0.08 20.69 0.65 ;
 RECT 0.185 0.08 0.345 0.84 ;
 RECT 1.07 0.08 1.21 0.96 ;
 RECT 10.58 0.08 10.72 0.785 ;
 RECT 4.29 0.08 4.43 0.32 ;
 RECT 14.825 0.08 14.965 0.815 ;
 RECT 7.94 0.08 8.08 0.78 ;
 RECT 2.63 0.08 2.77 0.96 ;
 RECT 12.095 0.08 12.235 0.575 ;
 RECT 13.185 0.08 13.325 0.865 ;
 RECT 9.395 0.08 9.535 0.555 ;
 RECT 5.995 0.08 6.135 0.555 ;
 RECT 17.83 0.08 17.97 0.22 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 21.405 1.4 21.745 1.765 ;
 RECT 17.83 2.235 21.56 2.375 ;
 RECT 17.785 1.47 18.015 1.61 ;
 RECT 20.505 1.395 20.645 2.235 ;
 RECT 21.42 1.765 21.56 2.235 ;
 RECT 17.83 1.61 17.97 2.235 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 15.955 0.81 16.335 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 19.445 0.865 19.825 0.965 ;
 RECT 2.405 0.51 2.505 2.45 ;
 RECT 2.38 2.45 2.61 2.66 ;
 RECT 13.47 0.385 13.57 2.405 ;
 RECT 13.37 2.405 13.6 2.635 ;
 RECT 9.675 0.33 9.775 1.175 ;
 RECT 9.675 1.395 9.775 2.235 ;
 RECT 9.415 1.175 9.775 1.395 ;
 RECT 18.54 0.865 19.265 0.965 ;
 RECT 18.54 0.735 18.77 0.865 ;
 RECT 19.165 0.275 19.265 0.865 ;
 RECT 9.135 0.33 9.235 2.135 ;
 RECT 9.015 2.135 9.245 2.365 ;
 RECT 4.05 0.38 4.15 1.23 ;
 RECT 4.05 1.46 4.15 2.34 ;
 RECT 4.05 1.23 4.28 1.46 ;
 RECT 2.885 1.58 2.985 2.56 ;
 RECT 2.885 0.515 2.985 1.37 ;
 RECT 2.735 1.37 2.985 1.58 ;
 RECT 13.78 1.835 13.88 2.425 ;
 RECT 13.77 1.605 14 1.835 ;
 RECT 10.87 0.365 10.97 1.16 ;
 RECT 10.675 1.16 10.97 1.22 ;
 RECT 10.87 1.39 10.97 2.47 ;
 RECT 10.675 1.32 10.97 1.39 ;
 RECT 10.675 1.22 11.88 1.32 ;
 RECT 11.78 0.105 11.88 1.22 ;
 RECT 11.78 1.32 11.88 2.75 ;
 RECT 7.065 1.445 7.165 2.285 ;
 RECT 6.98 2.285 7.21 2.515 ;
 RECT 12.36 0.105 15.735 0.205 ;
 RECT 12.36 0.205 12.46 0.87 ;
 RECT 14.265 0.205 14.365 0.925 ;
 RECT 15.505 0.205 15.735 0.4 ;
 RECT 12.36 1.085 12.46 2.755 ;
 RECT 12.215 0.87 12.46 1.085 ;
 RECT 14.14 0.925 14.37 1.135 ;
 RECT 5.775 0.84 6.02 0.87 ;
 RECT 5.775 0.97 6.02 1.06 ;
 RECT 5.775 0.38 5.875 0.84 ;
 RECT 6.25 0.38 6.35 0.87 ;
 RECT 5.775 0.87 6.35 0.97 ;
 RECT 4.545 0.1 7.24 0.2 ;
 RECT 7.14 0.42 7.24 0.95 ;
 RECT 6.94 0.2 7.24 0.42 ;
 RECT 4.545 0.2 4.645 0.97 ;
 RECT 7.67 0.37 7.77 1.21 ;
 RECT 7.67 1.42 7.77 2.16 ;
 RECT 7.67 1.21 7.955 1.42 ;
 RECT 2.1 0.635 2.2 1.45 ;
 RECT 1.63 1.55 1.73 2.55 ;
 RECT 1.97 0.405 2.2 0.635 ;
 RECT 1.63 1.45 2.2 1.55 ;
 RECT 1.195 1.33 1.425 1.395 ;
 RECT 1.195 1.495 1.425 1.56 ;
 RECT 0.855 1.395 1.425 1.495 ;
 RECT 1.325 0.51 1.425 1.33 ;
 RECT 1.325 1.56 1.425 2.55 ;
 RECT 0.855 0.51 0.955 1.395 ;
 RECT 0.855 1.495 0.955 2.55 ;
 RECT 20.2 0.275 20.3 1.025 ;
 RECT 20.2 1.255 20.3 1.86 ;
 RECT 20.2 1.025 20.48 1.255 ;
 RECT 8.22 0.37 8.32 2.68 ;
 RECT 10.09 2.475 10.32 2.68 ;
 RECT 8.22 2.68 10.32 2.78 ;
 RECT 4.945 0.38 5.045 0.945 ;
 RECT 4.945 1.175 5.045 2.36 ;
 RECT 4.825 0.945 5.055 1.175 ;
 RECT 6.24 1.75 6.34 2.585 ;
 RECT 6.11 1.53 6.34 1.63 ;
 RECT 6.11 1.73 6.34 1.75 ;
 RECT 5.77 1.73 5.87 2.34 ;
 RECT 5.77 1.63 6.34 1.73 ;
 RECT 14.31 2.605 15.66 2.695 ;
 RECT 14.315 2.695 15.66 2.705 ;
 RECT 14.31 1.425 14.41 2.605 ;
 RECT 13.775 0.385 13.875 1.325 ;
 RECT 13.775 1.325 14.41 1.425 ;
 RECT 15.43 2.475 15.66 2.605 ;
 RECT 4.635 1.76 4.735 2.34 ;
 RECT 4.515 1.53 4.745 1.76 ;
 RECT 1.63 0.5 1.73 1.04 ;
 RECT 1.63 1.04 1.86 1.27 ;
 RECT 20.805 0.27 20.905 0.745 ;
 RECT 20.805 0.975 20.905 1.855 ;
 RECT 20.66 0.745 20.905 0.975 ;
 RECT 5.47 1.34 5.7 1.45 ;
 RECT 5.47 0.38 5.57 1.24 ;
 RECT 5.47 1.45 5.57 2.345 ;
 RECT 6.565 0.38 6.665 1.24 ;
 RECT 6.565 1.34 6.665 2.585 ;
 RECT 5.47 1.24 6.665 1.34 ;
 RECT 1.91 1.73 2.2 1.96 ;
 RECT 2.1 1.96 2.2 2.55 ;
 RECT 14.61 0.385 14.71 1.215 ;
 RECT 14.61 1.215 14.885 1.27 ;
 RECT 14.61 1.425 14.71 2.425 ;
 RECT 14.61 1.37 14.885 1.425 ;
 RECT 15.085 1.045 15.185 1.27 ;
 RECT 15.085 1.37 15.185 2.425 ;
 RECT 14.61 1.27 15.185 1.37 ;
 RECT 17.535 1.045 17.635 1.76 ;
 RECT 15.085 0.385 15.185 0.945 ;
 RECT 15.085 0.945 17.635 1.045 ;
 RECT 16.045 0.84 16.275 0.945 ;
 RECT 16.045 1.045 16.275 1.07 ;
 RECT 19.725 1.145 19.825 2.09 ;
 RECT 17.535 0.145 17.635 0.945 ;
 RECT 18.69 1.86 18.79 2.09 ;
 RECT 18.56 1.545 18.79 1.76 ;
 RECT 18.69 2.09 19.825 2.19 ;
 RECT 17.535 1.76 18.79 1.86 ;
 RECT 18.115 0.965 18.215 1.145 ;
 RECT 18.115 1.145 19.545 1.245 ;
 RECT 19.445 0.965 19.545 1.145 ;
 RECT 19.255 1.245 19.355 1.86 ;
 RECT 19.725 0.275 19.825 0.865 ;
 RECT 18.115 0.735 18.345 0.965 ;
 LAYER CO ;
 RECT 0.2 1.97 0.33 2.1 ;
 RECT 0.2 2.23 0.33 2.36 ;
 RECT 17.835 0.225 17.965 0.355 ;
 RECT 7.37 0.6 7.5 0.73 ;
 RECT 7.775 1.25 7.905 1.38 ;
 RECT 2.785 1.41 2.915 1.54 ;
 RECT 11.53 2.105 11.66 2.235 ;
 RECT 12.1 2.34 12.23 2.47 ;
 RECT 14.19 0.965 14.32 1.095 ;
 RECT 0.2 1.71 0.33 1.84 ;
 RECT 2.43 2.49 2.56 2.62 ;
 RECT 20.555 0.47 20.685 0.6 ;
 RECT 20.51 1.455 20.64 1.585 ;
 RECT 19.95 1.435 20.08 1.565 ;
 RECT 19.95 0.505 20.08 0.635 ;
 RECT 19.475 1.415 19.605 1.545 ;
 RECT 19.475 0.505 19.605 0.635 ;
 RECT 18.915 1.415 19.045 1.545 ;
 RECT 18.915 0.505 19.045 0.635 ;
 RECT 12.58 0.555 12.71 0.685 ;
 RECT 10.585 2.01 10.715 2.14 ;
 RECT 10.725 1.21 10.855 1.34 ;
 RECT 10.585 0.605 10.715 0.735 ;
 RECT 11.145 2.025 11.275 2.155 ;
 RECT 11.145 0.605 11.275 0.735 ;
 RECT 9.465 1.215 9.595 1.345 ;
 RECT 7.03 2.335 7.16 2.465 ;
 RECT 6.99 0.24 7.12 0.37 ;
 RECT 6.16 1.57 6.29 1.7 ;
 RECT 5.83 0.89 5.96 1.02 ;
 RECT 5.52 1.28 5.65 1.41 ;
 RECT 4.565 1.58 4.695 1.71 ;
 RECT 4.875 0.995 5.005 1.125 ;
 RECT 1.96 1.78 2.09 1.91 ;
 RECT 10.025 0.56 10.155 0.69 ;
 RECT 10.025 1.83 10.155 1.96 ;
 RECT 9.4 0.56 9.53 0.69 ;
 RECT 8.885 0.57 9.015 0.7 ;
 RECT 8.885 1.48 9.015 1.61 ;
 RECT 9.41 2.375 9.54 2.505 ;
 RECT 7.93 2.63 8.06 2.76 ;
 RECT 3.48 1.935 3.61 2.065 ;
 RECT 3.68 0.6 3.81 0.73 ;
 RECT 7.37 1.48 7.5 1.61 ;
 RECT 6.81 0.6 6.94 0.73 ;
 RECT 6 0.555 6.13 0.685 ;
 RECT 5.2 0.6 5.33 0.73 ;
 RECT 3.11 2.14 3.24 2.27 ;
 RECT 3.11 0.76 3.24 0.89 ;
 RECT 2.635 0.76 2.765 0.89 ;
 RECT 2.635 2.14 2.765 2.27 ;
 RECT 1.85 2.14 1.98 2.27 ;
 RECT 1.85 0.76 1.98 0.89 ;
 RECT 1.075 0.76 1.205 0.89 ;
 RECT 0.605 0.76 0.735 0.89 ;
 RECT 0.605 2.14 0.735 2.27 ;
 RECT 15.555 0.225 15.685 0.355 ;
 RECT 17.835 1.475 17.965 1.605 ;
 RECT 4.1 1.28 4.23 1.41 ;
 RECT 2.02 0.455 2.15 0.585 ;
 RECT 1.68 1.09 1.81 1.22 ;
 RECT 1.68 1.09 1.81 1.22 ;
 RECT 1.245 1.38 1.375 1.51 ;
 RECT 17.23 1.255 17.36 1.385 ;
 RECT 17.185 0.505 17.315 0.635 ;
 RECT 15.48 2.525 15.61 2.655 ;
 RECT 13.42 2.455 13.55 2.585 ;
 RECT 13.82 1.655 13.95 1.785 ;
 RECT 15.31 0.635 15.44 0.765 ;
 RECT 14.83 0.635 14.96 0.765 ;
 RECT 6.81 1.67 6.94 1.8 ;
 RECT 4.295 2.515 4.425 2.645 ;
 RECT 5.97 2.515 6.1 2.645 ;
 RECT 5.2 1.52 5.33 1.65 ;
 RECT 1.075 2.2 1.205 2.33 ;
 RECT 8.505 1.705 8.635 1.835 ;
 RECT 8.505 0.6 8.635 0.73 ;
 RECT 7.945 0.6 8.075 0.73 ;
 RECT 14.83 2.075 14.96 2.205 ;
 RECT 14.015 2.05 14.145 2.18 ;
 RECT 14.015 0.635 14.145 0.765 ;
 RECT 18.59 0.785 18.72 0.915 ;
 RECT 20.71 0.795 20.84 0.925 ;
 RECT 20.3 1.075 20.43 1.205 ;
 RECT 21.035 0.505 21.165 0.635 ;
 RECT 21.035 1.44 21.165 1.57 ;
 RECT 13.19 0.635 13.32 0.765 ;
 RECT 13.14 2.06 13.27 2.19 ;
 RECT 15.31 2.065 15.44 2.195 ;
 RECT 11.53 1.715 11.66 1.845 ;
 RECT 10.14 2.525 10.27 2.655 ;
 RECT 12.265 0.915 12.395 1.045 ;
 RECT 12.58 1.6 12.71 1.73 ;
 RECT 12.1 0.395 12.23 0.525 ;
 RECT 11.53 0.585 11.66 0.715 ;
 RECT 9.065 2.185 9.195 2.315 ;
 RECT 16.095 0.89 16.225 1.02 ;
 RECT 18.61 1.595 18.74 1.725 ;
 RECT 14.705 1.255 14.835 1.385 ;
 RECT 18.165 0.785 18.295 0.915 ;
 RECT 4.295 0.12 4.425 0.25 ;
 RECT 21.455 1.44 21.585 1.57 ;
 RECT 0.2 0.36 0.33 0.49 ;
 RECT 0.2 0.62 0.33 0.75 ;
 LAYER M1 ;
 RECT 18.605 0.92 18.745 1.785 ;
 RECT 18.52 0.78 18.77 0.92 ;
 RECT 14.45 1.845 14.59 2.45 ;
 RECT 13.415 2.385 13.555 2.45 ;
 RECT 13.415 2.45 14.59 2.59 ;
 RECT 13.415 2.59 13.555 2.65 ;
 RECT 15.305 0.585 15.445 1.705 ;
 RECT 14.45 1.705 15.445 1.845 ;
 RECT 15.305 1.845 15.445 2.265 ;
 RECT 14.61 1.17 14.95 1.51 ;
 RECT 11.14 0.385 11.28 2.21 ;
 RECT 11.14 0.24 11.28 0.245 ;
 RECT 11.805 0.385 11.945 0.75 ;
 RECT 11.14 0.245 11.945 0.385 ;
 RECT 12.26 0.89 12.4 1.095 ;
 RECT 11.805 0.75 12.4 0.89 ;
 RECT 10.86 1.775 11 2.435 ;
 RECT 10.3 1.635 11 1.775 ;
 RECT 10.3 1.775 10.44 2.52 ;
 RECT 10.07 2.52 10.44 2.66 ;
 RECT 11.815 2.135 11.955 2.435 ;
 RECT 10.86 2.435 11.955 2.575 ;
 RECT 12.855 1.86 12.995 1.995 ;
 RECT 11.815 1.995 12.995 2.135 ;
 RECT 13.53 2.045 14.195 2.185 ;
 RECT 13.53 1.86 13.67 2.045 ;
 RECT 13.53 0.63 14.195 0.77 ;
 RECT 13.53 0.77 13.67 1.72 ;
 RECT 12.855 1.72 13.67 1.86 ;
 RECT 13.815 1.095 13.955 1.835 ;
 RECT 14.14 0.925 14.37 0.955 ;
 RECT 13.815 0.955 14.37 1.095 ;
 RECT 14.14 1.095 14.37 1.135 ;
 RECT 7.725 1.21 7.955 1.245 ;
 RECT 7.725 1.385 7.955 1.42 ;
 RECT 7.725 1.245 8.64 1.385 ;
 RECT 8.5 0.55 8.64 1.245 ;
 RECT 8.5 1.385 8.64 1.9 ;
 RECT 7.365 0.55 7.505 1.475 ;
 RECT 7.3 1.475 7.57 1.615 ;
 RECT 6.325 0.375 6.465 1.26 ;
 RECT 7.655 0.375 7.795 0.93 ;
 RECT 6.155 1.26 6.465 1.4 ;
 RECT 6.155 1.4 6.295 1.77 ;
 RECT 6.325 0.235 7.795 0.375 ;
 RECT 8.22 0.24 9.02 0.38 ;
 RECT 8.88 0.38 9.02 1.66 ;
 RECT 8.22 0.38 8.36 0.93 ;
 RECT 7.655 0.93 8.36 1.07 ;
 RECT 3.77 1.13 3.91 2.42 ;
 RECT 3.11 2.32 3.25 2.42 ;
 RECT 3.105 2.14 3.25 2.32 ;
 RECT 3.105 0.67 3.245 2.14 ;
 RECT 3.11 2.42 3.91 2.56 ;
 RECT 3.77 0.99 5.055 1.13 ;
 RECT 17.505 0.36 17.645 0.5 ;
 RECT 15.455 0.22 17.645 0.36 ;
 RECT 17.505 0.5 19.05 0.64 ;
 RECT 18.91 0.435 19.05 0.5 ;
 RECT 18.91 0.64 19.05 1.61 ;
 RECT 17.225 0.64 17.365 0.78 ;
 RECT 17.225 0.92 17.365 1.455 ;
 RECT 17.12 0.5 17.365 0.64 ;
 RECT 17.225 0.78 18.36 0.92 ;
 RECT 8.78 1.94 8.92 2.05 ;
 RECT 7.02 2.05 8.92 2.19 ;
 RECT 7.02 1.805 7.16 2.05 ;
 RECT 6.735 1.665 7.16 1.805 ;
 RECT 6.805 0.545 6.945 1.665 ;
 RECT 10.3 0.365 10.44 1.205 ;
 RECT 9.74 0.365 9.88 1.8 ;
 RECT 9.74 0.225 10.44 0.365 ;
 RECT 8.78 1.8 9.88 1.94 ;
 RECT 10.3 1.205 10.925 1.345 ;
 RECT 21.03 0.435 21.17 1.07 ;
 RECT 21.03 1.21 21.17 1.64 ;
 RECT 20.23 1.07 21.17 1.21 ;
 RECT 9.06 2.23 9.2 2.33 ;
 RECT 6.69 2.33 9.2 2.47 ;
 RECT 6.69 2.085 6.83 2.33 ;
 RECT 4.555 1.945 6.83 2.085 ;
 RECT 5.825 0.835 5.965 1.945 ;
 RECT 4.56 1.715 4.7 1.945 ;
 RECT 4.49 1.575 4.765 1.715 ;
 RECT 9.06 2.09 10.16 2.23 ;
 RECT 10.02 0.505 10.16 2.09 ;
 RECT 15.4 2.52 17.645 2.65 ;
 RECT 15.4 2.65 17.635 2.66 ;
 RECT 17.505 1.33 17.645 2.52 ;
 RECT 19.945 0.64 20.085 1.925 ;
 RECT 18.155 1.33 18.295 1.925 ;
 RECT 19.88 0.5 20.13 0.64 ;
 RECT 18.155 1.925 20.085 2.065 ;
 RECT 17.505 1.19 18.295 1.33 ;
 RECT 2.235 1.545 2.375 2.135 ;
 RECT 2.235 0.895 2.375 1.405 ;
 RECT 1.78 2.135 2.375 2.275 ;
 RECT 1.78 0.755 2.375 0.895 ;
 RECT 2.735 1.37 2.965 1.405 ;
 RECT 2.235 1.405 2.965 1.545 ;
 RECT 2.735 1.545 2.965 1.58 ;
 RECT 5.195 0.55 5.335 1.275 ;
 RECT 4.05 1.275 5.335 1.415 ;
 RECT 5.195 1.415 5.335 1.71 ;
 RECT 19.47 0.36 19.61 1.41 ;
 RECT 20.27 0.36 20.41 0.79 ;
 RECT 19.405 1.41 19.675 1.55 ;
 RECT 19.47 0.22 20.41 0.36 ;
 RECT 20.27 0.79 20.89 0.93 ;
 RECT 3.475 0.6 3.88 0.735 ;
 RECT 3.475 0.735 3.615 2.13 ;
 RECT 4.755 0.6 4.895 0.61 ;
 RECT 4.755 0.41 4.895 0.46 ;
 RECT 3.475 0.595 4.895 0.6 ;
 RECT 3.68 0.46 4.895 0.595 ;
 RECT 4.755 0.275 5.655 0.41 ;
 RECT 5.515 0.41 5.655 1.475 ;
 RECT 4.755 0.27 5.59 0.275 ;
 RECT 0.6 0.71 0.74 1.805 ;
 RECT 0.6 1.945 0.74 2.32 ;
 RECT 1.37 1.945 1.51 2.415 ;
 RECT 0.6 1.805 1.51 1.945 ;
 RECT 1.37 2.415 2.61 2.555 ;
 RECT 2.38 2.555 2.61 2.66 ;
 END
END RSDFFNX1

MACRO RSDFFNX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 23.68 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.88 1.285 1.27 1.625 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.61 1.06 1.84 1.275 ;
 RECT 1.64 1.62 2.095 1.965 ;
 RECT 1.64 1.275 1.78 1.62 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.775 0.63 2.165 0.92 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.2 1.145 9.6 1.415 ;
 END
 ANTENNAGATEAREA 0.05 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.185 1.09 12.605 1.5 ;
 RECT 12.185 1.5 12.325 1.855 ;
 RECT 12.185 0.525 12.325 1.09 ;
 END
 ANTENNADIFFAREA 0.618 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.23 1.005 13.565 1.35 ;
 RECT 13.235 1.35 13.375 1.855 ;
 RECT 13.235 0.48 13.375 1.005 ;
 END
 ANTENNADIFFAREA 0.6 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 23.68 2.96 ;
 RECT 7.875 2.615 8.11 2.8 ;
 RECT 5.92 2.51 6.15 2.65 ;
 RECT 4.225 2.51 4.495 2.65 ;
 RECT 9.34 2.37 9.61 2.51 ;
 RECT 2.585 2.135 2.965 2.275 ;
 RECT 0.185 1.64 0.345 2.8 ;
 RECT 11.705 2.275 11.845 2.8 ;
 RECT 10.58 1.94 10.72 2.8 ;
 RECT 15.47 2.025 15.61 2.8 ;
 RECT 13.715 2.275 13.855 2.8 ;
 RECT 1.07 2.14 1.21 2.8 ;
 RECT 12.71 2.275 12.85 2.8 ;
 RECT 5.965 2.65 6.105 2.8 ;
 RECT 4.29 2.65 4.43 2.8 ;
 RECT 9.405 2.51 9.545 2.8 ;
 RECT 2.825 2.275 2.965 2.8 ;
 RECT 2.825 2.08 2.965 2.135 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 23.68 0.08 ;
 RECT 1.025 0.31 1.255 0.45 ;
 RECT 9.33 0.565 9.6 0.705 ;
 RECT 2.585 0.31 2.815 0.45 ;
 RECT 5.93 0.555 6.18 0.695 ;
 RECT 18.43 0.22 18.68 0.36 ;
 RECT 13.71 0.08 13.85 0.575 ;
 RECT 7.94 0.08 8.08 0.78 ;
 RECT 21.195 0.08 21.335 0.65 ;
 RECT 11.625 0.08 11.765 0.575 ;
 RECT 15.47 0.08 15.61 0.815 ;
 RECT 10.58 0.08 10.72 0.785 ;
 RECT 12.755 0.08 12.895 0.575 ;
 RECT 0.185 0.08 0.345 0.84 ;
 RECT 4.29 0.08 4.43 0.32 ;
 RECT 1.07 0.45 1.21 0.49 ;
 RECT 1.07 0.08 1.21 0.31 ;
 RECT 9.395 0.08 9.535 0.565 ;
 RECT 2.63 0.45 2.77 0.485 ;
 RECT 2.63 0.08 2.77 0.31 ;
 RECT 5.995 0.08 6.135 0.555 ;
 RECT 18.475 0.08 18.615 0.22 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 22.05 1.4 22.39 1.765 ;
 RECT 18.475 2.225 22.215 2.385 ;
 RECT 18.43 1.47 18.66 1.61 ;
 RECT 21.15 1.395 21.29 2.225 ;
 RECT 22.065 1.765 22.205 2.225 ;
 RECT 18.475 1.61 18.615 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 16.6 0.81 16.98 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 9.415 1.16 9.775 1.395 ;
 RECT 14.425 1.835 14.525 2.425 ;
 RECT 14.415 1.605 14.645 1.835 ;
 RECT 7.065 1.445 7.165 2.285 ;
 RECT 6.98 2.285 7.21 2.515 ;
 RECT 2.1 1.965 2.2 2.55 ;
 RECT 1.91 1.735 2.2 1.965 ;
 RECT 4.945 0.38 5.045 0.945 ;
 RECT 4.945 1.175 5.045 2.36 ;
 RECT 4.825 0.945 5.055 1.175 ;
 RECT 21.45 0.27 21.55 0.745 ;
 RECT 21.45 0.975 21.55 1.855 ;
 RECT 21.305 0.745 21.55 0.975 ;
 RECT 14.115 0.385 14.215 2.405 ;
 RECT 14.015 2.405 14.245 2.635 ;
 RECT 2.885 0.095 2.985 1.525 ;
 RECT 2.735 1.525 2.985 1.735 ;
 RECT 2.885 1.735 2.985 2.55 ;
 RECT 2.405 0.095 2.505 2.45 ;
 RECT 2.395 2.45 2.625 2.66 ;
 RECT 8.22 0.37 8.32 2.68 ;
 RECT 10.09 2.475 10.32 2.68 ;
 RECT 8.22 2.68 10.32 2.78 ;
 RECT 5.47 1.34 5.7 1.45 ;
 RECT 5.47 1.45 5.57 2.345 ;
 RECT 6.565 0.38 6.665 1.24 ;
 RECT 5.47 1.24 6.665 1.34 ;
 RECT 6.565 1.34 6.665 2.62 ;
 RECT 5.47 0.38 5.57 1.24 ;
 RECT 7.67 0.37 7.77 1.21 ;
 RECT 7.67 1.42 7.77 2.16 ;
 RECT 7.67 1.21 7.955 1.42 ;
 RECT 1.63 0.095 1.73 1.045 ;
 RECT 1.61 1.045 1.84 1.275 ;
 RECT 9.135 0.33 9.235 2.135 ;
 RECT 9.015 2.135 9.245 2.365 ;
 RECT 5.775 0.38 5.875 0.84 ;
 RECT 5.775 0.87 6.35 0.97 ;
 RECT 6.25 0.38 6.35 0.87 ;
 RECT 5.775 0.84 6.02 0.87 ;
 RECT 5.775 0.97 6.02 1.06 ;
 RECT 6.24 1.75 6.34 2.62 ;
 RECT 6.11 1.53 6.34 1.63 ;
 RECT 6.11 1.73 6.34 1.75 ;
 RECT 5.77 1.73 5.87 2.34 ;
 RECT 5.77 1.63 6.34 1.73 ;
 RECT 4.545 0.1 7.24 0.2 ;
 RECT 7.14 0.42 7.24 0.95 ;
 RECT 6.94 0.2 7.24 0.42 ;
 RECT 4.545 0.2 4.645 0.97 ;
 RECT 4.635 1.76 4.735 2.34 ;
 RECT 4.515 1.53 4.745 1.76 ;
 RECT 0.855 1.32 1.145 1.385 ;
 RECT 0.855 0.095 0.955 1.32 ;
 RECT 0.855 1.485 1.145 1.55 ;
 RECT 0.855 1.55 0.955 2.55 ;
 RECT 1.325 0.095 1.425 1.385 ;
 RECT 1.325 1.485 1.425 2.55 ;
 RECT 0.855 1.385 1.425 1.485 ;
 RECT 2.1 0.845 2.2 1.455 ;
 RECT 2.1 0.095 2.2 0.615 ;
 RECT 1.63 1.555 1.73 2.55 ;
 RECT 1.63 1.455 2.2 1.555 ;
 RECT 1.92 0.615 2.2 0.845 ;
 RECT 4.05 0.38 4.15 1.23 ;
 RECT 4.05 1.46 4.15 2.34 ;
 RECT 4.05 1.23 4.28 1.46 ;
 RECT 20.845 0.275 20.945 1.025 ;
 RECT 20.845 1.255 20.945 1.86 ;
 RECT 20.845 1.025 21.125 1.255 ;
 RECT 10.675 1.22 12.54 1.32 ;
 RECT 10.675 1.16 10.97 1.22 ;
 RECT 10.87 0.365 10.97 1.16 ;
 RECT 12.44 0.105 12.54 0.94 ;
 RECT 12.44 1.04 12.54 1.22 ;
 RECT 11.97 0.095 12.07 0.94 ;
 RECT 10.675 1.32 10.97 1.39 ;
 RECT 10.87 1.39 10.97 2.47 ;
 RECT 12.44 1.32 12.54 2.75 ;
 RECT 11.97 1.32 12.07 2.77 ;
 RECT 11.97 0.94 12.54 1.04 ;
 RECT 14.955 1.425 15.055 2.605 ;
 RECT 14.42 0.385 14.52 1.325 ;
 RECT 14.42 1.325 15.055 1.425 ;
 RECT 14.955 2.605 16.305 2.705 ;
 RECT 16.075 2.475 16.305 2.605 ;
 RECT 15.255 1.215 15.53 1.27 ;
 RECT 15.255 1.37 15.53 1.425 ;
 RECT 15.255 1.27 15.83 1.37 ;
 RECT 15.73 1.045 15.83 1.27 ;
 RECT 15.73 1.37 15.83 2.425 ;
 RECT 18.18 1.045 18.28 1.76 ;
 RECT 15.255 0.385 15.355 1.215 ;
 RECT 15.255 1.425 15.355 2.425 ;
 RECT 16.69 0.84 16.92 0.945 ;
 RECT 16.69 1.045 16.92 1.07 ;
 RECT 15.73 0.385 15.83 0.945 ;
 RECT 15.73 0.945 18.28 1.045 ;
 RECT 18.18 0.145 18.28 0.945 ;
 RECT 19.335 1.86 19.435 2.09 ;
 RECT 19.205 1.545 19.435 1.76 ;
 RECT 20.37 1.145 20.47 2.09 ;
 RECT 18.18 1.76 19.435 1.86 ;
 RECT 19.335 2.09 20.47 2.19 ;
 RECT 14.91 0.205 15.01 0.925 ;
 RECT 13.02 0.105 13.12 0.87 ;
 RECT 12.875 0.87 13.12 0.88 ;
 RECT 12.875 0.88 13.59 0.98 ;
 RECT 13.49 0.205 13.59 0.88 ;
 RECT 16.15 0.205 16.38 0.4 ;
 RECT 13.02 1.085 13.12 1.23 ;
 RECT 13.02 1.23 13.59 1.33 ;
 RECT 13.02 1.33 13.12 2.755 ;
 RECT 13.49 1.33 13.59 2.77 ;
 RECT 12.875 0.98 13.12 1.085 ;
 RECT 13.49 0.105 16.38 0.205 ;
 RECT 14.785 0.925 15.015 1.135 ;
 RECT 18.76 0.965 18.86 1.145 ;
 RECT 18.76 1.145 20.19 1.245 ;
 RECT 20.09 0.965 20.19 1.145 ;
 RECT 19.9 1.245 20 1.86 ;
 RECT 20.37 0.275 20.47 0.865 ;
 RECT 18.76 0.735 18.99 0.965 ;
 RECT 20.09 0.865 20.47 0.965 ;
 RECT 19.185 0.865 19.91 0.965 ;
 RECT 19.185 0.735 19.415 0.865 ;
 RECT 19.81 0.275 19.91 0.865 ;
 RECT 9.675 0.33 9.775 1.16 ;
 RECT 9.675 1.395 9.775 2.235 ;
 LAYER CO ;
 RECT 12.925 0.915 13.055 1.045 ;
 RECT 13.24 1.675 13.37 1.805 ;
 RECT 12.715 2.34 12.845 2.47 ;
 RECT 15.35 1.255 15.48 1.385 ;
 RECT 2.445 2.49 2.575 2.62 ;
 RECT 11.63 0.395 11.76 0.525 ;
 RECT 11.71 2.34 11.84 2.47 ;
 RECT 19.235 0.785 19.365 0.915 ;
 RECT 21.355 0.795 21.485 0.925 ;
 RECT 20.945 1.075 21.075 1.205 ;
 RECT 21.68 0.505 21.81 0.635 ;
 RECT 21.68 1.44 21.81 1.57 ;
 RECT 21.2 0.47 21.33 0.6 ;
 RECT 21.155 1.455 21.285 1.585 ;
 RECT 20.595 1.435 20.725 1.565 ;
 RECT 20.595 0.505 20.725 0.635 ;
 RECT 20.12 1.415 20.25 1.545 ;
 RECT 20.12 0.505 20.25 0.635 ;
 RECT 19.56 1.415 19.69 1.545 ;
 RECT 19.56 0.505 19.69 0.635 ;
 RECT 13.24 0.555 13.37 0.685 ;
 RECT 10.585 2.01 10.715 2.14 ;
 RECT 10.725 1.21 10.855 1.34 ;
 RECT 10.585 0.605 10.715 0.735 ;
 RECT 11.145 2.025 11.275 2.155 ;
 RECT 11.145 0.605 11.275 0.735 ;
 RECT 9.455 1.215 9.585 1.345 ;
 RECT 7.03 2.335 7.16 2.465 ;
 RECT 6.99 0.24 7.12 0.37 ;
 RECT 6.16 1.57 6.29 1.7 ;
 RECT 5.83 0.89 5.96 1.02 ;
 RECT 5.52 1.28 5.65 1.41 ;
 RECT 4.565 1.58 4.695 1.71 ;
 RECT 4.875 0.995 5.005 1.125 ;
 RECT 4.1 1.28 4.23 1.41 ;
 RECT 1.97 0.665 2.1 0.795 ;
 RECT 1.66 1.095 1.79 1.225 ;
 RECT 0.96 1.37 1.09 1.5 ;
 RECT 1.96 1.785 2.09 1.915 ;
 RECT 10.025 0.57 10.155 0.7 ;
 RECT 10.025 1.845 10.155 1.975 ;
 RECT 9.4 0.57 9.53 0.7 ;
 RECT 8.885 0.57 9.015 0.7 ;
 RECT 8.885 1.48 9.015 1.61 ;
 RECT 9.41 2.375 9.54 2.505 ;
 RECT 7.93 2.63 8.06 2.76 ;
 RECT 3.48 1.935 3.61 2.065 ;
 RECT 3.68 0.6 3.81 0.73 ;
 RECT 6.81 1.67 6.94 1.8 ;
 RECT 4.295 2.515 4.425 2.645 ;
 RECT 5.97 2.515 6.1 2.645 ;
 RECT 5.2 1.52 5.33 1.65 ;
 RECT 1.075 2.19 1.205 2.32 ;
 RECT 8.505 1.705 8.635 1.835 ;
 RECT 8.505 0.6 8.635 0.73 ;
 RECT 7.945 0.6 8.075 0.73 ;
 RECT 7.37 0.6 7.5 0.73 ;
 RECT 7.37 1.48 7.5 1.61 ;
 RECT 6.81 0.6 6.94 0.73 ;
 RECT 6 0.555 6.13 0.685 ;
 RECT 5.2 0.6 5.33 0.73 ;
 RECT 3.11 2.14 3.24 2.27 ;
 RECT 3.11 0.315 3.24 0.445 ;
 RECT 2.635 0.315 2.765 0.445 ;
 RECT 2.635 2.14 2.765 2.27 ;
 RECT 1.85 2.14 1.98 2.27 ;
 RECT 1.85 0.315 1.98 0.445 ;
 RECT 1.075 0.315 1.205 0.445 ;
 RECT 0.605 0.315 0.735 0.445 ;
 RECT 0.605 2.14 0.735 2.27 ;
 RECT 16.2 0.225 16.33 0.355 ;
 RECT 18.48 1.475 18.61 1.605 ;
 RECT 17.875 1.255 18.005 1.385 ;
 RECT 17.83 0.505 17.96 0.635 ;
 RECT 16.125 2.525 16.255 2.655 ;
 RECT 14.065 2.455 14.195 2.585 ;
 RECT 14.465 1.655 14.595 1.785 ;
 RECT 15.955 0.615 16.085 0.745 ;
 RECT 15.475 0.615 15.605 0.745 ;
 RECT 15.475 2.075 15.605 2.205 ;
 RECT 14.66 2.05 14.79 2.18 ;
 RECT 14.66 0.615 14.79 0.745 ;
 RECT 15.955 2.065 16.085 2.195 ;
 RECT 12.19 1.675 12.32 1.805 ;
 RECT 10.14 2.525 10.27 2.655 ;
 RECT 12.76 0.395 12.89 0.525 ;
 RECT 12.19 0.585 12.32 0.715 ;
 RECT 14.835 0.965 14.965 1.095 ;
 RECT 7.775 1.25 7.905 1.38 ;
 RECT 2.785 1.565 2.915 1.695 ;
 RECT 13.715 0.395 13.845 0.525 ;
 RECT 13.72 2.34 13.85 2.47 ;
 RECT 9.065 2.185 9.195 2.315 ;
 RECT 16.74 0.89 16.87 1.02 ;
 RECT 19.255 1.595 19.385 1.725 ;
 RECT 18.81 0.785 18.94 0.915 ;
 RECT 4.295 0.12 4.425 0.25 ;
 RECT 22.1 1.44 22.23 1.57 ;
 RECT 0.2 0.36 0.33 0.49 ;
 RECT 0.2 0.62 0.33 0.75 ;
 RECT 0.2 1.71 0.33 1.84 ;
 RECT 0.2 1.97 0.33 2.1 ;
 RECT 0.2 2.23 0.33 2.36 ;
 RECT 18.48 0.225 18.61 0.355 ;
 LAYER M1 ;
 RECT 15.255 1.17 15.595 1.51 ;
 RECT 5.195 0.55 5.335 1.275 ;
 RECT 4.05 1.275 5.335 1.415 ;
 RECT 5.195 1.415 5.335 1.71 ;
 RECT 7.365 0.55 7.505 1.475 ;
 RECT 7.3 1.475 7.57 1.615 ;
 RECT 11.905 0.385 12.045 0.88 ;
 RECT 11.14 0.88 12.045 1.02 ;
 RECT 11.14 0.55 11.28 0.88 ;
 RECT 11.14 1.02 11.28 2.21 ;
 RECT 12.465 0.385 12.605 0.75 ;
 RECT 11.905 0.245 12.605 0.385 ;
 RECT 12.92 0.89 13.06 1.095 ;
 RECT 12.465 0.75 13.06 0.89 ;
 RECT 2.305 0.45 2.445 1.56 ;
 RECT 2.305 1.7 2.445 2.135 ;
 RECT 1.78 0.31 2.445 0.45 ;
 RECT 1.78 2.135 2.445 2.275 ;
 RECT 2.735 1.525 2.965 1.56 ;
 RECT 2.735 1.7 2.965 1.735 ;
 RECT 2.305 1.56 2.965 1.7 ;
 RECT 21.675 0.435 21.815 1.07 ;
 RECT 20.875 1.07 21.815 1.21 ;
 RECT 21.675 1.21 21.815 1.64 ;
 RECT 0.6 0.275 0.74 0.31 ;
 RECT 0.6 0.45 0.74 1.86 ;
 RECT 0.6 2 0.74 2.365 ;
 RECT 0.555 0.31 0.785 0.45 ;
 RECT 1.36 2 1.5 2.52 ;
 RECT 0.6 1.86 1.5 2 ;
 RECT 1.36 2.52 2.625 2.66 ;
 RECT 2.395 2.45 2.625 2.52 ;
 RECT 15.095 1.845 15.235 2.45 ;
 RECT 14.06 2.385 14.2 2.45 ;
 RECT 14.06 2.45 15.235 2.59 ;
 RECT 14.06 2.59 14.2 2.65 ;
 RECT 15.95 0.55 16.09 1.705 ;
 RECT 15.095 1.705 16.09 1.845 ;
 RECT 15.95 1.845 16.09 2.265 ;
 RECT 7.725 1.21 7.955 1.245 ;
 RECT 7.725 1.385 7.955 1.42 ;
 RECT 7.725 1.245 8.64 1.385 ;
 RECT 8.5 0.55 8.64 1.245 ;
 RECT 8.5 1.385 8.64 1.9 ;
 RECT 14.785 0.925 15.015 0.955 ;
 RECT 14.46 0.955 15.015 1.095 ;
 RECT 14.785 1.095 15.015 1.135 ;
 RECT 14.46 1.095 14.6 1.835 ;
 RECT 3.77 1.13 3.91 2.42 ;
 RECT 3.105 0.275 3.245 0.31 ;
 RECT 3.105 0.45 3.245 2.42 ;
 RECT 3.105 2.42 3.91 2.56 ;
 RECT 3.06 0.31 3.29 0.45 ;
 RECT 3.77 0.99 5.055 1.13 ;
 RECT 17.87 0.64 18.01 0.78 ;
 RECT 17.87 0.92 18.01 1.455 ;
 RECT 17.765 0.5 18.01 0.64 ;
 RECT 17.87 0.78 19.005 0.92 ;
 RECT 19.25 0.92 19.39 1.785 ;
 RECT 19.165 0.78 19.415 0.92 ;
 RECT 10.86 1.775 11 2.435 ;
 RECT 11.42 2.135 11.56 2.435 ;
 RECT 10.3 1.635 11 1.775 ;
 RECT 10.86 2.435 11.56 2.575 ;
 RECT 10.3 1.775 10.44 2.52 ;
 RECT 10.07 2.52 10.44 2.66 ;
 RECT 13.515 1.86 13.655 1.995 ;
 RECT 11.42 1.995 13.655 2.135 ;
 RECT 14.175 0.75 14.315 1.72 ;
 RECT 14.175 2.045 14.84 2.185 ;
 RECT 14.175 1.86 14.315 2.045 ;
 RECT 13.515 1.72 14.315 1.86 ;
 RECT 14.175 0.61 14.86 0.75 ;
 RECT 18.15 0.36 18.29 0.5 ;
 RECT 16.1 0.22 18.29 0.36 ;
 RECT 19.555 0.435 19.695 0.5 ;
 RECT 19.555 0.64 19.695 1.61 ;
 RECT 18.15 0.5 19.695 0.64 ;
 RECT 6.325 0.375 6.465 1.26 ;
 RECT 7.655 0.375 7.795 0.93 ;
 RECT 6.155 1.26 6.465 1.4 ;
 RECT 6.155 1.4 6.295 1.77 ;
 RECT 6.325 0.235 7.795 0.375 ;
 RECT 8.22 0.38 8.36 0.93 ;
 RECT 8.88 0.38 9.02 1.66 ;
 RECT 8.22 0.24 9.02 0.38 ;
 RECT 7.655 0.93 8.36 1.07 ;
 RECT 16.045 2.52 18.29 2.66 ;
 RECT 18.15 1.33 18.29 2.52 ;
 RECT 20.59 0.64 20.73 1.925 ;
 RECT 18.8 1.33 18.94 1.925 ;
 RECT 20.525 0.5 20.775 0.64 ;
 RECT 18.8 1.925 20.73 2.065 ;
 RECT 18.15 1.19 18.94 1.33 ;
 RECT 8.78 1.94 8.92 2.05 ;
 RECT 7.02 2.05 8.92 2.19 ;
 RECT 7.02 1.805 7.16 2.05 ;
 RECT 6.805 0.545 6.945 1.665 ;
 RECT 6.735 1.665 7.16 1.805 ;
 RECT 10.3 0.365 10.44 1.205 ;
 RECT 9.74 0.365 9.88 1.8 ;
 RECT 9.74 0.225 10.44 0.365 ;
 RECT 8.78 1.8 9.88 1.94 ;
 RECT 10.3 1.205 10.925 1.345 ;
 RECT 6.69 2.085 6.83 2.33 ;
 RECT 4.555 1.945 6.83 2.085 ;
 RECT 5.825 0.835 5.965 1.945 ;
 RECT 4.56 1.715 4.7 1.945 ;
 RECT 4.49 1.575 4.765 1.715 ;
 RECT 9.06 2.23 9.2 2.33 ;
 RECT 6.69 2.33 9.2 2.47 ;
 RECT 9.06 2.09 10.16 2.23 ;
 RECT 10.02 0.52 10.16 2.09 ;
 RECT 20.915 0.36 21.055 0.79 ;
 RECT 20.115 0.36 20.255 1.41 ;
 RECT 20.115 0.22 21.055 0.36 ;
 RECT 20.05 1.41 20.32 1.55 ;
 RECT 20.915 0.79 21.535 0.93 ;
 RECT 3.475 0.6 3.88 0.735 ;
 RECT 3.475 0.735 3.615 2.13 ;
 RECT 4.755 0.41 4.895 0.46 ;
 RECT 4.755 0.275 5.655 0.41 ;
 RECT 5.515 0.41 5.655 1.475 ;
 RECT 4.755 0.27 5.59 0.275 ;
 RECT 3.475 0.595 4.895 0.6 ;
 RECT 3.68 0.46 4.895 0.595 ;
 RECT 4.755 0.6 4.895 0.61 ;
 END
END RSDFFNX2

MACRO ANTENNA
 CLASS CORE ANTENNACELL ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 1.6 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 1.6 2.96 ;
 RECT 1.06 1.92 1.2 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 1.6 0.08 ;
 RECT 1.085 0.08 1.225 0.76 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 1.16 0.47 1.4 ;
 RECT 0.33 1.4 0.47 1.715 ;
 RECT 0.33 0.74 0.47 1.16 ;
 END
 ANTENNADIFFAREA 0.526 ;
 END INP

 OBS
 LAYER CO ;
 RECT 1.065 1.97 1.195 2.1 ;
 RECT 1.09 0.575 1.22 0.705 ;
 RECT 1.09 0.315 1.22 0.445 ;
 RECT 0.335 0.79 0.465 0.92 ;
 RECT 0.335 1.535 0.465 1.665 ;
 RECT 1.065 2.23 1.195 2.36 ;
 END
END ANTENNA

MACRO AOBUFX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 5.76 ;
 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 2.31 1.62 2.45 1.76 ;
 RECT 2.365 2.15 2.505 2.66 ;
 RECT 2.265 1.9 2.585 2.15 ;
 RECT 1.9 1.76 2.585 1.9 ;
 RECT 1.9 1.625 2.04 1.76 ;
 END
 END VDDG

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.67 0.8 2.04 1.145 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END INP

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.895 4.36 2.36 4.6 ;
 RECT 1.895 4.6 2.035 5.27 ;
 RECT 1.895 3.65 2.035 4.36 ;
 END
 ANTENNADIFFAREA 0.483 ;
 END Z

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 2.31 0.08 2.45 0.765 ;
 RECT 1.9 0.08 2.04 0.53 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 3.84 5.84 ;
 RECT 1.425 5.19 1.565 5.68 ;
 RECT 2.31 4.975 2.45 5.68 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 2.32 2.425 2.785 3.37 ;
 RECT 1.525 2.415 1.78 2.645 ;
 RECT 1.68 2.645 1.78 5.665 ;
 RECT 1.68 0.1 1.78 0.845 ;
 RECT 1.68 0.845 1.94 1.075 ;
 RECT 1.68 1.075 1.78 2.185 ;
 LAYER CO ;
 RECT 2.315 5.31 2.445 5.44 ;
 RECT 2.315 5.035 2.445 5.165 ;
 RECT 2.37 2.47 2.5 2.6 ;
 RECT 2.37 3.19 2.5 3.32 ;
 RECT 1.575 2.465 1.705 2.595 ;
 RECT 1.9 5.075 2.03 5.205 ;
 RECT 1.43 5.26 1.56 5.39 ;
 RECT 1.43 3.375 1.56 3.505 ;
 RECT 1.9 3.715 2.03 3.845 ;
 RECT 1.9 4.015 2.03 4.145 ;
 RECT 1.905 0.33 2.035 0.46 ;
 RECT 1.905 1.695 2.035 1.825 ;
 RECT 1.76 0.895 1.89 1.025 ;
 RECT 1.43 1.685 1.56 1.815 ;
 RECT 1.43 0.33 1.56 0.46 ;
 RECT 2.315 0.305 2.445 0.435 ;
 RECT 2.315 0.565 2.445 0.695 ;
 RECT 2.315 1.69 2.445 1.82 ;
 RECT 2.315 1.95 2.445 2.08 ;
 LAYER M1 ;
 RECT 2.365 3.12 2.505 3.37 ;
 RECT 1.355 3.37 2.505 3.51 ;
 RECT 1.425 1.435 1.565 2.46 ;
 RECT 1.425 0.26 1.565 0.52 ;
 RECT 1.36 0.52 1.565 0.66 ;
 RECT 1.36 0.66 1.5 1.295 ;
 RECT 1.36 1.295 1.565 1.435 ;
 RECT 1.425 2.46 1.76 2.6 ;
 END
END AOBUFX1

MACRO AOBUFX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 5.76 ;
 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 2.31 1.62 2.45 1.76 ;
 RECT 2.365 2.465 3.135 2.605 ;
 RECT 2.265 1.9 2.585 2.15 ;
 RECT 2.365 2.15 2.505 2.465 ;
 RECT 1.9 1.76 2.585 1.9 ;
 RECT 1.9 1.625 2.04 1.76 ;
 END
 END VDDG

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.68 0.84 2.04 1.08 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END INP

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.895 4.6 2.035 5.27 ;
 RECT 1.895 4.36 2.36 4.6 ;
 RECT 1.895 3.695 2.035 4.36 ;
 END
 ANTENNADIFFAREA 0.616 ;
 END Z

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 2.31 0.08 2.45 0.765 ;
 RECT 1.9 0.08 2.04 0.53 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 3.84 5.84 ;
 RECT 1.425 5.19 1.565 5.68 ;
 RECT 2.37 5.185 2.51 5.68 ;
 RECT 0.855 4.905 0.995 5.68 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 2.89 2.425 3.48 3.37 ;
 RECT 1.68 2.645 1.78 4.715 ;
 RECT 1.68 4.815 1.78 5.665 ;
 RECT 1.68 4.715 2.25 4.815 ;
 RECT 2.15 3.005 2.25 4.715 ;
 RECT 2.15 4.815 2.25 5.665 ;
 RECT 1.525 2.415 1.78 2.645 ;
 RECT 1.68 0.1 1.78 0.845 ;
 RECT 1.68 1.075 1.78 2.235 ;
 RECT 1.68 0.845 1.91 1.075 ;
 LAYER CO ;
 RECT 0.86 4.975 0.99 5.105 ;
 RECT 0.86 5.235 0.99 5.365 ;
 RECT 2.375 5.255 2.505 5.385 ;
 RECT 2.375 3.89 2.505 4.02 ;
 RECT 1.43 3.74 1.56 3.87 ;
 RECT 1.43 4.105 1.56 4.235 ;
 RECT 2.375 3.375 2.505 3.505 ;
 RECT 2.94 2.47 3.07 2.6 ;
 RECT 2.94 3.19 3.07 3.32 ;
 RECT 1.575 2.465 1.705 2.595 ;
 RECT 1.9 5.075 2.03 5.205 ;
 RECT 1.43 5.27 1.56 5.4 ;
 RECT 1.43 3.375 1.56 3.505 ;
 RECT 1.9 3.77 2.03 3.9 ;
 RECT 1.9 4.07 2.03 4.2 ;
 RECT 1.905 0.33 2.035 0.46 ;
 RECT 1.905 1.695 2.035 1.825 ;
 RECT 1.73 0.895 1.86 1.025 ;
 RECT 1.43 1.685 1.56 1.815 ;
 RECT 1.43 0.33 1.56 0.46 ;
 RECT 2.315 0.305 2.445 0.435 ;
 RECT 2.315 0.565 2.445 0.695 ;
 RECT 2.315 1.69 2.445 1.82 ;
 RECT 2.315 1.95 2.445 2.08 ;
 LAYER M1 ;
 RECT 1.425 3.51 1.565 4.315 ;
 RECT 2.37 3.51 2.51 4.09 ;
 RECT 2.935 3.12 3.075 3.37 ;
 RECT 1.355 3.37 3.075 3.51 ;
 RECT 1.425 1.435 1.565 2.46 ;
 RECT 1.425 0.26 1.565 0.52 ;
 RECT 1.36 0.52 1.565 0.66 ;
 RECT 1.36 0.66 1.5 1.295 ;
 RECT 1.36 1.295 1.565 1.435 ;
 RECT 1.425 2.46 1.76 2.6 ;
 END
END AOBUFX2

MACRO AOBUFX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 5.76 ;
 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 2.31 1.62 2.45 1.69 ;
 RECT 2.365 2.465 3.855 2.605 ;
 RECT 2.265 1.83 2.585 2.15 ;
 RECT 2.365 2.15 2.505 2.465 ;
 RECT 1.9 1.69 2.585 1.83 ;
 RECT 1.9 1.83 2.04 1.9 ;
 RECT 1.9 1.625 2.04 1.69 ;
 END
 END VDDG

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.68 0.84 2.04 1.08 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END INP

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 2.31 0.08 2.45 0.765 ;
 RECT 1.9 0.08 2.04 0.53 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 4.8 5.84 ;
 RECT 1.425 5.19 1.565 5.68 ;
 RECT 0.855 4.905 0.995 5.68 ;
 RECT 2.365 5.19 2.505 5.68 ;
 RECT 3.31 5.185 3.45 5.68 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 END
 END VDD

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.835 3.695 2.975 4.36 ;
 RECT 2.835 4.36 3.325 4.54 ;
 RECT 1.895 4.54 3.325 4.6 ;
 RECT 1.895 4.68 2.035 5.27 ;
 RECT 1.895 4.6 2.975 4.68 ;
 RECT 2.835 4.68 2.975 5.27 ;
 RECT 1.895 3.695 2.035 4.54 ;
 END
 ANTENNADIFFAREA 1.128 ;
 END Z

 OBS
 LAYER PO ;
 RECT 3.625 2.425 4.14 3.37 ;
 RECT 2.62 2.635 2.72 4.715 ;
 RECT 1.68 2.645 1.78 4.715 ;
 RECT 1.68 4.815 1.78 5.665 ;
 RECT 1.68 4.715 2.25 4.815 ;
 RECT 3.09 3.005 3.19 4.715 ;
 RECT 3.09 4.815 3.19 5.665 ;
 RECT 2.62 4.715 3.19 4.815 ;
 RECT 2.62 4.815 2.72 5.665 ;
 RECT 1.525 2.415 1.78 2.535 ;
 RECT 1.525 2.535 2.72 2.635 ;
 RECT 1.525 2.635 1.78 2.645 ;
 RECT 2.15 3.005 2.25 4.715 ;
 RECT 2.15 4.815 2.25 5.665 ;
 RECT 1.68 0.1 1.78 0.845 ;
 RECT 1.68 1.075 1.78 2.235 ;
 RECT 1.68 0.845 1.91 1.075 ;
 LAYER CO ;
 RECT 3.315 3.89 3.445 4.02 ;
 RECT 3.315 3.375 3.445 3.505 ;
 RECT 2.84 5.075 2.97 5.205 ;
 RECT 2.37 5.27 2.5 5.4 ;
 RECT 2.84 3.77 2.97 3.9 ;
 RECT 3.315 5.255 3.445 5.385 ;
 RECT 2.84 4.07 2.97 4.2 ;
 RECT 0.86 4.975 0.99 5.105 ;
 RECT 0.86 5.235 0.99 5.365 ;
 RECT 2.37 3.89 2.5 4.02 ;
 RECT 1.43 3.74 1.56 3.87 ;
 RECT 1.43 4.105 1.56 4.235 ;
 RECT 2.37 3.375 2.5 3.505 ;
 RECT 3.675 2.47 3.805 2.6 ;
 RECT 3.675 3.19 3.805 3.32 ;
 RECT 1.575 2.465 1.705 2.595 ;
 RECT 1.9 5.075 2.03 5.205 ;
 RECT 1.43 5.27 1.56 5.4 ;
 RECT 1.43 3.375 1.56 3.505 ;
 RECT 1.9 3.77 2.03 3.9 ;
 RECT 1.9 4.07 2.03 4.2 ;
 RECT 1.905 0.33 2.035 0.46 ;
 RECT 1.905 1.695 2.035 1.825 ;
 RECT 1.73 0.895 1.86 1.025 ;
 RECT 1.43 1.685 1.56 1.815 ;
 RECT 1.43 0.33 1.56 0.46 ;
 RECT 2.315 0.305 2.445 0.435 ;
 RECT 2.315 0.565 2.445 0.695 ;
 RECT 2.315 1.69 2.445 1.82 ;
 RECT 2.315 1.95 2.445 2.08 ;
 LAYER M1 ;
 RECT 2.365 3.51 2.505 4.09 ;
 RECT 1.425 3.51 1.565 4.315 ;
 RECT 1.355 3.37 3.81 3.51 ;
 RECT 3.31 3.51 3.45 4.09 ;
 RECT 3.67 3.12 3.81 3.37 ;
 RECT 1.425 1.435 1.565 2.46 ;
 RECT 1.425 0.26 1.565 0.52 ;
 RECT 1.36 0.52 1.565 0.66 ;
 RECT 1.36 0.66 1.5 1.295 ;
 RECT 1.36 1.295 1.565 1.435 ;
 RECT 1.425 2.46 1.76 2.6 ;
 END
END AOBUFX4

MACRO RDFFSRSSRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 28.48 BY 2.88 ;
 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.76 1.16 10.055 1.505 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 21.725 0.59 22.095 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.45 1.255 17.69 1.495 ;
 RECT 17.55 0.915 17.69 1.255 ;
 RECT 17.55 1.7 18.685 1.84 ;
 RECT 17.55 1.84 17.69 1.9 ;
 RECT 17.55 1.495 17.69 1.7 ;
 RECT 18.545 1.84 18.685 1.9 ;
 RECT 18.545 0.915 18.685 1.7 ;
 END
 ANTENNADIFFAREA 0.961 ;
 END Q

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.2 1.475 4.53 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.08 1.135 19.335 1.375 ;
 RECT 19.195 0.55 19.335 1.135 ;
 RECT 20.255 1.905 20.395 1.91 ;
 RECT 19.195 1.765 20.395 1.905 ;
 RECT 20.255 0.56 20.395 1.765 ;
 RECT 19.195 1.905 19.335 1.915 ;
 RECT 19.195 1.375 19.335 1.765 ;
 END
 ANTENNADIFFAREA 0.725 ;
 END QN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 28.48 0.08 ;
 RECT 25.395 0.08 25.635 0.26 ;
 RECT 10.305 0.59 10.58 0.73 ;
 RECT 17.985 0.335 18.25 0.495 ;
 RECT 1.345 0.08 1.645 0.26 ;
 RECT 0.35 0.08 0.49 0.775 ;
 RECT 4.15 0.08 4.29 1.055 ;
 RECT 4.895 0.08 5.035 0.39 ;
 RECT 7.495 0.08 7.73 0.595 ;
 RECT 14.23 0.08 14.37 0.945 ;
 RECT 15.735 0.08 15.875 0.525 ;
 RECT 23.045 0.08 23.185 0.36 ;
 RECT 19.755 0.08 19.895 0.82 ;
 RECT 24.26 0.08 24.4 0.35 ;
 RECT 10.37 0.08 10.51 0.59 ;
 RECT 18.04 0.08 18.18 0.335 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 28.48 2.96 ;
 RECT 0.41 1.74 0.55 2.8 ;
 RECT 1.45 1.98 1.59 2.8 ;
 RECT 4.825 2.34 5.075 2.8 ;
 RECT 4.15 1.98 4.29 2.8 ;
 RECT 10.18 2.375 10.32 2.8 ;
 RECT 8.08 2.07 8.22 2.8 ;
 RECT 14.83 2.57 14.97 2.8 ;
 RECT 17.955 2.57 18.095 2.8 ;
 RECT 19.67 2.57 19.81 2.8 ;
 RECT 15.73 2.57 15.87 2.8 ;
 RECT 15.19 2.54 15.42 2.8 ;
 END
 END VDD

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.955 1.435 27.295 1.8 ;
 RECT 25.275 1.99 27.14 2.13 ;
 RECT 23.045 2.22 25.415 2.36 ;
 RECT 25.275 1.435 25.415 1.99 ;
 RECT 27 1.8 27.14 1.99 ;
 RECT 23.045 1.39 23.185 2.22 ;
 RECT 24.43 1.37 24.57 2.22 ;
 RECT 25.275 2.13 25.415 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.06 1.455 2.44 1.735 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.43 0.22 3.73 0.535 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.165 1.48 1.48 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SETB

 OBS
 LAYER PO ;
 RECT 14.615 0.47 14.78 0.625 ;
 RECT 13.76 0.455 14.78 0.47 ;
 RECT 13.76 0.47 13.99 0.665 ;
 RECT 13.84 0.37 14.78 0.455 ;
 RECT 14.615 0.625 14.845 0.835 ;
 RECT 22.83 0.21 22.93 0.755 ;
 RECT 22.83 0.855 22.93 2.2 ;
 RECT 25.695 1.125 25.795 2.2 ;
 RECT 21.865 0.755 23.4 0.84 ;
 RECT 21.865 0.84 23.395 0.855 ;
 RECT 23.3 0.215 23.4 0.755 ;
 RECT 21.865 0.595 22.095 0.755 ;
 RECT 22.83 2.2 25.795 2.3 ;
 RECT 20.035 0.32 20.135 1.33 ;
 RECT 19.44 1.2 19.65 1.33 ;
 RECT 19.44 1.43 19.65 1.435 ;
 RECT 19.44 1.33 20.135 1.43 ;
 RECT 19.455 0.4 19.555 1.2 ;
 RECT 19.455 1.435 19.555 2.585 ;
 RECT 20.035 1.43 20.135 2.58 ;
 RECT 21.285 0.32 21.515 0.43 ;
 RECT 20.035 0.22 21.515 0.32 ;
 RECT 11.025 2.69 12.935 2.695 ;
 RECT 12.835 2.54 12.935 2.69 ;
 RECT 11.815 2.695 12.935 2.79 ;
 RECT 11.025 0.655 11.125 2.595 ;
 RECT 11.025 2.595 11.915 2.69 ;
 RECT 12.835 2.33 13.065 2.54 ;
 RECT 26.705 0.195 26.805 2.665 ;
 RECT 25.695 0.095 26.805 0.195 ;
 RECT 22.07 1.245 22.17 2.665 ;
 RECT 22.07 1.2 22.355 1.245 ;
 RECT 25.695 0.195 25.795 0.945 ;
 RECT 22.125 1.035 22.355 1.1 ;
 RECT 22.07 2.665 26.805 2.765 ;
 RECT 22.07 1.1 22.4 1.2 ;
 RECT 8.81 1.575 8.91 2.485 ;
 RECT 9.32 1.41 9.55 1.475 ;
 RECT 9.32 1.575 9.55 1.62 ;
 RECT 8.81 1.475 9.55 1.575 ;
 RECT 26.005 2.27 26.29 2.48 ;
 RECT 26.005 1.2 26.105 2.27 ;
 RECT 26.005 0.375 26.105 0.99 ;
 RECT 26.005 0.99 26.255 1.2 ;
 RECT 23.305 1.245 23.405 2.02 ;
 RECT 23.175 1.035 23.405 1.245 ;
 RECT 24.52 0.38 24.62 0.96 ;
 RECT 24.52 1.06 24.62 1.14 ;
 RECT 24.885 0.22 25.115 0.28 ;
 RECT 24.52 0.28 25.115 0.38 ;
 RECT 24.885 0.38 25.115 0.43 ;
 RECT 24.52 1.14 24.79 1.24 ;
 RECT 24.69 1.24 24.79 1.84 ;
 RECT 24.1 0.935 24.33 0.96 ;
 RECT 24.1 1.06 24.33 1.145 ;
 RECT 24.1 0.96 24.62 1.06 ;
 RECT 15.985 1.635 16.085 1.66 ;
 RECT 15.985 1.66 16.24 1.87 ;
 RECT 15.985 1.87 16.085 2.565 ;
 RECT 13.035 0.795 13.2 0.925 ;
 RECT 12.355 0.885 12.585 0.925 ;
 RECT 12.355 1.025 12.585 1.095 ;
 RECT 12.355 0.925 13.2 1.025 ;
 RECT 13.035 0.585 13.265 0.795 ;
 RECT 10.63 0.655 10.73 1.24 ;
 RECT 10.5 1.24 10.73 1.475 ;
 RECT 7.005 0.695 7.105 1.61 ;
 RECT 7.04 1.71 7.14 2.48 ;
 RECT 7.005 1.61 7.14 1.71 ;
 RECT 6.885 0.465 7.125 0.695 ;
 RECT 8.17 1.61 8.435 1.82 ;
 RECT 8.335 1.82 8.435 2.49 ;
 RECT 7.965 0.66 8.065 1.51 ;
 RECT 7.965 1.51 8.435 1.61 ;
 RECT 6.565 1.33 6.705 1.475 ;
 RECT 6.565 1.71 6.665 2.475 ;
 RECT 6.605 0.65 6.705 1.33 ;
 RECT 6.565 1.475 6.795 1.71 ;
 RECT 4.75 1.52 5.35 1.62 ;
 RECT 6.115 0.47 6.4 0.705 ;
 RECT 6.115 0.705 6.215 1.165 ;
 RECT 5.185 1.62 5.285 2.69 ;
 RECT 7.865 1.79 7.965 2.69 ;
 RECT 5.25 0.585 5.35 1.165 ;
 RECT 5.25 1.265 5.35 1.52 ;
 RECT 4.75 1.44 4.995 1.52 ;
 RECT 4.75 1.62 4.995 1.69 ;
 RECT 5.185 2.69 7.965 2.79 ;
 RECT 5.25 1.165 6.215 1.265 ;
 RECT 2.175 0.745 2.275 1.475 ;
 RECT 2.175 1.71 2.275 2.465 ;
 RECT 2.13 1.475 2.36 1.71 ;
 RECT 1.705 1.775 1.805 2.675 ;
 RECT 0.79 2.375 1.02 2.675 ;
 RECT 0.79 2.675 1.805 2.775 ;
 RECT 2.645 0.745 2.745 1.28 ;
 RECT 2.645 1.28 3.155 1.515 ;
 RECT 1.235 0.74 1.335 1.485 ;
 RECT 1.235 1.72 1.335 2.465 ;
 RECT 1.2 1.485 1.43 1.72 ;
 RECT 4.41 0.655 4.51 1.495 ;
 RECT 4.215 1.495 4.51 1.745 ;
 RECT 4.41 1.745 4.51 2.37 ;
 RECT 6.07 1.595 6.17 2.48 ;
 RECT 5.53 1.445 5.775 1.495 ;
 RECT 5.53 1.495 6.17 1.595 ;
 RECT 5.53 1.595 5.775 1.69 ;
 RECT 3.34 0.23 3.44 0.295 ;
 RECT 3.34 0.295 3.695 0.465 ;
 RECT 1.705 0.465 3.695 0.505 ;
 RECT 1.705 0.505 3.44 0.565 ;
 RECT 1.705 0.565 1.805 1.325 ;
 RECT 3.34 0.565 3.44 1.71 ;
 RECT 2.645 1.81 2.745 2.465 ;
 RECT 2.645 1.71 3.44 1.81 ;
 RECT 3.935 0.27 4.035 2.4 ;
 RECT 3.78 2.4 4.035 2.61 ;
 RECT 17.815 0.39 17.915 1.17 ;
 RECT 17.815 1.27 17.915 2.375 ;
 RECT 18.33 0.38 18.43 1.17 ;
 RECT 18.33 1.27 18.43 2.375 ;
 RECT 16.565 0.225 16.795 0.29 ;
 RECT 16.565 0.39 16.795 0.435 ;
 RECT 16.565 0.29 17.915 0.39 ;
 RECT 17.815 1.17 18.43 1.27 ;
 RECT 16.26 1.25 16.52 1.3 ;
 RECT 16.42 0.61 16.52 1.25 ;
 RECT 16.26 1.4 16.52 1.46 ;
 RECT 16.42 1.46 16.52 2.56 ;
 RECT 16.95 0.84 17.05 1.3 ;
 RECT 16.26 1.3 17.05 1.4 ;
 RECT 16.935 0.63 17.165 0.84 ;
 RECT 12.06 0.19 12.16 1.29 ;
 RECT 5.57 0.185 12.16 0.19 ;
 RECT 12.955 1.39 13.15 1.405 ;
 RECT 5.57 0.285 5.67 0.51 ;
 RECT 5.57 0.19 7.405 0.285 ;
 RECT 7.305 0.285 7.405 1.24 ;
 RECT 7.305 0.09 12.16 0.185 ;
 RECT 12.06 1.29 13.15 1.39 ;
 RECT 5.53 0.51 5.775 0.755 ;
 RECT 12.955 1.405 13.185 1.615 ;
 RECT 15.085 0.81 15.185 2.54 ;
 RECT 15.085 2.54 15.42 2.75 ;
 RECT 15.045 0.6 15.275 0.81 ;
 RECT 9.735 1.45 9.835 1.655 ;
 RECT 9.735 1.755 9.835 2.57 ;
 RECT 9.735 1.655 10.695 1.755 ;
 RECT 10.595 1.755 10.695 2.355 ;
 RECT 9.735 0.655 9.835 1.13 ;
 RECT 9.735 1.23 9.835 1.24 ;
 RECT 8.82 0.66 8.92 1.13 ;
 RECT 9.735 1.24 9.99 1.45 ;
 RECT 8.82 1.13 9.835 1.23 ;
 RECT 23.61 0.215 23.71 0.995 ;
 RECT 23.61 0.995 23.85 1.205 ;
 RECT 23.61 1.205 23.71 2 ;
 RECT 8.355 0.47 8.54 0.5 ;
 RECT 15.99 0.19 16.09 1.18 ;
 RECT 13.45 0.19 13.55 1.91 ;
 RECT 12.63 1.71 12.73 1.91 ;
 RECT 11.545 0.47 11.645 1.61 ;
 RECT 11.545 1.61 12.73 1.71 ;
 RECT 11.545 1.71 11.645 1.725 ;
 RECT 12.095 1.71 12.195 2.445 ;
 RECT 13.45 0.09 16.09 0.19 ;
 RECT 12.63 1.91 13.55 2.01 ;
 RECT 8.355 0.37 11.645 0.47 ;
 RECT 8.31 0.5 8.54 0.71 ;
 RECT 14.615 0.835 14.715 2.21 ;
 LAYER CO ;
 RECT 16.615 0.265 16.745 0.395 ;
 RECT 26.11 2.31 26.24 2.44 ;
 RECT 16.31 1.29 16.44 1.42 ;
 RECT 13.005 1.445 13.135 1.575 ;
 RECT 15.095 0.64 15.225 0.77 ;
 RECT 14.665 0.665 14.795 0.795 ;
 RECT 9.81 1.28 9.94 1.41 ;
 RECT 23.67 1.035 23.8 1.165 ;
 RECT 8.36 0.54 8.49 0.67 ;
 RECT 13.81 0.495 13.94 0.625 ;
 RECT 21.915 0.635 22.045 0.765 ;
 RECT 21.335 0.26 21.465 0.39 ;
 RECT 12.885 2.37 13.015 2.5 ;
 RECT 22.175 1.075 22.305 1.205 ;
 RECT 9.37 1.45 9.5 1.58 ;
 RECT 26.075 1.03 26.205 1.16 ;
 RECT 23.225 1.075 23.355 1.205 ;
 RECT 13.085 0.625 13.215 0.755 ;
 RECT 24.15 0.975 24.28 1.105 ;
 RECT 16.06 1.7 16.19 1.83 ;
 RECT 12.405 0.925 12.535 1.055 ;
 RECT 24.435 1.445 24.565 1.575 ;
 RECT 23.83 0.435 23.96 0.565 ;
 RECT 11.81 1.9 11.94 2.03 ;
 RECT 4.76 0.875 4.89 1.005 ;
 RECT 9.485 1.995 9.615 2.125 ;
 RECT 17.555 1.705 17.685 1.835 ;
 RECT 10.375 0.595 10.505 0.725 ;
 RECT 7.615 2.125 7.745 2.255 ;
 RECT 19.2 0.62 19.33 0.75 ;
 RECT 6.615 1.525 6.745 1.655 ;
 RECT 27.005 1.475 27.135 1.605 ;
 RECT 11.285 0.875 11.415 1.005 ;
 RECT 24.265 0.12 24.395 0.25 ;
 RECT 18.55 1.705 18.68 1.835 ;
 RECT 20.26 1.71 20.39 1.84 ;
 RECT 7.545 0.455 7.675 0.585 ;
 RECT 14.235 0.745 14.365 0.875 ;
 RECT 5.82 2.105 5.95 2.235 ;
 RECT 17.555 0.975 17.685 1.105 ;
 RECT 12.315 0.595 12.445 0.725 ;
 RECT 19.48 1.25 19.61 1.38 ;
 RECT 25.28 1.49 25.41 1.62 ;
 RECT 9.04 2.07 9.17 2.2 ;
 RECT 7.265 1.825 7.395 1.955 ;
 RECT 16.64 0.83 16.77 0.96 ;
 RECT 8.555 0.93 8.685 1.06 ;
 RECT 0.355 0.56 0.485 0.69 ;
 RECT 5.405 1.825 5.535 1.955 ;
 RECT 23.83 1.485 23.96 1.615 ;
 RECT 10.55 1.28 10.68 1.41 ;
 RECT 3.685 2.115 3.815 2.245 ;
 RECT 18.045 0.36 18.175 0.49 ;
 RECT 14.835 2.64 14.965 2.77 ;
 RECT 12.315 1.87 12.445 2 ;
 RECT 9.485 0.88 9.615 1.01 ;
 RECT 6.94 0.515 7.07 0.645 ;
 RECT 0.415 1.825 0.545 1.955 ;
 RECT 0.415 2.085 0.545 2.215 ;
 RECT 0.415 2.345 0.545 2.475 ;
 RECT 1.925 0.97 2.055 1.1 ;
 RECT 4.9 0.21 5.03 0.34 ;
 RECT 22.58 1.425 22.71 1.555 ;
 RECT 0.355 0.3 0.485 0.43 ;
 RECT 18.55 0.975 18.68 1.105 ;
 RECT 11.285 1.945 11.415 2.075 ;
 RECT 20.26 0.63 20.39 0.76 ;
 RECT 6.785 2.125 6.915 2.255 ;
 RECT 24.91 1.405 25.04 1.535 ;
 RECT 14.365 1.7 14.495 1.83 ;
 RECT 22.33 0.505 22.46 0.635 ;
 RECT 4.895 2.345 5.025 2.475 ;
 RECT 3.685 0.875 3.815 1.005 ;
 RECT 10.185 2.445 10.315 2.575 ;
 RECT 6.335 0.88 6.465 1.01 ;
 RECT 5.585 1.49 5.715 1.62 ;
 RECT 24.77 0.595 24.9 0.725 ;
 RECT 6.315 2.07 6.445 2.2 ;
 RECT 26.225 1.465 26.355 1.595 ;
 RECT 17.96 2.64 18.09 2.77 ;
 RECT 23.05 1.475 23.18 1.605 ;
 RECT 19.2 1.725 19.33 1.855 ;
 RECT 4.155 2.05 4.285 2.18 ;
 RECT 6.22 0.525 6.35 0.655 ;
 RECT 15.34 0.96 15.47 1.09 ;
 RECT 11.81 0.595 11.94 0.725 ;
 RECT 8.085 2.135 8.215 2.265 ;
 RECT 19.76 0.62 19.89 0.75 ;
 RECT 4.155 0.875 4.285 1.005 ;
 RECT 25.445 0.12 25.575 0.25 ;
 RECT 8.225 1.63 8.355 1.76 ;
 RECT 4.81 1.495 4.94 1.625 ;
 RECT 26.225 0.595 26.355 0.725 ;
 RECT 15.305 1.705 15.435 1.835 ;
 RECT 9.04 0.88 9.17 1.01 ;
 RECT 4.63 1.995 4.76 2.125 ;
 RECT 5.47 0.905 5.6 1.035 ;
 RECT 15.735 2.64 15.865 2.77 ;
 RECT 19.675 2.64 19.805 2.77 ;
 RECT 5.865 0.88 5.995 1.01 ;
 RECT 1.925 2.05 2.055 2.18 ;
 RECT 2.975 1.335 3.105 1.465 ;
 RECT 2.18 1.53 2.31 1.66 ;
 RECT 0.985 2.05 1.115 2.18 ;
 RECT 0.985 0.97 1.115 1.1 ;
 RECT 1.455 2.05 1.585 2.18 ;
 RECT 2.865 0.97 2.995 1.1 ;
 RECT 1.25 1.54 1.38 1.67 ;
 RECT 2.395 2.05 2.525 2.18 ;
 RECT 0.84 2.43 0.97 2.56 ;
 RECT 2.865 2.05 2.995 2.18 ;
 RECT 2.395 0.97 2.525 1.1 ;
 RECT 1.465 0.125 1.595 0.255 ;
 RECT 15.74 0.33 15.87 0.46 ;
 RECT 8.555 2.015 8.685 2.145 ;
 RECT 4.275 1.55 4.405 1.68 ;
 RECT 16.64 1.78 16.77 1.91 ;
 RECT 23.05 0.135 23.18 0.265 ;
 RECT 5.585 0.555 5.715 0.685 ;
 RECT 3.515 0.335 3.645 0.465 ;
 RECT 3.83 2.44 3.96 2.57 ;
 RECT 15.24 2.58 15.37 2.71 ;
 RECT 16.985 0.67 17.115 0.8 ;
 RECT 24.935 0.26 25.065 0.39 ;
 LAYER M1 ;
 RECT 24.7 0.59 24.975 0.73 ;
 RECT 26.025 0.99 26.255 1.04 ;
 RECT 24.765 1.04 26.255 1.18 ;
 RECT 26.025 1.18 26.255 1.2 ;
 RECT 24.885 0.29 25.255 0.43 ;
 RECT 25.115 0.43 25.255 0.71 ;
 RECT 24.885 0.22 25.115 0.29 ;
 RECT 26.535 0.85 26.675 1.385 ;
 RECT 26.22 1.525 26.36 1.73 ;
 RECT 25.115 0.71 26.675 0.85 ;
 RECT 26.22 0.51 26.36 0.71 ;
 RECT 26.22 1.385 26.675 1.525 ;
 RECT 22.125 1.225 22.355 1.245 ;
 RECT 22.125 1.195 22.715 1.225 ;
 RECT 22.265 1.015 22.575 1.035 ;
 RECT 22.125 1.035 22.575 1.055 ;
 RECT 22.4 0.64 22.54 1.015 ;
 RECT 22.575 1.225 22.715 1.75 ;
 RECT 22.28 0.5 22.54 0.64 ;
 RECT 23.175 1.035 23.405 1.055 ;
 RECT 23.175 1.195 23.405 1.245 ;
 RECT 22.125 1.055 23.405 1.195 ;
 RECT 24.145 1.145 24.285 1.345 ;
 RECT 23.825 1.485 23.965 1.76 ;
 RECT 24.145 0.73 24.285 0.935 ;
 RECT 23.825 0.355 23.965 0.59 ;
 RECT 23.825 1.345 24.285 1.485 ;
 RECT 24.1 0.935 24.33 1.145 ;
 RECT 23.825 0.59 24.285 0.73 ;
 RECT 21.285 0.36 21.515 0.43 ;
 RECT 22.68 0.36 22.82 0.565 ;
 RECT 21.285 0.22 22.82 0.36 ;
 RECT 23.42 0.705 23.56 0.75 ;
 RECT 23.545 0.995 23.85 1.205 ;
 RECT 23.545 0.89 23.685 0.995 ;
 RECT 23.42 0.75 23.685 0.89 ;
 RECT 22.68 0.565 23.56 0.705 ;
 RECT 16.935 0.63 17.165 0.635 ;
 RECT 16.935 0.775 17.165 0.84 ;
 RECT 18.45 0.37 18.59 0.635 ;
 RECT 16.93 0.635 18.59 0.775 ;
 RECT 19.475 0.37 19.615 1.46 ;
 RECT 18.445 0.23 19.615 0.37 ;
 RECT 9.035 0.82 9.175 2.33 ;
 RECT 9.035 2.47 9.175 2.475 ;
 RECT 9.885 2.165 10.025 2.33 ;
 RECT 9.885 2.47 10.025 2.475 ;
 RECT 9.035 2.33 10.025 2.47 ;
 RECT 10.965 2.165 11.105 2.295 ;
 RECT 11.28 0.765 11.42 2.295 ;
 RECT 11.28 2.435 11.42 2.44 ;
 RECT 11.805 0.525 11.945 2.295 ;
 RECT 11.805 2.435 11.945 2.44 ;
 RECT 9.885 2.025 11.105 2.165 ;
 RECT 10.965 2.295 11.945 2.435 ;
 RECT 12.31 0.525 12.45 0.885 ;
 RECT 12.31 1.095 12.45 2.065 ;
 RECT 12.31 0.885 12.585 1.095 ;
 RECT 15.415 0.36 15.555 0.665 ;
 RECT 14.615 0.22 15.56 0.36 ;
 RECT 14.615 0.36 14.845 0.835 ;
 RECT 16.635 0.22 16.775 0.225 ;
 RECT 16.635 0.435 16.775 0.665 ;
 RECT 15.415 0.665 16.775 0.805 ;
 RECT 16.635 0.805 16.775 1.98 ;
 RECT 16.565 0.225 16.795 0.435 ;
 RECT 13.76 0.455 13.99 0.49 ;
 RECT 13.035 0.49 13.99 0.63 ;
 RECT 13.76 0.63 13.99 0.665 ;
 RECT 13.035 0.63 13.265 0.795 ;
 RECT 9.365 0.36 9.505 0.525 ;
 RECT 7.87 0.36 8.01 0.735 ;
 RECT 7.87 0.22 9.505 0.36 ;
 RECT 6.935 0.735 8.01 0.875 ;
 RECT 6.935 0.695 7.125 0.735 ;
 RECT 6.935 0.445 7.075 0.465 ;
 RECT 6.9 0.465 7.125 0.695 ;
 RECT 10.745 0.385 10.885 0.87 ;
 RECT 12.755 0.385 12.895 1.09 ;
 RECT 10.745 0.255 12.895 0.385 ;
 RECT 10.745 0.245 12.89 0.255 ;
 RECT 10.025 0.87 10.885 1.01 ;
 RECT 10.745 1.01 10.885 1.015 ;
 RECT 10.025 0.665 10.165 0.87 ;
 RECT 9.365 0.525 10.165 0.665 ;
 RECT 14.985 0.6 15.275 0.81 ;
 RECT 14.985 0.81 15.125 1.09 ;
 RECT 12.755 1.09 15.125 1.23 ;
 RECT 5.465 0.5 5.72 0.965 ;
 RECT 5.465 1.67 5.605 1.82 ;
 RECT 5.465 1.96 5.605 2.65 ;
 RECT 5.465 0.965 5.605 1.44 ;
 RECT 5.465 1.44 5.72 1.67 ;
 RECT 5.335 1.82 5.605 1.96 ;
 RECT 6.15 0.52 6.75 0.66 ;
 RECT 6.61 0.66 6.75 1.015 ;
 RECT 8.155 0.505 8.54 0.71 ;
 RECT 8.31 0.5 8.54 0.505 ;
 RECT 8.155 0.71 8.295 1.015 ;
 RECT 6.61 1.015 8.295 1.155 ;
 RECT 3.46 1.01 3.6 1.195 ;
 RECT 3.46 1.335 3.6 2.11 ;
 RECT 3.46 2.25 3.6 2.255 ;
 RECT 3.46 0.87 3.885 1.01 ;
 RECT 3.46 2.11 3.885 2.25 ;
 RECT 4.43 0.67 4.57 1.195 ;
 RECT 3.46 1.195 4.57 1.335 ;
 RECT 5.86 0.36 6 2.035 ;
 RECT 4.43 0.53 5.315 0.67 ;
 RECT 5.175 0.22 6 0.36 ;
 RECT 5.815 2.17 5.955 2.305 ;
 RECT 5.815 2.035 6 2.17 ;
 RECT 5.175 0.36 5.315 0.53 ;
 RECT 0.835 1.105 0.975 2.045 ;
 RECT 0.835 0.54 0.975 0.965 ;
 RECT 0.835 2.185 0.975 2.66 ;
 RECT 0.835 2.045 1.175 2.185 ;
 RECT 0.835 0.965 1.185 1.105 ;
 RECT 2.86 1.33 3.28 1.47 ;
 RECT 3.14 0.54 3.28 1.33 ;
 RECT 0.835 0.4 3.28 0.54 ;
 RECT 12.835 2.4 13.065 2.54 ;
 RECT 21.72 2.4 21.86 2.52 ;
 RECT 12.835 2.26 21.86 2.4 ;
 RECT 26.06 2.48 26.2 2.52 ;
 RECT 21.72 2.52 26.2 2.66 ;
 RECT 26.06 2.27 26.29 2.48 ;
 RECT 14.36 1.51 14.5 1.695 ;
 RECT 15.335 1.095 15.475 1.37 ;
 RECT 16.26 1.25 16.49 1.37 ;
 RECT 15.3 1.51 15.44 1.7 ;
 RECT 14.36 1.37 16.49 1.51 ;
 RECT 14.29 1.695 14.57 1.835 ;
 RECT 15.265 0.955 15.545 1.095 ;
 RECT 15.235 1.7 15.51 1.84 ;
 RECT 12.97 2.05 13.11 2.055 ;
 RECT 16.01 1.87 16.195 1.98 ;
 RECT 12.97 1.915 14.145 1.98 ;
 RECT 12.97 1.91 14.14 1.915 ;
 RECT 12.97 1.615 13.11 1.91 ;
 RECT 12.97 1.98 16.195 2.05 ;
 RECT 14 2.05 16.195 2.12 ;
 RECT 16.01 1.66 16.24 1.87 ;
 RECT 12.955 1.405 13.185 1.615 ;
 RECT 6.715 2.12 7.815 2.26 ;
 RECT 9.48 1.62 9.62 1.735 ;
 RECT 9.48 1.875 9.62 2.18 ;
 RECT 9.48 0.81 9.62 1.41 ;
 RECT 9.32 1.41 9.62 1.62 ;
 RECT 10.54 1.415 10.68 1.735 ;
 RECT 9.48 1.735 10.68 1.875 ;
 RECT 10.48 1.275 10.75 1.415 ;
 RECT 7.275 1.44 7.415 1.52 ;
 RECT 6.545 1.52 7.415 1.66 ;
 RECT 8.55 0.865 8.69 1.3 ;
 RECT 7.275 1.3 8.69 1.44 ;
 RECT 8.55 1.44 8.69 2.215 ;
 RECT 4.67 1.63 4.81 1.99 ;
 RECT 4.755 0.825 4.895 1.475 ;
 RECT 4.67 1.475 5.015 1.63 ;
 RECT 4.56 1.99 4.81 2.13 ;
 RECT 7.595 1.79 7.735 1.82 ;
 RECT 6.24 1.96 6.52 2.215 ;
 RECT 6.155 1.22 6.47 1.36 ;
 RECT 6.33 0.805 6.47 1.22 ;
 RECT 6.155 1.82 7.735 1.96 ;
 RECT 6.155 1.36 6.295 1.82 ;
 RECT 8.17 1.58 8.41 1.65 ;
 RECT 7.595 1.65 8.41 1.79 ;
 RECT 8.17 1.79 8.41 1.835 ;
 RECT 3.14 2.435 4.01 2.565 ;
 RECT 3.195 2.565 4.01 2.575 ;
 RECT 3.14 1.81 3.28 2.435 ;
 RECT 2.58 1.81 2.72 1.9 ;
 RECT 2.39 2.04 2.53 2.255 ;
 RECT 2.315 0.965 2.72 1.105 ;
 RECT 2.58 1.105 2.72 1.67 ;
 RECT 3.78 2.4 4.01 2.435 ;
 RECT 3.78 2.575 4.01 2.61 ;
 RECT 2.39 1.9 2.72 2.04 ;
 RECT 2.58 1.67 3.285 1.81 ;
 RECT 1.92 2.465 3 2.605 ;
 RECT 2.86 1.98 3 2.465 ;
 RECT 1.92 1.98 2.06 2.465 ;
 RECT 1.92 0.825 2.06 0.965 ;
 RECT 1.92 0.685 3 0.825 ;
 RECT 2.86 0.825 3 1.16 ;
 RECT 1.845 0.965 2.13 1.105 ;
 RECT 24.765 0.73 24.905 1.04 ;
 RECT 24.905 1.18 25.045 1.605 ;
 END
END RDFFSRSSRX1

MACRO RDFFSRSSRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 32 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 32 0.08 ;
 RECT 28.585 0.08 28.825 0.26 ;
 RECT 11.265 0.595 11.54 0.735 ;
 RECT 20.135 0.335 20.4 0.495 ;
 RECT 18.945 0.335 19.21 0.495 ;
 RECT 1.61 0.08 1.91 0.26 ;
 RECT 0.43 0.08 0.57 0.775 ;
 RECT 8.455 0.08 8.69 0.595 ;
 RECT 5.11 0.08 5.25 1.055 ;
 RECT 5.855 0.08 5.995 0.39 ;
 RECT 15.19 0.08 15.33 0.945 ;
 RECT 16.695 0.08 16.835 0.525 ;
 RECT 21.87 0.08 22.01 0.82 ;
 RECT 26.235 0.08 26.375 0.36 ;
 RECT 27.45 0.08 27.59 0.35 ;
 RECT 11.33 0.08 11.47 0.595 ;
 RECT 20.19 0.08 20.33 0.335 ;
 RECT 19 0.08 19.14 0.335 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 32 2.96 ;
 RECT 15.72 2.52 15.995 2.66 ;
 RECT 1.715 1.98 1.855 2.8 ;
 RECT 0.435 1.74 0.575 2.8 ;
 RECT 5.785 2.34 6.035 2.8 ;
 RECT 5.11 1.98 5.25 2.8 ;
 RECT 11.14 2.375 11.28 2.8 ;
 RECT 9.04 2.07 9.18 2.8 ;
 RECT 16.69 2.5 16.83 2.8 ;
 RECT 18.915 2.5 19.055 2.8 ;
 RECT 20.145 2.5 20.285 2.8 ;
 RECT 21.705 2.5 21.845 2.8 ;
 RECT 22.91 2.5 23.05 2.8 ;
 RECT 16.135 2.5 16.365 2.8 ;
 RECT 15.79 2.66 15.93 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.16 1.475 5.49 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.49 1.905 19.63 1.91 ;
 RECT 19.49 0.915 19.63 1.765 ;
 RECT 20.75 1.905 20.89 1.91 ;
 RECT 18.51 1.765 20.89 1.905 ;
 RECT 20.75 0.915 20.89 1.765 ;
 RECT 18.51 0.915 18.65 1.765 ;
 END
 ANTENNADIFFAREA 1.311 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 21.07 1.22 21.37 1.46 ;
 RECT 21.23 1.765 23.845 1.905 ;
 RECT 21.16 0.94 21.44 1.08 ;
 RECT 22.345 1.905 22.485 1.91 ;
 RECT 22.345 0.56 22.485 1.765 ;
 RECT 21.23 1.905 21.37 1.915 ;
 RECT 21.23 1.46 21.37 1.765 ;
 RECT 21.23 1.08 21.37 1.22 ;
 RECT 21.23 0.915 21.37 0.94 ;
 END
 ANTENNADIFFAREA 1.473 ;
 END QN

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.72 1.16 11.015 1.505 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 30.145 1.435 30.485 1.8 ;
 RECT 28.465 1.99 30.33 2.13 ;
 RECT 26.235 2.22 28.605 2.36 ;
 RECT 30.19 1.8 30.33 1.99 ;
 RECT 28.465 1.435 28.605 1.99 ;
 RECT 26.235 1.39 26.375 2.22 ;
 RECT 27.62 1.37 27.76 2.22 ;
 RECT 28.465 2.13 28.605 2.22 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 24.835 0.745 25.16 1.09 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.07 1.455 2.625 1.735 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.43 1.48 1.745 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SETB

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.685 0.465 3.99 0.675 ;
 RECT 3.69 0.675 3.99 0.76 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END RSTB

 OBS
 LAYER PO ;
 RECT 13.315 0.885 13.545 0.925 ;
 RECT 13.315 1.025 13.545 1.095 ;
 RECT 13.315 0.925 14.16 1.025 ;
 RECT 13.995 0.585 14.225 0.795 ;
 RECT 16.945 1.635 17.045 1.66 ;
 RECT 16.945 1.66 17.2 1.87 ;
 RECT 16.945 1.87 17.045 2.565 ;
 RECT 18.775 0.39 18.875 1.31 ;
 RECT 18.775 1.41 18.875 2.27 ;
 RECT 20.48 0.395 20.58 1.31 ;
 RECT 19.93 0.395 20.03 1.31 ;
 RECT 19.255 0.395 19.355 1.31 ;
 RECT 18.775 1.31 20.58 1.41 ;
 RECT 20.48 1.41 20.58 2.27 ;
 RECT 19.93 1.41 20.03 2.27 ;
 RECT 19.255 1.41 19.355 2.27 ;
 RECT 17.525 0.225 17.755 0.29 ;
 RECT 17.525 0.39 17.755 0.435 ;
 RECT 17.525 0.29 18.875 0.39 ;
 RECT 17.22 1.25 17.48 1.3 ;
 RECT 17.38 0.61 17.48 1.25 ;
 RECT 17.22 1.4 17.48 1.46 ;
 RECT 17.38 1.46 17.48 2.56 ;
 RECT 17.91 0.84 18.01 1.3 ;
 RECT 17.22 1.3 18.01 1.4 ;
 RECT 17.895 0.63 18.125 0.84 ;
 RECT 16.045 0.81 16.145 2.5 ;
 RECT 16.045 2.5 16.365 2.71 ;
 RECT 16.005 0.6 16.235 0.81 ;
 RECT 14.72 0.455 15.74 0.47 ;
 RECT 14.8 0.37 15.74 0.455 ;
 RECT 14.72 0.47 14.95 0.665 ;
 RECT 15.575 0.47 15.74 0.625 ;
 RECT 15.575 0.835 15.675 2.21 ;
 RECT 15.575 0.625 15.805 0.835 ;
 RECT 11.985 2.69 13.895 2.695 ;
 RECT 13.795 2.54 13.895 2.69 ;
 RECT 12.775 2.695 13.895 2.79 ;
 RECT 11.985 0.655 12.085 2.595 ;
 RECT 11.985 2.595 12.875 2.69 ;
 RECT 13.795 2.33 14.025 2.54 ;
 RECT 13.02 0.19 13.12 1.29 ;
 RECT 6.53 0.185 13.12 0.19 ;
 RECT 13.915 1.39 14.11 1.405 ;
 RECT 6.53 0.285 6.63 0.51 ;
 RECT 6.53 0.19 8.365 0.285 ;
 RECT 8.265 0.285 8.365 1.24 ;
 RECT 8.265 0.09 13.12 0.185 ;
 RECT 13.02 1.29 14.11 1.39 ;
 RECT 6.49 0.51 6.735 0.755 ;
 RECT 13.915 1.405 14.145 1.615 ;
 RECT 9.315 0.475 9.5 0.5 ;
 RECT 16.95 0.19 17.05 1.18 ;
 RECT 14.41 0.09 17.05 0.19 ;
 RECT 14.41 0.19 14.51 1.91 ;
 RECT 13.59 1.71 13.69 1.91 ;
 RECT 12.505 0.475 12.605 1.61 ;
 RECT 12.505 1.61 13.69 1.71 ;
 RECT 12.505 1.71 12.605 1.725 ;
 RECT 13.055 1.71 13.155 2.445 ;
 RECT 13.59 1.91 14.51 2.01 ;
 RECT 9.315 0.375 12.605 0.475 ;
 RECT 9.27 0.5 9.5 0.71 ;
 RECT 9.77 1.575 9.87 2.485 ;
 RECT 10.28 1.41 10.51 1.475 ;
 RECT 10.28 1.575 10.51 1.62 ;
 RECT 9.77 1.475 10.51 1.575 ;
 RECT 1.5 0.74 1.6 1.485 ;
 RECT 1.5 1.72 1.6 2.465 ;
 RECT 1.465 1.485 1.695 1.72 ;
 RECT 2.91 0.745 3.01 1.28 ;
 RECT 2.91 1.28 3.42 1.515 ;
 RECT 1.97 1.775 2.07 2.675 ;
 RECT 1.055 2.375 1.285 2.675 ;
 RECT 1.055 2.675 2.07 2.775 ;
 RECT 2.44 0.745 2.54 1.475 ;
 RECT 2.44 1.71 2.54 2.465 ;
 RECT 2.395 1.475 2.625 1.71 ;
 RECT 7.965 0.695 8.065 1.61 ;
 RECT 8 1.71 8.1 2.48 ;
 RECT 7.965 1.61 8.1 1.71 ;
 RECT 7.845 0.465 8.085 0.695 ;
 RECT 9.13 1.61 9.395 1.82 ;
 RECT 9.295 1.82 9.395 2.49 ;
 RECT 8.925 0.66 9.025 1.51 ;
 RECT 8.925 1.51 9.395 1.61 ;
 RECT 7.03 1.595 7.13 2.48 ;
 RECT 6.49 1.445 6.735 1.495 ;
 RECT 6.49 1.595 6.735 1.69 ;
 RECT 6.49 1.495 7.13 1.595 ;
 RECT 11.59 0.655 11.69 1.24 ;
 RECT 11.46 1.24 11.69 1.475 ;
 RECT 5.37 0.655 5.47 1.495 ;
 RECT 5.175 1.495 5.47 1.745 ;
 RECT 5.37 1.745 5.47 2.37 ;
 RECT 4.895 0.52 4.995 2.465 ;
 RECT 4.655 0.27 4.995 0.52 ;
 RECT 7.525 1.33 7.665 1.475 ;
 RECT 7.525 1.71 7.625 2.475 ;
 RECT 7.565 0.65 7.665 1.33 ;
 RECT 7.525 1.475 7.755 1.71 ;
 RECT 6.145 1.62 6.245 2.69 ;
 RECT 7.075 0.47 7.36 0.705 ;
 RECT 7.075 0.705 7.175 1.165 ;
 RECT 6.21 0.585 6.31 1.165 ;
 RECT 6.21 1.265 6.31 1.52 ;
 RECT 5.71 1.44 5.955 1.52 ;
 RECT 5.71 1.62 5.955 1.69 ;
 RECT 5.71 1.52 6.31 1.62 ;
 RECT 8.825 1.79 8.925 2.69 ;
 RECT 6.21 1.165 7.175 1.265 ;
 RECT 6.145 2.69 8.925 2.79 ;
 RECT 3.605 0.685 3.705 1.71 ;
 RECT 2.91 1.81 3.01 2.465 ;
 RECT 1.97 0.465 3.915 0.565 ;
 RECT 3.605 0.565 3.915 0.685 ;
 RECT 1.97 0.565 2.07 1.325 ;
 RECT 2.91 1.71 3.705 1.81 ;
 RECT 21.49 0.4 21.59 1.2 ;
 RECT 21.49 1.2 21.76 1.33 ;
 RECT 22.13 0.26 22.23 1.33 ;
 RECT 22.13 1.43 22.23 2.565 ;
 RECT 23.315 0.39 23.415 1.33 ;
 RECT 22.625 1.43 22.725 2.565 ;
 RECT 21.49 1.43 21.76 1.435 ;
 RECT 21.49 1.435 21.59 2.57 ;
 RECT 21.49 1.33 23.415 1.43 ;
 RECT 23.315 1.43 23.415 2.565 ;
 RECT 24.35 0.235 24.58 0.29 ;
 RECT 24.35 0.39 24.58 0.445 ;
 RECT 23.315 0.29 24.58 0.39 ;
 RECT 29.195 2.27 29.48 2.48 ;
 RECT 29.195 1.2 29.295 2.27 ;
 RECT 29.195 0.375 29.295 0.99 ;
 RECT 29.195 0.99 29.445 1.2 ;
 RECT 27.71 1.06 27.81 1.14 ;
 RECT 27.71 0.38 27.81 0.96 ;
 RECT 27.71 1.14 27.98 1.24 ;
 RECT 27.88 1.24 27.98 1.84 ;
 RECT 27.29 0.935 27.52 0.96 ;
 RECT 27.29 0.96 27.81 1.06 ;
 RECT 27.29 1.06 27.52 1.145 ;
 RECT 28.075 0.22 28.305 0.28 ;
 RECT 28.075 0.38 28.305 0.43 ;
 RECT 27.71 0.28 28.305 0.38 ;
 RECT 26.8 0.215 26.9 0.995 ;
 RECT 26.8 0.995 27.04 1.205 ;
 RECT 26.8 1.205 26.9 2 ;
 RECT 25.26 1.1 25.545 1.245 ;
 RECT 29.895 0.195 29.995 2.665 ;
 RECT 28.885 0.095 29.995 0.195 ;
 RECT 25.26 1.245 25.36 2.665 ;
 RECT 28.885 0.195 28.985 0.945 ;
 RECT 25.315 1.035 25.545 1.1 ;
 RECT 25.26 2.665 29.995 2.765 ;
 RECT 26.02 0.21 26.12 0.755 ;
 RECT 26.02 0.855 26.12 2.2 ;
 RECT 28.885 1.125 28.985 2.2 ;
 RECT 24.835 0.755 26.59 0.84 ;
 RECT 24.835 0.84 26.585 0.855 ;
 RECT 26.49 0.215 26.59 0.755 ;
 RECT 24.835 0.855 25.065 0.965 ;
 RECT 26.02 2.2 28.985 2.3 ;
 RECT 26.495 1.245 26.595 2.02 ;
 RECT 26.365 1.035 26.595 1.245 ;
 RECT 10.695 1.45 10.795 1.655 ;
 RECT 10.695 1.755 10.795 2.57 ;
 RECT 10.695 1.655 11.655 1.755 ;
 RECT 11.555 1.755 11.655 2.355 ;
 RECT 10.695 0.655 10.795 1.13 ;
 RECT 10.695 1.23 10.795 1.24 ;
 RECT 9.78 0.66 9.88 1.13 ;
 RECT 10.695 1.24 10.95 1.45 ;
 RECT 9.78 1.13 10.795 1.23 ;
 RECT 13.995 0.795 14.16 0.925 ;
 LAYER CO ;
 RECT 28.125 0.26 28.255 0.39 ;
 RECT 26.86 1.035 26.99 1.165 ;
 RECT 25.365 1.075 25.495 1.205 ;
 RECT 24.885 0.795 25.015 0.925 ;
 RECT 26.415 1.075 26.545 1.205 ;
 RECT 10.77 1.28 10.9 1.41 ;
 RECT 14.77 0.495 14.9 0.625 ;
 RECT 14.045 0.625 14.175 0.755 ;
 RECT 13.365 0.925 13.495 1.055 ;
 RECT 17.945 0.67 18.075 0.8 ;
 RECT 17.02 1.7 17.15 1.83 ;
 RECT 17.575 0.265 17.705 0.395 ;
 RECT 17.27 1.29 17.4 1.42 ;
 RECT 16.055 0.64 16.185 0.77 ;
 RECT 15.625 0.665 15.755 0.795 ;
 RECT 13.845 2.37 13.975 2.5 ;
 RECT 13.965 1.445 14.095 1.575 ;
 RECT 9.32 0.54 9.45 0.67 ;
 RECT 10.33 1.45 10.46 1.58 ;
 RECT 21.59 1.25 21.72 1.38 ;
 RECT 21.875 0.62 22.005 0.75 ;
 RECT 3.13 2.05 3.26 2.18 ;
 RECT 3.24 1.335 3.37 1.465 ;
 RECT 2.445 1.53 2.575 1.66 ;
 RECT 1.25 0.97 1.38 1.1 ;
 RECT 1.73 0.125 1.86 0.255 ;
 RECT 3.13 0.97 3.26 1.1 ;
 RECT 1.105 2.43 1.235 2.56 ;
 RECT 2.66 2.05 2.79 2.18 ;
 RECT 2.66 0.97 2.79 1.1 ;
 RECT 2.19 0.97 2.32 1.1 ;
 RECT 1.72 2.05 1.85 2.18 ;
 RECT 1.25 2.05 1.38 2.18 ;
 RECT 1.515 1.54 1.645 1.67 ;
 RECT 2.19 2.05 2.32 2.18 ;
 RECT 23.63 1.77 23.76 1.9 ;
 RECT 20.755 0.97 20.885 1.1 ;
 RECT 20.755 1.705 20.885 1.835 ;
 RECT 22.915 2.57 23.045 2.7 ;
 RECT 20.195 0.36 20.325 0.49 ;
 RECT 20.15 2.57 20.28 2.7 ;
 RECT 18.92 2.57 19.05 2.7 ;
 RECT 21.235 0.95 21.365 1.08 ;
 RECT 15.195 0.745 15.325 0.875 ;
 RECT 17.6 0.83 17.73 0.96 ;
 RECT 16.7 0.33 16.83 0.46 ;
 RECT 17.6 1.78 17.73 1.91 ;
 RECT 16.695 2.57 16.825 2.7 ;
 RECT 16.3 0.96 16.43 1.09 ;
 RECT 16.265 1.665 16.395 1.795 ;
 RECT 15.795 2.525 15.925 2.655 ;
 RECT 15.325 1.665 15.455 1.795 ;
 RECT 11.145 2.445 11.275 2.575 ;
 RECT 5.59 1.995 5.72 2.125 ;
 RECT 7.575 1.525 7.705 1.655 ;
 RECT 6.825 0.88 6.955 1.01 ;
 RECT 9.515 0.93 9.645 1.06 ;
 RECT 7.18 0.525 7.31 0.655 ;
 RECT 10.445 1.995 10.575 2.125 ;
 RECT 10 0.88 10.13 1.01 ;
 RECT 5.77 1.495 5.9 1.625 ;
 RECT 12.245 0.875 12.375 1.005 ;
 RECT 9.185 1.63 9.315 1.76 ;
 RECT 18.515 0.975 18.645 1.105 ;
 RECT 13.275 0.595 13.405 0.725 ;
 RECT 13.275 1.87 13.405 2 ;
 RECT 12.77 0.595 12.9 0.725 ;
 RECT 12.77 1.9 12.9 2.03 ;
 RECT 25.77 1.425 25.9 1.555 ;
 RECT 28.1 1.405 28.23 1.535 ;
 RECT 30.195 1.475 30.325 1.605 ;
 RECT 29.415 0.595 29.545 0.725 ;
 RECT 26.24 1.475 26.37 1.605 ;
 RECT 28.635 0.12 28.765 0.25 ;
 RECT 29.415 1.465 29.545 1.595 ;
 RECT 28.47 1.49 28.6 1.62 ;
 RECT 27.96 0.595 28.09 0.725 ;
 RECT 26.24 0.135 26.37 0.265 ;
 RECT 27.625 1.445 27.755 1.575 ;
 RECT 27.02 1.485 27.15 1.615 ;
 RECT 27.02 0.435 27.15 0.565 ;
 RECT 25.52 0.505 25.65 0.635 ;
 RECT 27.455 0.12 27.585 0.25 ;
 RECT 22.35 0.63 22.48 0.76 ;
 RECT 22.35 1.71 22.48 1.84 ;
 RECT 21.71 2.57 21.84 2.7 ;
 RECT 19.005 0.36 19.135 0.49 ;
 RECT 19.495 0.97 19.625 1.1 ;
 RECT 19.495 1.705 19.625 1.835 ;
 RECT 18.515 1.705 18.645 1.835 ;
 RECT 21.235 1.725 21.365 1.855 ;
 RECT 6.365 1.825 6.495 1.955 ;
 RECT 11.51 1.28 11.64 1.41 ;
 RECT 9.515 2.015 9.645 2.145 ;
 RECT 0.44 2.085 0.57 2.215 ;
 RECT 10.445 0.88 10.575 1.01 ;
 RECT 12.245 1.945 12.375 2.075 ;
 RECT 0.435 0.33 0.565 0.46 ;
 RECT 11.335 0.595 11.465 0.725 ;
 RECT 0.44 2.345 0.57 2.475 ;
 RECT 7.9 0.515 8.03 0.645 ;
 RECT 7.275 2.07 7.405 2.2 ;
 RECT 5.115 0.875 5.245 1.005 ;
 RECT 8.505 0.455 8.635 0.585 ;
 RECT 6.545 1.49 6.675 1.62 ;
 RECT 6.545 0.555 6.675 0.685 ;
 RECT 7.295 0.88 7.425 1.01 ;
 RECT 4.715 0.325 4.845 0.455 ;
 RECT 4.645 0.875 4.775 1.005 ;
 RECT 9.045 2.135 9.175 2.265 ;
 RECT 5.855 2.345 5.985 2.475 ;
 RECT 10 2.07 10.13 2.2 ;
 RECT 0.435 0.59 0.565 0.72 ;
 RECT 4.645 2.115 4.775 2.245 ;
 RECT 7.745 2.125 7.875 2.255 ;
 RECT 6.43 0.905 6.56 1.035 ;
 RECT 6.78 2.105 6.91 2.235 ;
 RECT 5.72 0.875 5.85 1.005 ;
 RECT 5.115 2.05 5.245 2.18 ;
 RECT 8.225 1.825 8.355 1.955 ;
 RECT 5.235 1.55 5.365 1.68 ;
 RECT 5.86 0.21 5.99 0.34 ;
 RECT 0.44 1.825 0.57 1.955 ;
 RECT 8.575 2.125 8.705 2.255 ;
 RECT 3.735 0.505 3.865 0.635 ;
 RECT 16.185 2.54 16.315 2.67 ;
 RECT 24.4 0.275 24.53 0.405 ;
 RECT 29.3 2.31 29.43 2.44 ;
 RECT 27.34 0.975 27.47 1.105 ;
 RECT 29.265 1.03 29.395 1.16 ;
 LAYER M1 ;
 RECT 28.305 0.71 29.865 0.85 ;
 RECT 29.41 0.51 29.55 0.71 ;
 RECT 29.41 1.385 29.865 1.525 ;
 RECT 25.315 1.225 25.545 1.245 ;
 RECT 25.315 1.195 25.905 1.225 ;
 RECT 25.455 1.015 25.765 1.035 ;
 RECT 25.315 1.035 25.765 1.055 ;
 RECT 25.59 0.64 25.73 1.015 ;
 RECT 25.765 1.225 25.905 1.75 ;
 RECT 25.47 0.5 25.73 0.64 ;
 RECT 26.365 1.035 26.595 1.055 ;
 RECT 26.365 1.195 26.595 1.245 ;
 RECT 25.315 1.055 26.595 1.195 ;
 RECT 27.335 1.145 27.475 1.345 ;
 RECT 27.015 1.485 27.155 1.76 ;
 RECT 27.335 0.73 27.475 0.935 ;
 RECT 27.015 0.355 27.155 0.59 ;
 RECT 27.015 1.345 27.475 1.485 ;
 RECT 27.29 0.935 27.52 1.145 ;
 RECT 27.015 0.59 27.475 0.73 ;
 RECT 24.35 0.36 24.58 0.445 ;
 RECT 25.87 0.36 26.01 0.565 ;
 RECT 24.35 0.235 26.01 0.36 ;
 RECT 24.475 0.22 26.01 0.235 ;
 RECT 26.61 0.705 26.75 0.75 ;
 RECT 26.735 0.995 27.04 1.205 ;
 RECT 26.735 0.89 26.875 0.995 ;
 RECT 26.61 0.75 26.875 0.89 ;
 RECT 25.87 0.565 26.75 0.705 ;
 RECT 13.995 0.585 14.95 0.63 ;
 RECT 14.72 0.63 14.95 0.665 ;
 RECT 14.72 0.455 14.95 0.49 ;
 RECT 14.02 0.49 14.95 0.585 ;
 RECT 13.995 0.63 14.225 0.795 ;
 RECT 17.895 0.63 18.125 0.635 ;
 RECT 17.895 0.775 18.125 0.84 ;
 RECT 21.585 0.775 21.725 1.46 ;
 RECT 17.89 0.635 21.725 0.775 ;
 RECT 16.375 0.36 16.515 0.665 ;
 RECT 15.575 0.22 16.52 0.36 ;
 RECT 15.575 0.36 15.805 0.835 ;
 RECT 17.595 0.22 17.735 0.225 ;
 RECT 17.595 0.435 17.735 0.665 ;
 RECT 16.375 0.665 17.735 0.805 ;
 RECT 17.595 0.805 17.735 1.98 ;
 RECT 17.525 0.225 17.755 0.435 ;
 RECT 13.27 0.525 13.41 0.885 ;
 RECT 13.27 1.095 13.41 2.065 ;
 RECT 13.27 0.885 13.545 1.095 ;
 RECT 9.995 0.82 10.135 2.33 ;
 RECT 9.995 2.47 10.135 2.475 ;
 RECT 10.845 2.165 10.985 2.33 ;
 RECT 10.845 2.47 10.985 2.475 ;
 RECT 9.995 2.33 10.985 2.47 ;
 RECT 11.925 2.165 12.065 2.295 ;
 RECT 12.24 0.765 12.38 2.295 ;
 RECT 12.24 2.435 12.38 2.44 ;
 RECT 12.765 0.525 12.905 2.295 ;
 RECT 12.765 2.435 12.905 2.44 ;
 RECT 10.845 2.025 12.065 2.165 ;
 RECT 11.925 2.295 12.905 2.435 ;
 RECT 6.425 0.5 6.68 0.965 ;
 RECT 6.425 1.67 6.565 1.82 ;
 RECT 6.425 1.96 6.565 2.65 ;
 RECT 6.425 0.965 6.565 1.44 ;
 RECT 6.425 1.44 6.68 1.67 ;
 RECT 6.295 1.82 6.565 1.96 ;
 RECT 7.11 0.52 7.71 0.66 ;
 RECT 7.57 0.66 7.71 1.015 ;
 RECT 9.115 0.505 9.5 0.71 ;
 RECT 9.27 0.5 9.5 0.505 ;
 RECT 9.115 0.71 9.255 1.015 ;
 RECT 7.57 1.015 9.255 1.155 ;
 RECT 4.42 1.01 4.56 1.195 ;
 RECT 4.42 1.335 4.56 2.11 ;
 RECT 4.42 2.25 4.56 2.255 ;
 RECT 4.42 2.11 4.845 2.25 ;
 RECT 4.42 0.87 4.845 1.01 ;
 RECT 5.39 0.67 5.53 1.195 ;
 RECT 4.42 1.195 5.53 1.335 ;
 RECT 6.82 0.36 6.96 2.035 ;
 RECT 6.135 0.22 6.96 0.36 ;
 RECT 5.39 0.53 6.275 0.67 ;
 RECT 6.775 2.17 6.915 2.305 ;
 RECT 6.775 2.035 6.96 2.17 ;
 RECT 6.135 0.36 6.275 0.53 ;
 RECT 10.325 0.36 10.465 0.525 ;
 RECT 8.83 0.36 8.97 0.735 ;
 RECT 8.83 0.22 10.465 0.36 ;
 RECT 7.895 0.735 8.97 0.875 ;
 RECT 7.895 0.695 8.085 0.735 ;
 RECT 7.895 0.445 8.035 0.465 ;
 RECT 7.86 0.465 8.085 0.695 ;
 RECT 11.705 0.385 11.845 0.875 ;
 RECT 13.715 0.385 13.855 1.09 ;
 RECT 11.705 0.255 13.855 0.385 ;
 RECT 11.705 0.245 13.85 0.255 ;
 RECT 10.73 0.875 11.845 1.015 ;
 RECT 10.73 0.665 10.87 0.875 ;
 RECT 10.325 0.525 10.87 0.665 ;
 RECT 15.945 0.6 16.235 0.81 ;
 RECT 15.945 0.81 16.085 1.09 ;
 RECT 13.715 1.09 16.085 1.23 ;
 RECT 1.1 1.105 1.24 2.045 ;
 RECT 1.1 0.54 1.24 0.965 ;
 RECT 1.1 2.185 1.24 2.63 ;
 RECT 1.1 2.045 1.44 2.185 ;
 RECT 1.1 0.965 1.45 1.105 ;
 RECT 3.125 1.33 3.545 1.47 ;
 RECT 3.405 0.54 3.545 1.33 ;
 RECT 1.1 0.4 3.545 0.54 ;
 RECT 2.845 1.82 2.985 1.9 ;
 RECT 2.655 2.04 2.795 2.255 ;
 RECT 2.58 0.965 2.985 1.105 ;
 RECT 2.845 1.105 2.985 1.68 ;
 RECT 2.655 1.9 2.985 2.04 ;
 RECT 4.135 0.455 4.275 1.68 ;
 RECT 4.605 0.22 4.97 0.315 ;
 RECT 4.605 0.455 4.97 0.615 ;
 RECT 2.845 1.68 4.28 1.82 ;
 RECT 4.135 0.315 4.97 0.455 ;
 RECT 13.795 2.36 14.025 2.54 ;
 RECT 24.91 2.36 25.05 2.52 ;
 RECT 13.795 2.22 25.05 2.36 ;
 RECT 29.25 2.48 29.39 2.52 ;
 RECT 24.91 2.52 29.39 2.66 ;
 RECT 29.25 2.27 29.48 2.48 ;
 RECT 16.295 1.095 16.435 1.37 ;
 RECT 16.26 1.51 16.4 1.66 ;
 RECT 15.32 1.51 15.46 1.66 ;
 RECT 15.32 1.37 17.45 1.51 ;
 RECT 17.22 1.25 17.45 1.37 ;
 RECT 16.225 0.955 16.505 1.095 ;
 RECT 16.195 1.66 16.47 1.8 ;
 RECT 15.25 1.66 15.53 1.8 ;
 RECT 13.93 2.05 14.07 2.055 ;
 RECT 16.97 1.87 17.155 1.94 ;
 RECT 13.93 1.615 14.07 1.91 ;
 RECT 13.93 1.94 17.155 2.05 ;
 RECT 13.93 1.91 15.1 1.94 ;
 RECT 14.965 2.05 17.155 2.08 ;
 RECT 16.97 1.66 17.2 1.87 ;
 RECT 13.915 1.405 14.145 1.615 ;
 RECT 10.44 1.62 10.58 1.735 ;
 RECT 10.44 1.875 10.58 2.18 ;
 RECT 10.44 0.81 10.58 1.41 ;
 RECT 10.28 1.41 10.58 1.62 ;
 RECT 11.49 1.415 11.63 1.735 ;
 RECT 10.44 1.735 11.63 1.875 ;
 RECT 11.46 1.275 11.71 1.415 ;
 RECT 8.235 1.44 8.375 1.52 ;
 RECT 7.505 1.52 8.375 1.66 ;
 RECT 9.51 0.865 9.65 1.3 ;
 RECT 8.235 1.3 9.65 1.44 ;
 RECT 9.51 1.44 9.65 2.215 ;
 RECT 7.675 2.12 8.775 2.26 ;
 RECT 5.63 1.63 5.77 1.99 ;
 RECT 5.63 1.475 5.975 1.63 ;
 RECT 5.715 0.825 5.855 1.475 ;
 RECT 5.52 1.99 5.77 2.13 ;
 RECT 7.115 1.82 8.695 1.96 ;
 RECT 8.555 1.79 8.695 1.82 ;
 RECT 7.115 1.22 7.43 1.36 ;
 RECT 7.29 0.805 7.43 1.22 ;
 RECT 7.2 1.96 7.48 2.215 ;
 RECT 7.115 1.36 7.255 1.82 ;
 RECT 9.13 1.58 9.37 1.65 ;
 RECT 8.555 1.65 9.37 1.79 ;
 RECT 9.13 1.79 9.37 1.835 ;
 RECT 2.185 2.465 3.265 2.605 ;
 RECT 3.125 1.98 3.265 2.465 ;
 RECT 2.185 1.98 2.325 2.465 ;
 RECT 2.185 0.825 2.325 0.965 ;
 RECT 2.185 0.685 3.265 0.825 ;
 RECT 3.125 0.825 3.265 1.16 ;
 RECT 2.11 0.965 2.395 1.105 ;
 RECT 27.955 0.73 28.095 1.04 ;
 RECT 28.095 1.18 28.235 1.605 ;
 RECT 27.89 0.59 28.165 0.73 ;
 RECT 29.215 0.99 29.445 1.04 ;
 RECT 27.955 1.04 29.445 1.18 ;
 RECT 29.215 1.18 29.445 1.2 ;
 RECT 28.075 0.29 28.445 0.43 ;
 RECT 28.305 0.43 28.445 0.71 ;
 RECT 28.075 0.22 28.305 0.29 ;
 RECT 29.725 0.85 29.865 1.385 ;
 RECT 29.41 1.525 29.55 1.73 ;
 END
END RDFFSRSSRX2

MACRO RDFFSRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 24.96 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 15.52 1.16 15.885 1.4 ;
 RECT 15.745 0.695 15.885 1.16 ;
 RECT 16.805 1.905 16.945 1.91 ;
 RECT 15.745 1.765 16.945 1.905 ;
 RECT 16.805 0.71 16.945 1.765 ;
 RECT 15.745 1.4 15.885 1.765 ;
 END
 ANTENNADIFFAREA 0.717 ;
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 24.96 0.08 ;
 RECT 14.655 0.28 14.92 0.44 ;
 RECT 2.18 0.08 2.32 1.055 ;
 RECT 21.785 0.08 22.025 0.31 ;
 RECT 5.525 0.08 5.76 0.595 ;
 RECT 0.68 0.08 0.82 0.775 ;
 RECT 11.575 0.08 11.715 1.155 ;
 RECT 2.925 0.08 3.065 0.39 ;
 RECT 16.305 0.08 16.445 0.965 ;
 RECT 8.4 0.08 8.54 0.815 ;
 RECT 20.65 0.08 20.79 0.325 ;
 RECT 12.65 0.08 12.79 0.525 ;
 RECT 19.435 0.08 19.575 0.31 ;
 RECT 14.71 0.08 14.85 0.28 ;
 END
 END VSS

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.005 0.57 18.485 0.78 ;
 RECT 18.005 0.78 18.375 0.865 ;
 RECT 18.005 0.565 18.375 0.57 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.79 1.16 8.12 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 23.345 1.41 23.685 1.775 ;
 RECT 21.665 1.965 23.53 2.105 ;
 RECT 19.435 2.195 21.805 2.335 ;
 RECT 21.665 1.41 21.805 1.965 ;
 RECT 23.39 1.775 23.53 1.965 ;
 RECT 19.435 1.365 19.575 2.195 ;
 RECT 20.82 1.345 20.96 2.195 ;
 RECT 21.665 2.105 21.805 2.195 ;
 END
 END VDDG

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.23 1.475 2.56 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 24.96 2.96 ;
 RECT 2.855 2.34 3.105 2.8 ;
 RECT 6.11 2.07 6.25 2.8 ;
 RECT 8.21 2.375 8.35 2.8 ;
 RECT 14.705 2.57 14.845 2.8 ;
 RECT 11.8 2.57 11.94 2.8 ;
 RECT 2.18 1.98 2.32 2.8 ;
 RECT 16.22 2.57 16.36 2.8 ;
 RECT 0.725 1.74 0.865 2.8 ;
 RECT 12.645 2.57 12.785 2.8 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.22 1.7 15.365 1.75 ;
 RECT 14.005 1.84 14.36 1.99 ;
 RECT 14.005 1.75 15.365 1.84 ;
 RECT 14.22 0.905 14.36 1.7 ;
 RECT 15.225 0.915 15.365 1.7 ;
 RECT 15.225 1.84 15.365 1.92 ;
 END
 ANTENNADIFFAREA 0.531 ;
 END QN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.675 0.22 2.04 0.615 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 20 0.97 20.24 1.18 ;
 RECT 20 1.18 20.1 1.975 ;
 RECT 12.9 1.635 13 1.66 ;
 RECT 12.9 1.66 13.155 1.87 ;
 RECT 12.9 1.87 13 2.565 ;
 RECT 7.765 1.45 7.865 1.655 ;
 RECT 7.765 1.755 7.865 2.57 ;
 RECT 7.765 0.655 7.865 1.13 ;
 RECT 7.765 1.23 7.865 1.24 ;
 RECT 6.85 0.66 6.95 1.13 ;
 RECT 7.765 1.655 8.725 1.755 ;
 RECT 8.625 1.755 8.725 2.355 ;
 RECT 7.765 1.24 8.02 1.45 ;
 RECT 6.85 1.13 7.865 1.23 ;
 RECT 13.175 1.25 13.435 1.3 ;
 RECT 13.335 0.61 13.435 1.25 ;
 RECT 13.865 0.84 13.965 1.3 ;
 RECT 13.335 1.46 13.435 2.56 ;
 RECT 13.175 1.4 13.435 1.46 ;
 RECT 13.175 1.3 13.965 1.4 ;
 RECT 13.85 0.63 14.08 0.84 ;
 RECT 6.84 1.575 6.94 2.485 ;
 RECT 7.35 1.41 7.58 1.475 ;
 RECT 7.35 1.575 7.58 1.62 ;
 RECT 6.84 1.475 7.58 1.575 ;
 RECT 19.22 0.87 19.32 2.175 ;
 RECT 18.255 0.77 19.79 0.78 ;
 RECT 19.22 0.73 19.79 0.77 ;
 RECT 21.92 1.125 22.02 2.175 ;
 RECT 18.26 0.78 19.79 0.83 ;
 RECT 18.26 0.83 19.32 0.87 ;
 RECT 19.69 0.19 19.79 0.73 ;
 RECT 19.22 0.185 19.32 0.73 ;
 RECT 18.255 0.57 18.485 0.77 ;
 RECT 19.22 2.175 22.02 2.275 ;
 RECT 22.395 0.37 22.495 1.01 ;
 RECT 22.395 1.01 22.645 1.22 ;
 RECT 22.395 1.22 22.495 2.245 ;
 RECT 22.395 2.245 22.68 2.455 ;
 RECT 1.965 0.52 2.065 2.465 ;
 RECT 1.725 0.27 2.065 0.52 ;
 RECT 8.66 0.655 8.76 1.24 ;
 RECT 8.53 1.24 8.76 1.475 ;
 RECT 4.635 1.475 4.945 1.71 ;
 RECT 4.635 0.65 4.735 1.475 ;
 RECT 4.635 1.71 4.735 2.475 ;
 RECT 18.46 1.175 18.745 1.305 ;
 RECT 18.46 1.305 18.56 2.64 ;
 RECT 23.095 0.19 23.195 2.64 ;
 RECT 22.085 0.09 23.195 0.19 ;
 RECT 22.085 0.19 22.185 0.94 ;
 RECT 18.46 1.075 18.79 1.175 ;
 RECT 18.46 2.64 23.195 2.74 ;
 RECT 9.055 2.69 10.705 2.695 ;
 RECT 10.53 2.54 10.705 2.69 ;
 RECT 9.845 2.695 10.705 2.79 ;
 RECT 9.055 0.655 9.155 2.595 ;
 RECT 9.055 2.595 9.945 2.69 ;
 RECT 10.53 2.33 10.76 2.54 ;
 RECT 20.91 0.355 21.01 0.985 ;
 RECT 20.91 0.255 21.645 0.355 ;
 RECT 21.415 0.355 21.645 0.465 ;
 RECT 21.08 1.215 21.18 1.815 ;
 RECT 20.52 1.115 21.18 1.215 ;
 RECT 20.52 0.985 21.01 1.115 ;
 RECT 14.485 0.39 14.585 1.4 ;
 RECT 13.48 0.225 13.71 0.29 ;
 RECT 13.48 0.39 13.71 0.435 ;
 RECT 13.48 0.29 14.585 0.39 ;
 RECT 14.485 1.5 14.585 2.35 ;
 RECT 14.975 0.505 15.075 1.4 ;
 RECT 14.975 1.5 15.075 2.35 ;
 RECT 14.485 1.4 15.075 1.5 ;
 RECT 5.895 1.79 5.995 2.465 ;
 RECT 5.68 2.465 5.995 2.71 ;
 RECT 6.2 1.61 6.465 1.82 ;
 RECT 6.365 1.82 6.465 2.49 ;
 RECT 5.995 0.66 6.095 1.51 ;
 RECT 5.995 1.51 6.465 1.61 ;
 RECT 2.44 0.57 2.54 1.495 ;
 RECT 2.245 1.495 2.54 1.745 ;
 RECT 2.44 1.745 2.54 2.37 ;
 RECT 11.29 0.19 11.39 1.795 ;
 RECT 11.29 0.09 13.005 0.19 ;
 RECT 6.385 0.47 6.57 0.5 ;
 RECT 10.595 1.71 10.695 1.795 ;
 RECT 12.905 0.19 13.005 1.18 ;
 RECT 10.595 1.795 11.39 1.895 ;
 RECT 9.575 0.47 9.675 1.61 ;
 RECT 10.125 1.71 10.225 2.445 ;
 RECT 6.34 0.5 6.57 0.71 ;
 RECT 6.385 0.37 9.675 0.47 ;
 RECT 9.575 1.61 10.695 1.71 ;
 RECT 15.99 1.285 16.685 1.385 ;
 RECT 15.99 1.385 16.2 1.435 ;
 RECT 16.585 0.26 17.485 0.36 ;
 RECT 16.585 0.36 16.685 1.285 ;
 RECT 15.99 1.2 16.2 1.285 ;
 RECT 16.005 0.47 16.105 1.2 ;
 RECT 16.005 1.435 16.105 2.645 ;
 RECT 16.585 1.385 16.685 2.645 ;
 RECT 17.255 0.185 17.485 0.26 ;
 RECT 17.255 0.36 17.485 0.435 ;
 RECT 3.215 2.415 3.64 2.66 ;
 RECT 4.145 0.47 4.43 0.51 ;
 RECT 3.215 1.62 3.315 2.415 ;
 RECT 3.28 0.61 3.38 1.52 ;
 RECT 2.78 1.52 3.38 1.62 ;
 RECT 4.145 0.705 4.245 1.255 ;
 RECT 4.145 0.61 4.43 0.705 ;
 RECT 3.28 0.51 4.43 0.61 ;
 RECT 3.28 0.505 3.38 0.51 ;
 RECT 2.78 1.44 3.025 1.52 ;
 RECT 2.78 1.62 3.025 1.69 ;
 RECT 4.1 1.61 4.2 2.655 ;
 RECT 5.335 0.19 5.435 2.655 ;
 RECT 10.09 1.29 11.11 1.39 ;
 RECT 10.09 0.19 10.19 1.29 ;
 RECT 3.56 1.27 3.805 1.51 ;
 RECT 10.88 1.285 11.11 1.29 ;
 RECT 10.88 1.39 11.11 1.615 ;
 RECT 3.56 1.51 4.2 1.61 ;
 RECT 4.1 2.655 5.435 2.755 ;
 RECT 5.335 0.09 10.19 0.19 ;
 RECT 12.055 0.64 12.155 1.26 ;
 RECT 11.85 1.26 12.155 1.47 ;
 RECT 12.055 1.47 12.155 2.21 ;
 RECT 19.56 1.01 19.795 1.22 ;
 RECT 19.695 1.22 19.795 1.995 ;
 RECT 20 0.19 20.1 0.97 ;
 LAYER CO ;
 RECT 17.305 0.265 17.435 0.395 ;
 RECT 11.9 1.3 12.03 1.43 ;
 RECT 3.615 1.365 3.745 1.495 ;
 RECT 19.61 1.05 19.74 1.18 ;
 RECT 10.93 1.445 11.06 1.575 ;
 RECT 20.57 1.025 20.7 1.155 ;
 RECT 13.225 1.29 13.355 1.42 ;
 RECT 10.58 2.37 10.71 2.5 ;
 RECT 13.53 0.265 13.66 0.395 ;
 RECT 20.06 1.01 20.19 1.14 ;
 RECT 12.975 1.7 13.105 1.83 ;
 RECT 21.465 0.295 21.595 0.425 ;
 RECT 7.84 1.28 7.97 1.41 ;
 RECT 6.39 0.54 6.52 0.67 ;
 RECT 22.465 1.05 22.595 1.18 ;
 RECT 13.9 0.67 14.03 0.8 ;
 RECT 7.4 1.45 7.53 1.58 ;
 RECT 18.305 0.61 18.435 0.74 ;
 RECT 18.565 1.135 18.695 1.265 ;
 RECT 3.44 2.47 3.57 2.6 ;
 RECT 1.715 2.115 1.845 2.245 ;
 RECT 10.345 0.595 10.475 0.725 ;
 RECT 7.515 0.88 7.645 1.01 ;
 RECT 8.58 1.28 8.71 1.41 ;
 RECT 12.655 0.33 12.785 0.46 ;
 RECT 12.275 1.705 12.405 1.835 ;
 RECT 4.25 0.525 4.38 0.655 ;
 RECT 16.225 2.64 16.355 2.77 ;
 RECT 1.715 0.79 1.845 0.92 ;
 RECT 8.405 0.62 8.535 0.75 ;
 RECT 22.5 2.285 22.63 2.415 ;
 RECT 16.31 0.77 16.44 0.9 ;
 RECT 13.555 1.78 13.685 1.91 ;
 RECT 5.575 0.455 5.705 0.585 ;
 RECT 14.225 0.975 14.355 1.105 ;
 RECT 9.315 0.875 9.445 1.005 ;
 RECT 3.85 2.105 3.98 2.235 ;
 RECT 3.435 1.825 3.565 1.955 ;
 RECT 2.185 0.79 2.315 0.92 ;
 RECT 2.925 2.345 3.055 2.475 ;
 RECT 13.555 0.83 13.685 0.96 ;
 RECT 15.75 0.77 15.88 0.9 ;
 RECT 14.225 1.72 14.355 1.85 ;
 RECT 15.75 1.725 15.88 1.855 ;
 RECT 2.84 1.495 2.97 1.625 ;
 RECT 3.895 0.88 4.025 1.01 ;
 RECT 16.03 1.25 16.16 1.38 ;
 RECT 11.805 2.64 11.935 2.77 ;
 RECT 0.685 0.33 0.815 0.46 ;
 RECT 2.93 0.21 3.06 0.34 ;
 RECT 20.655 0.11 20.785 0.24 ;
 RECT 4.365 0.88 4.495 1.01 ;
 RECT 4.345 2.07 4.475 2.2 ;
 RECT 12.65 2.64 12.78 2.77 ;
 RECT 14.71 2.64 14.84 2.77 ;
 RECT 9.315 1.945 9.445 2.075 ;
 RECT 7.515 1.885 7.645 2.015 ;
 RECT 18.72 0.505 18.85 0.635 ;
 RECT 0.73 1.825 0.86 1.955 ;
 RECT 19.44 1.45 19.57 1.58 ;
 RECT 5.645 2.125 5.775 2.255 ;
 RECT 15.23 1.72 15.36 1.85 ;
 RECT 9.84 0.595 9.97 0.725 ;
 RECT 7.07 2.07 7.2 2.2 ;
 RECT 1.785 0.325 1.915 0.455 ;
 RECT 6.255 1.63 6.385 1.76 ;
 RECT 21.135 0.59 21.265 0.72 ;
 RECT 21.67 1.465 21.8 1.595 ;
 RECT 2.305 1.55 2.435 1.68 ;
 RECT 0.73 2.085 0.86 2.215 ;
 RECT 6.115 2.135 6.245 2.265 ;
 RECT 6.585 0.93 6.715 1.06 ;
 RECT 2.185 2.05 2.315 2.18 ;
 RECT 10.345 1.87 10.475 2 ;
 RECT 16.81 0.78 16.94 0.91 ;
 RECT 21.3 1.38 21.43 1.51 ;
 RECT 7.07 0.88 7.2 1.01 ;
 RECT 21.835 0.115 21.965 0.245 ;
 RECT 23.395 1.45 23.525 1.58 ;
 RECT 20.22 0.41 20.35 0.54 ;
 RECT 3.5 0.905 3.63 1.035 ;
 RECT 2.79 0.88 2.92 1.01 ;
 RECT 15.23 0.975 15.36 1.105 ;
 RECT 9.84 1.9 9.97 2.03 ;
 RECT 4.765 1.525 4.895 1.655 ;
 RECT 20.825 1.42 20.955 1.55 ;
 RECT 4.855 2.125 4.985 2.255 ;
 RECT 16.81 1.71 16.94 1.84 ;
 RECT 18.97 1.4 19.1 1.53 ;
 RECT 14.715 0.305 14.845 0.435 ;
 RECT 20.22 1.46 20.35 1.59 ;
 RECT 8.215 2.445 8.345 2.575 ;
 RECT 11.58 0.955 11.71 1.085 ;
 RECT 0.685 0.59 0.815 0.72 ;
 RECT 19.44 0.11 19.57 0.24 ;
 RECT 5.72 2.515 5.85 2.645 ;
 RECT 22.615 1.44 22.745 1.57 ;
 RECT 12.275 0.96 12.405 1.09 ;
 RECT 2.66 1.995 2.79 2.125 ;
 RECT 0.73 2.345 0.86 2.475 ;
 RECT 22.615 0.59 22.745 0.72 ;
 RECT 6.585 2.015 6.715 2.145 ;
 LAYER M1 ;
 RECT 6.58 1.44 6.72 2.215 ;
 RECT 5.305 1.3 6.72 1.44 ;
 RECT 4.745 2.12 5.845 2.26 ;
 RECT 3.495 1.535 3.635 1.82 ;
 RECT 3.495 0.73 3.635 1.325 ;
 RECT 3.495 1.325 3.795 1.535 ;
 RECT 3.365 1.82 3.635 1.96 ;
 RECT 20.52 1.195 20.66 1.32 ;
 RECT 20.215 1.46 20.355 1.735 ;
 RECT 20.535 0.705 20.675 0.985 ;
 RECT 20.215 0.33 20.355 0.565 ;
 RECT 20.215 1.32 20.66 1.46 ;
 RECT 20.215 0.565 20.675 0.705 ;
 RECT 20.52 0.985 20.75 1.195 ;
 RECT 12.27 1.37 13.405 1.46 ;
 RECT 12.27 1.095 12.41 1.37 ;
 RECT 12.27 1.46 13.4 1.51 ;
 RECT 12.27 1.51 12.41 1.7 ;
 RECT 13.175 1.25 13.405 1.37 ;
 RECT 12.205 1.7 12.48 1.84 ;
 RECT 12.2 0.955 12.47 1.095 ;
 RECT 11.855 0.805 11.995 1.26 ;
 RECT 11.85 1.26 12.08 1.295 ;
 RECT 11.85 1.435 12.08 1.47 ;
 RECT 11.26 1.295 12.08 1.435 ;
 RECT 11.26 1.105 11.4 1.295 ;
 RECT 10.34 0.525 10.48 0.965 ;
 RECT 10.34 1.105 10.48 2.065 ;
 RECT 10.34 0.965 11.4 1.105 ;
 RECT 13.55 0.435 13.69 0.665 ;
 RECT 13.55 0.805 13.69 1.98 ;
 RECT 11.855 0.665 13.69 0.805 ;
 RECT 13.55 0.22 13.69 0.225 ;
 RECT 13.48 0.225 13.71 0.435 ;
 RECT 21.505 0.465 21.645 0.685 ;
 RECT 21.415 0.255 21.645 0.465 ;
 RECT 21.505 0.685 23.065 0.825 ;
 RECT 22.925 0.825 23.065 1.36 ;
 RECT 22.61 1.5 22.75 1.705 ;
 RECT 22.61 0.485 22.75 0.685 ;
 RECT 22.61 1.36 23.065 1.5 ;
 RECT 13.85 0.72 14.08 0.84 ;
 RECT 15.12 0.37 15.26 0.58 ;
 RECT 13.85 0.63 15.26 0.72 ;
 RECT 13.86 0.58 15.26 0.63 ;
 RECT 16.025 0.37 16.165 1.46 ;
 RECT 15.12 0.23 16.165 0.37 ;
 RECT 7.51 1.62 7.65 1.735 ;
 RECT 7.51 1.875 7.65 2.085 ;
 RECT 7.51 0.81 7.65 1.41 ;
 RECT 7.35 1.41 7.65 1.62 ;
 RECT 8.57 1.415 8.71 1.735 ;
 RECT 7.51 1.735 8.71 1.875 ;
 RECT 8.515 1.275 8.78 1.415 ;
 RECT 10.53 2.42 10.76 2.54 ;
 RECT 10.53 2.28 18.135 2.42 ;
 RECT 17.995 2.42 18.135 2.505 ;
 RECT 22.45 2.455 22.59 2.505 ;
 RECT 17.995 2.505 22.59 2.645 ;
 RECT 22.45 2.245 22.68 2.455 ;
 RECT 17.255 0.36 17.485 0.435 ;
 RECT 19.07 0.36 19.21 0.54 ;
 RECT 17.255 0.225 19.21 0.36 ;
 RECT 17.29 0.22 19.21 0.225 ;
 RECT 19.935 0.535 20.075 0.54 ;
 RECT 19.935 0.68 20.075 0.97 ;
 RECT 19.935 0.97 20.24 1.18 ;
 RECT 19.07 0.54 20.075 0.68 ;
 RECT 7.065 0.82 7.205 2.225 ;
 RECT 7.915 2.165 8.055 2.225 ;
 RECT 7.065 2.225 8.055 2.365 ;
 RECT 9.835 0.525 9.975 2.025 ;
 RECT 9.31 0.765 9.45 2.025 ;
 RECT 7.915 2.025 9.975 2.165 ;
 RECT 21.13 0.48 21.27 1.08 ;
 RECT 21.295 1.22 21.435 1.58 ;
 RECT 22.415 1.01 22.645 1.08 ;
 RECT 21.13 1.08 22.645 1.22 ;
 RECT 2.7 1.63 2.84 1.99 ;
 RECT 2.7 1.475 3.045 1.63 ;
 RECT 2.785 0.81 2.925 1.475 ;
 RECT 2.59 1.99 2.84 2.13 ;
 RECT 4.18 0.52 4.78 0.66 ;
 RECT 4.64 0.66 4.78 1.015 ;
 RECT 6.185 0.505 6.57 0.71 ;
 RECT 4.64 1.015 6.325 1.155 ;
 RECT 6.34 0.5 6.57 0.505 ;
 RECT 6.185 0.71 6.325 1.015 ;
 RECT 3.38 2.41 3.645 2.51 ;
 RECT 3.38 2.65 3.645 2.655 ;
 RECT 3.38 2.51 5.97 2.65 ;
 RECT 18.79 0.64 18.93 0.99 ;
 RECT 18.515 1.17 19.105 1.2 ;
 RECT 18.965 1.2 19.105 1.725 ;
 RECT 18.655 0.99 18.965 1.03 ;
 RECT 18.515 1.2 18.745 1.305 ;
 RECT 18.67 0.5 18.93 0.64 ;
 RECT 19.56 1.01 19.79 1.03 ;
 RECT 18.51 1.03 19.79 1.17 ;
 RECT 19.56 1.17 19.79 1.22 ;
 RECT 1.49 1.335 1.63 2.11 ;
 RECT 1.49 0.925 1.63 1.195 ;
 RECT 1.49 2.11 1.915 2.25 ;
 RECT 1.49 0.785 1.915 0.925 ;
 RECT 1.49 1.195 2.6 1.335 ;
 RECT 2.46 0.67 2.6 1.195 ;
 RECT 3.205 0.22 4.03 0.36 ;
 RECT 3.89 0.36 4.03 0.9 ;
 RECT 3.965 1.08 4.105 1.945 ;
 RECT 2.46 0.53 3.345 0.67 ;
 RECT 3.205 0.36 3.345 0.53 ;
 RECT 3.89 0.9 4.105 1.08 ;
 RECT 3.845 1.945 4.105 2.17 ;
 RECT 3.845 2.17 3.985 2.305 ;
 RECT 5.625 1.79 5.765 1.82 ;
 RECT 4.27 1.96 4.55 2.215 ;
 RECT 4.27 1.82 5.765 1.96 ;
 RECT 4.36 0.805 4.5 1.82 ;
 RECT 6.2 1.58 6.44 1.65 ;
 RECT 5.625 1.65 6.44 1.79 ;
 RECT 6.2 1.79 6.44 1.835 ;
 RECT 10.875 1.43 11.11 1.615 ;
 RECT 10.875 1.615 11.015 1.985 ;
 RECT 10.88 1.405 11.11 1.43 ;
 RECT 10.875 1.985 13.11 2.125 ;
 RECT 12.925 1.87 13.11 1.985 ;
 RECT 12.925 1.66 13.155 1.87 ;
 RECT 4.695 1.52 5.445 1.66 ;
 RECT 5.305 1.44 5.445 1.52 ;
 RECT 6.58 0.865 6.72 1.3 ;
 END
END RDFFSRX1

MACRO RDFFSRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 24.64 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.585 0.57 18.065 0.78 ;
 RECT 17.585 0.78 17.955 0.865 ;
 RECT 17.585 0.565 17.955 0.57 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 24.64 0.08 ;
 RECT 13.645 0.28 13.91 0.44 ;
 RECT 4.85 0.08 5.085 0.595 ;
 RECT 21.365 0.08 21.605 0.31 ;
 RECT 1.505 0.08 1.645 1.055 ;
 RECT 10.34 0.08 10.48 1.155 ;
 RECT 16.575 0.08 16.715 0.965 ;
 RECT 11.415 0.08 11.555 0.525 ;
 RECT 15.63 0.08 15.77 0.965 ;
 RECT 19.015 0.08 19.155 0.31 ;
 RECT 2.25 0.08 2.39 0.39 ;
 RECT 0.47 0.08 0.61 0.775 ;
 RECT 7.725 0.08 7.865 0.815 ;
 RECT 20.23 0.08 20.37 0.325 ;
 RECT 13.7 0.08 13.84 0.28 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.01 1.205 13.365 1.445 ;
 RECT 12.615 1.705 14.77 1.845 ;
 RECT 13.22 0.88 13.36 1.205 ;
 RECT 14.23 0.89 14.37 1.705 ;
 RECT 13.22 1.445 13.36 1.705 ;
 END
 ANTENNADIFFAREA 0.815 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.845 1.16 15.2 1.4 ;
 RECT 14.97 0.695 15.11 1.16 ;
 RECT 14.97 1.765 17.185 1.905 ;
 RECT 14.97 1.4 15.11 1.765 ;
 RECT 17.045 0.71 17.185 1.765 ;
 RECT 16.1 0.71 16.24 1.765 ;
 END
 ANTENNADIFFAREA 1.132 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 24.64 2.96 ;
 RECT 2.18 2.34 2.43 2.8 ;
 RECT 7.535 2.375 7.675 2.8 ;
 RECT 14.095 2.57 14.235 2.8 ;
 RECT 15.445 2.57 15.585 2.8 ;
 RECT 13.145 2.57 13.285 2.8 ;
 RECT 5.435 2.07 5.575 2.8 ;
 RECT 11.41 2.57 11.55 2.8 ;
 RECT 10.565 2.57 10.705 2.8 ;
 RECT 16.43 2.57 16.57 2.8 ;
 RECT 0.505 1.74 0.645 2.8 ;
 RECT 1.505 1.98 1.645 2.8 ;
 END
 END VDD

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.115 1.235 7.4 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 22.925 1.41 23.265 1.775 ;
 RECT 21.245 1.965 23.11 2.105 ;
 RECT 19.015 2.195 21.385 2.335 ;
 RECT 22.97 1.775 23.11 1.965 ;
 RECT 21.245 1.41 21.385 1.965 ;
 RECT 19.015 1.365 19.155 2.195 ;
 RECT 20.4 1.345 20.54 2.195 ;
 RECT 21.245 2.105 21.385 2.195 ;
 END
 END VDDG

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 1.475 1.885 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 0.22 1.365 0.615 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 6.165 1.475 6.905 1.575 ;
 RECT 7.09 1.45 7.19 1.655 ;
 RECT 7.09 1.755 7.19 2.57 ;
 RECT 7.09 1.655 8.05 1.755 ;
 RECT 7.95 1.755 8.05 2.355 ;
 RECT 7.09 0.655 7.19 1.13 ;
 RECT 7.09 1.23 7.19 1.24 ;
 RECT 6.175 0.66 6.275 1.13 ;
 RECT 7.09 1.24 7.345 1.45 ;
 RECT 6.175 1.13 7.19 1.23 ;
 RECT 10.82 0.64 10.92 1.26 ;
 RECT 10.615 1.26 10.92 1.47 ;
 RECT 10.82 1.47 10.92 2.21 ;
 RECT 19.58 0.19 19.68 0.97 ;
 RECT 19.58 0.97 19.82 1.18 ;
 RECT 19.58 1.18 19.68 1.975 ;
 RECT 12.63 0.84 12.73 1.095 ;
 RECT 12.1 0.61 12.2 1.095 ;
 RECT 12.1 1.195 12.2 1.25 ;
 RECT 11.945 1.25 12.2 1.46 ;
 RECT 12.1 1.46 12.2 2.56 ;
 RECT 12.615 0.63 12.845 0.84 ;
 RECT 12.1 1.095 12.73 1.195 ;
 RECT 19.14 1.01 19.375 1.22 ;
 RECT 19.275 1.22 19.375 1.995 ;
 RECT 18.8 0.87 18.9 2.175 ;
 RECT 17.835 0.77 19.37 0.78 ;
 RECT 18.8 0.73 19.37 0.77 ;
 RECT 21.5 1.125 21.6 2.175 ;
 RECT 17.84 0.78 19.37 0.83 ;
 RECT 17.84 0.83 18.9 0.87 ;
 RECT 19.27 0.19 19.37 0.73 ;
 RECT 18.8 0.185 18.9 0.73 ;
 RECT 17.835 0.57 18.065 0.77 ;
 RECT 18.8 2.175 21.6 2.275 ;
 RECT 21.975 0.37 22.075 1.01 ;
 RECT 21.975 1.01 22.225 1.22 ;
 RECT 21.975 1.22 22.075 2.245 ;
 RECT 21.975 2.245 22.26 2.455 ;
 RECT 11.665 1.635 11.765 1.66 ;
 RECT 11.665 1.66 11.92 1.87 ;
 RECT 11.665 1.87 11.765 2.565 ;
 RECT 7.985 0.655 8.085 1.24 ;
 RECT 7.855 1.24 8.085 1.475 ;
 RECT 1.765 0.57 1.865 1.495 ;
 RECT 1.57 1.495 1.865 1.745 ;
 RECT 1.765 1.745 1.865 2.37 ;
 RECT 18.04 1.075 18.325 1.305 ;
 RECT 18.04 1.305 18.14 2.64 ;
 RECT 21.665 0.19 21.765 0.94 ;
 RECT 21.665 0.09 22.775 0.19 ;
 RECT 22.675 0.19 22.775 2.64 ;
 RECT 18.04 2.64 22.775 2.74 ;
 RECT 5.525 1.61 5.79 1.82 ;
 RECT 5.69 1.82 5.79 2.49 ;
 RECT 5.32 0.66 5.42 1.51 ;
 RECT 5.32 1.51 5.79 1.61 ;
 RECT 16.83 0.31 16.93 1.285 ;
 RECT 17.125 0.31 17.355 0.435 ;
 RECT 16.83 0.21 17.36 0.31 ;
 RECT 15.225 1.2 15.525 1.285 ;
 RECT 15.225 1.285 16.935 1.385 ;
 RECT 15.225 1.385 15.525 1.435 ;
 RECT 16.21 1.385 16.31 2.625 ;
 RECT 16.355 0.525 16.455 1.285 ;
 RECT 15.715 1.385 15.815 2.625 ;
 RECT 16.685 1.385 16.785 2.625 ;
 RECT 15.885 0.52 15.985 1.285 ;
 RECT 15.225 0.525 15.325 1.2 ;
 RECT 15.225 1.435 15.325 2.625 ;
 RECT 5.22 1.79 5.32 2.465 ;
 RECT 5.005 2.465 5.32 2.71 ;
 RECT 3.96 1.475 4.27 1.71 ;
 RECT 3.96 0.65 4.06 1.475 ;
 RECT 3.96 1.71 4.06 2.475 ;
 RECT 8.38 2.69 10.03 2.695 ;
 RECT 9.855 2.54 10.03 2.69 ;
 RECT 9.17 2.695 10.03 2.79 ;
 RECT 8.38 0.655 8.48 2.595 ;
 RECT 8.38 2.595 9.27 2.69 ;
 RECT 9.855 2.33 10.085 2.54 ;
 RECT 2.605 0.57 2.705 1.52 ;
 RECT 2.54 1.62 2.64 2.395 ;
 RECT 3.47 0.705 3.57 1.255 ;
 RECT 3.47 0.57 3.755 0.705 ;
 RECT 2.605 0.47 3.755 0.57 ;
 RECT 2.105 1.44 2.35 1.52 ;
 RECT 2.105 1.62 2.35 1.69 ;
 RECT 2.105 1.52 2.705 1.62 ;
 RECT 2.54 2.395 2.92 2.705 ;
 RECT 1.05 0.27 1.39 0.52 ;
 RECT 1.29 0.52 1.39 2.465 ;
 RECT 13.885 1.5 13.985 2.275 ;
 RECT 12.605 0.29 13.575 0.39 ;
 RECT 13.475 0.39 13.575 1.4 ;
 RECT 12.605 0.22 12.835 0.29 ;
 RECT 12.605 0.39 12.835 0.43 ;
 RECT 13.955 0.37 14.055 1.4 ;
 RECT 13.41 1.5 13.51 2.275 ;
 RECT 12.935 1.4 14.45 1.5 ;
 RECT 12.935 1.5 13.035 2.275 ;
 RECT 14.35 1.5 14.45 2.275 ;
 RECT 9.415 0.19 9.515 1.29 ;
 RECT 9.415 1.29 10.32 1.39 ;
 RECT 4.66 0.19 4.76 2.655 ;
 RECT 3.425 1.665 3.525 2.655 ;
 RECT 10.09 1.39 10.32 1.82 ;
 RECT 2.885 1.35 3.13 1.565 ;
 RECT 4.66 0.09 9.515 0.19 ;
 RECT 3.425 2.655 4.76 2.755 ;
 RECT 2.885 1.565 3.525 1.665 ;
 RECT 20.49 0.355 20.59 0.985 ;
 RECT 20.66 1.215 20.76 1.815 ;
 RECT 20.1 1.115 20.76 1.215 ;
 RECT 20.49 0.255 21.225 0.355 ;
 RECT 20.995 0.355 21.225 0.465 ;
 RECT 20.1 0.985 20.59 1.115 ;
 RECT 5.71 0.47 5.895 0.5 ;
 RECT 9.45 1.71 9.55 2.445 ;
 RECT 8.765 0.47 9 0.59 ;
 RECT 8.9 0.59 9 1.61 ;
 RECT 5.665 0.5 5.895 0.71 ;
 RECT 8.9 1.61 9.55 1.71 ;
 RECT 5.71 0.37 9 0.47 ;
 RECT 9.955 0.09 11.77 0.19 ;
 RECT 11.67 0.19 11.77 1.18 ;
 RECT 9.955 0.19 10.185 0.45 ;
 RECT 6.165 1.575 6.265 2.485 ;
 RECT 6.675 1.41 6.905 1.475 ;
 RECT 6.675 1.575 6.905 1.62 ;
 LAYER CO ;
 RECT 16.105 0.79 16.235 0.92 ;
 RECT 5.91 2.015 6.04 2.145 ;
 RECT 5.91 0.93 6.04 1.06 ;
 RECT 16.435 2.64 16.565 2.77 ;
 RECT 12.655 0.26 12.785 0.39 ;
 RECT 6.725 1.45 6.855 1.58 ;
 RECT 9.905 2.37 10.035 2.5 ;
 RECT 20.15 1.025 20.28 1.155 ;
 RECT 7.165 1.28 7.295 1.41 ;
 RECT 10.665 1.3 10.795 1.43 ;
 RECT 22.045 1.05 22.175 1.18 ;
 RECT 12.665 0.67 12.795 0.8 ;
 RECT 10.14 1.65 10.27 1.78 ;
 RECT 21.045 0.295 21.175 0.425 ;
 RECT 5.715 0.54 5.845 0.67 ;
 RECT 19.64 1.01 19.77 1.14 ;
 RECT 11.995 1.29 12.125 1.42 ;
 RECT 19.19 1.05 19.32 1.18 ;
 RECT 17.885 0.61 18.015 0.74 ;
 RECT 2.94 1.445 3.07 1.575 ;
 RECT 22.08 2.285 22.21 2.415 ;
 RECT 17.175 0.265 17.305 0.395 ;
 RECT 11.74 1.7 11.87 1.83 ;
 RECT 18.145 1.135 18.275 1.265 ;
 RECT 2.675 2.485 2.805 2.615 ;
 RECT 13.635 1.71 13.765 1.84 ;
 RECT 2.165 1.495 2.295 1.625 ;
 RECT 13.225 0.95 13.355 1.08 ;
 RECT 4.9 0.455 5.03 0.585 ;
 RECT 18.3 0.505 18.43 0.635 ;
 RECT 1.51 2.05 1.64 2.18 ;
 RECT 22.195 0.59 22.325 0.72 ;
 RECT 13.705 0.305 13.835 0.435 ;
 RECT 8.64 1.945 8.77 2.075 ;
 RECT 14.975 1.725 15.105 1.855 ;
 RECT 9.67 1.87 9.8 2 ;
 RECT 14.975 0.77 15.105 0.9 ;
 RECT 2.825 0.905 2.955 1.035 ;
 RECT 17.05 0.78 17.18 0.91 ;
 RECT 8.64 0.875 8.77 1.005 ;
 RECT 15.45 2.64 15.58 2.77 ;
 RECT 9.165 1.9 9.295 2.03 ;
 RECT 16.58 0.78 16.71 0.91 ;
 RECT 22.195 1.44 22.325 1.57 ;
 RECT 3.575 0.525 3.705 0.655 ;
 RECT 15.95 1.77 16.08 1.9 ;
 RECT 9.165 0.595 9.295 0.725 ;
 RECT 11.04 0.96 11.17 1.09 ;
 RECT 13.15 2.64 13.28 2.77 ;
 RECT 20.235 0.11 20.365 0.24 ;
 RECT 15.355 1.25 15.485 1.38 ;
 RECT 19.02 0.11 19.15 0.24 ;
 RECT 0.475 0.33 0.605 0.46 ;
 RECT 3.175 2.105 3.305 2.235 ;
 RECT 7.73 0.62 7.86 0.75 ;
 RECT 21.25 1.465 21.38 1.595 ;
 RECT 2.76 1.825 2.89 1.955 ;
 RECT 1.51 0.79 1.64 0.92 ;
 RECT 3.69 0.88 3.82 1.01 ;
 RECT 4.09 1.525 4.22 1.655 ;
 RECT 1.04 2.115 1.17 2.245 ;
 RECT 6.84 1.885 6.97 2.015 ;
 RECT 6.395 0.88 6.525 1.01 ;
 RECT 11.04 1.705 11.17 1.835 ;
 RECT 1.985 1.995 2.115 2.125 ;
 RECT 16.91 1.77 17.04 1.9 ;
 RECT 20.715 0.59 20.845 0.72 ;
 RECT 11.415 2.64 11.545 2.77 ;
 RECT 15.635 0.77 15.765 0.9 ;
 RECT 3.22 0.88 3.35 1.01 ;
 RECT 22.975 1.45 23.105 1.58 ;
 RECT 2.25 2.345 2.38 2.475 ;
 RECT 1.11 0.325 1.24 0.455 ;
 RECT 2.255 0.21 2.385 0.34 ;
 RECT 19.8 1.46 19.93 1.59 ;
 RECT 5.44 2.135 5.57 2.265 ;
 RECT 19.8 0.41 19.93 0.54 ;
 RECT 10.57 2.64 10.7 2.77 ;
 RECT 11.42 0.33 11.55 0.46 ;
 RECT 10.345 0.955 10.475 1.085 ;
 RECT 14.235 0.96 14.365 1.09 ;
 RECT 7.54 2.445 7.67 2.575 ;
 RECT 4.18 2.125 4.31 2.255 ;
 RECT 5.045 2.515 5.175 2.645 ;
 RECT 1.04 0.79 1.17 0.92 ;
 RECT 12.32 0.83 12.45 0.96 ;
 RECT 20.88 1.38 21.01 1.51 ;
 RECT 20.405 1.42 20.535 1.55 ;
 RECT 6.84 0.88 6.97 1.01 ;
 RECT 3.67 2.07 3.8 2.2 ;
 RECT 0.51 2.085 0.64 2.215 ;
 RECT 9.67 0.595 9.8 0.725 ;
 RECT 12.685 1.71 12.815 1.84 ;
 RECT 14.57 1.71 14.7 1.84 ;
 RECT 12.32 1.78 12.45 1.91 ;
 RECT 0.51 2.345 0.64 2.475 ;
 RECT 7.905 1.28 8.035 1.41 ;
 RECT 18.55 1.4 18.68 1.53 ;
 RECT 5.58 1.63 5.71 1.76 ;
 RECT 19.02 1.45 19.15 1.58 ;
 RECT 21.415 0.115 21.545 0.245 ;
 RECT 2.115 0.88 2.245 1.01 ;
 RECT 4.97 2.125 5.1 2.255 ;
 RECT 14.1 2.64 14.23 2.77 ;
 RECT 6.395 2.07 6.525 2.2 ;
 RECT 0.475 0.59 0.605 0.72 ;
 RECT 1.63 1.55 1.76 1.68 ;
 RECT 0.51 1.825 0.64 1.955 ;
 RECT 8.815 0.42 8.945 0.55 ;
 RECT 10.005 0.28 10.135 0.41 ;
 LAYER M1 ;
 RECT 4.63 1.44 4.77 1.52 ;
 RECT 4.02 1.52 4.77 1.66 ;
 RECT 5.905 0.865 6.045 1.3 ;
 RECT 4.63 1.3 6.045 1.44 ;
 RECT 5.905 1.44 6.045 2.215 ;
 RECT 4.07 2.12 5.17 2.26 ;
 RECT 6.39 0.82 6.53 2.225 ;
 RECT 7.24 2.165 7.38 2.225 ;
 RECT 6.39 2.225 7.38 2.365 ;
 RECT 8.635 0.765 8.775 2.025 ;
 RECT 9.16 0.525 9.3 2.025 ;
 RECT 7.24 2.025 9.3 2.165 ;
 RECT 6.835 1.62 6.975 1.735 ;
 RECT 6.835 1.875 6.975 2.085 ;
 RECT 6.835 0.81 6.975 1.41 ;
 RECT 6.675 1.41 6.975 1.62 ;
 RECT 7.585 1.415 7.725 1.735 ;
 RECT 6.835 1.735 7.725 1.875 ;
 RECT 7.585 1.275 8.105 1.415 ;
 RECT 20.115 0.705 20.255 0.985 ;
 RECT 19.795 0.33 19.935 0.565 ;
 RECT 20.1 1.195 20.24 1.32 ;
 RECT 19.795 1.46 19.935 1.735 ;
 RECT 19.795 0.565 20.255 0.705 ;
 RECT 19.795 1.32 20.24 1.46 ;
 RECT 20.1 0.985 20.33 1.195 ;
 RECT 10.62 0.805 10.76 1.26 ;
 RECT 10.615 1.26 10.845 1.3 ;
 RECT 10.615 1.44 10.845 1.47 ;
 RECT 9.665 1.3 10.845 1.44 ;
 RECT 9.665 0.525 9.805 1.3 ;
 RECT 9.665 1.44 9.805 2.065 ;
 RECT 12.315 0.43 12.455 0.665 ;
 RECT 10.62 0.665 12.455 0.805 ;
 RECT 12.315 0.805 12.455 1.98 ;
 RECT 12.315 0.22 12.835 0.43 ;
 RECT 12.615 0.72 12.845 0.84 ;
 RECT 14.11 0.37 14.25 0.58 ;
 RECT 12.615 0.58 14.25 0.72 ;
 RECT 15.35 0.37 15.49 1.46 ;
 RECT 14.11 0.23 15.49 0.37 ;
 RECT 21.085 0.465 21.225 0.685 ;
 RECT 20.995 0.255 21.225 0.465 ;
 RECT 22.505 0.825 22.645 1.36 ;
 RECT 21.085 0.685 22.645 0.825 ;
 RECT 22.19 1.5 22.33 1.705 ;
 RECT 22.19 0.485 22.33 0.685 ;
 RECT 22.19 1.36 22.645 1.5 ;
 RECT 11.035 1.095 11.175 1.255 ;
 RECT 11.035 1.255 12.175 1.395 ;
 RECT 11.035 1.395 11.175 1.7 ;
 RECT 11.945 1.25 12.175 1.255 ;
 RECT 11.945 1.395 12.175 1.46 ;
 RECT 10.97 1.7 11.245 1.84 ;
 RECT 10.965 0.955 11.235 1.095 ;
 RECT 2.82 1.615 2.96 1.82 ;
 RECT 2.82 0.795 2.96 1.405 ;
 RECT 2.82 1.405 3.12 1.615 ;
 RECT 2.69 1.82 2.96 1.96 ;
 RECT 9.855 2.42 10.085 2.54 ;
 RECT 9.855 2.28 17.715 2.42 ;
 RECT 17.575 2.42 17.715 2.505 ;
 RECT 22.03 2.455 22.17 2.505 ;
 RECT 17.575 2.505 22.17 2.645 ;
 RECT 22.03 2.245 22.26 2.455 ;
 RECT 17.125 0.36 17.355 0.435 ;
 RECT 18.65 0.36 18.79 0.54 ;
 RECT 17.115 0.22 18.79 0.36 ;
 RECT 19.515 0.97 19.82 1.18 ;
 RECT 19.515 0.68 19.655 0.97 ;
 RECT 18.65 0.54 19.655 0.68 ;
 RECT 19.515 0.535 19.655 0.54 ;
 RECT 20.71 0.48 20.85 1.08 ;
 RECT 20.875 1.22 21.015 1.58 ;
 RECT 21.995 1.01 22.225 1.08 ;
 RECT 20.71 1.08 22.225 1.22 ;
 RECT 10.12 1.82 10.26 1.985 ;
 RECT 10.12 1.985 11.875 2.125 ;
 RECT 11.69 1.87 11.875 1.985 ;
 RECT 10.09 1.61 10.32 1.82 ;
 RECT 11.69 1.66 11.92 1.87 ;
 RECT 3.505 0.52 4.105 0.66 ;
 RECT 3.965 0.66 4.105 1.015 ;
 RECT 5.51 0.505 5.895 0.71 ;
 RECT 3.965 1.015 5.65 1.155 ;
 RECT 5.665 0.5 5.895 0.505 ;
 RECT 5.51 0.71 5.65 1.015 ;
 RECT 18.37 0.64 18.51 0.99 ;
 RECT 18.095 1.17 18.685 1.2 ;
 RECT 18.095 0.99 18.545 1.03 ;
 RECT 18.545 1.2 18.685 1.725 ;
 RECT 18.095 1.2 18.325 1.305 ;
 RECT 18.25 0.5 18.51 0.64 ;
 RECT 19.14 1.01 19.37 1.03 ;
 RECT 18.095 1.03 19.37 1.17 ;
 RECT 19.14 1.17 19.37 1.22 ;
 RECT 0.815 0.925 0.955 1.195 ;
 RECT 0.815 1.335 0.955 2.11 ;
 RECT 0.815 0.785 1.24 0.925 ;
 RECT 0.815 2.11 1.24 2.25 ;
 RECT 0.815 1.195 1.925 1.335 ;
 RECT 1.785 0.67 1.925 1.195 ;
 RECT 3.215 0.36 3.355 0.9 ;
 RECT 3.29 1.08 3.43 1.945 ;
 RECT 2.53 0.22 3.355 0.36 ;
 RECT 3.17 2.17 3.31 2.305 ;
 RECT 3.17 1.945 3.43 2.17 ;
 RECT 3.215 0.9 3.43 1.08 ;
 RECT 2.53 0.36 2.67 0.53 ;
 RECT 1.785 0.53 2.67 0.67 ;
 RECT 2.025 1.63 2.165 1.99 ;
 RECT 2.025 1.475 2.37 1.63 ;
 RECT 2.11 0.81 2.25 1.475 ;
 RECT 1.915 1.99 2.165 2.13 ;
 RECT 4.95 1.79 5.09 1.82 ;
 RECT 3.685 0.805 3.825 1.82 ;
 RECT 3.595 1.96 3.875 2.215 ;
 RECT 3.595 1.82 5.09 1.96 ;
 RECT 5.525 1.58 5.765 1.65 ;
 RECT 4.95 1.65 5.765 1.79 ;
 RECT 5.525 1.79 5.765 1.835 ;
 RECT 2.575 2.41 2.91 2.51 ;
 RECT 2.575 2.65 2.91 2.66 ;
 RECT 2.575 2.51 5.295 2.65 ;
 RECT 9.955 0.38 10.185 0.45 ;
 RECT 8.765 0.38 8.995 0.59 ;
 RECT 8.765 0.24 10.2 0.38 ;
 END
END RDFFSRX2

MACRO LSDNENCLX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.36 BY 5.76 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.02 2.17 5.38 2.55 ;
 END
 ANTENNAGATEAREA 0.36 ;
 END ENB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 2.24 2.8 7.36 2.96 ;
 RECT 4.385 2.96 4.525 3.72 ;
 RECT 3.075 2.96 3.215 3.705 ;
 RECT 6.615 2.96 6.755 3.745 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.065 3.85 3.385 4.24 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END D

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 7.36 5.2 ;
 RECT 1.885 4.225 2.025 5.04 ;
 RECT 1.37 4 1.51 5.04 ;
 END
 END VDDH

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.36 0.08 ;
 RECT 3.405 0.08 3.545 2.195 ;
 RECT 5.455 0.08 5.595 1.03 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 7.36 5.84 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.03 3.88 4.995 4.02 ;
 RECT 3.85 3.515 4.17 3.655 ;
 RECT 4.855 3.2 6.285 3.34 ;
 RECT 5.815 3.34 6.285 3.425 ;
 RECT 5.815 3.105 6.285 3.2 ;
 RECT 4.03 3.655 4.17 3.88 ;
 RECT 4.855 3.34 4.995 3.88 ;
 END
 ANTENNADIFFAREA 0.864 ;
 END Q

 OBS
 LAYER PO ;
 RECT 3.33 4.1 3.43 4.67 ;
 RECT 2.14 3.8 2.24 4.67 ;
 RECT 3.33 3.275 3.43 3.87 ;
 RECT 3.085 3.87 3.43 4.1 ;
 RECT 2.14 4.67 3.43 4.77 ;
 RECT 4.17 2.26 4.27 3.11 ;
 RECT 4.64 0.39 4.74 2.16 ;
 RECT 4.17 0.39 4.27 2.16 ;
 RECT 4.17 2.16 4.74 2.26 ;
 RECT 3.95 3.11 4.27 3.34 ;
 RECT 4.17 3.34 4.27 3.97 ;
 RECT 6 2.645 6.1 3.11 ;
 RECT 6 2.415 6.23 2.645 ;
 RECT 5.945 3.11 6.175 3.34 ;
 RECT 5.075 2.275 5.335 2.455 ;
 RECT 4.64 2.555 4.74 4.05 ;
 RECT 5.715 0.39 5.815 2.455 ;
 RECT 5.235 0.39 5.335 2.275 ;
 RECT 4.64 2.455 5.815 2.555 ;
 LAYER CO ;
 RECT 6.05 2.465 6.18 2.595 ;
 RECT 3.92 3.52 4.05 3.65 ;
 RECT 3.08 3.525 3.21 3.655 ;
 RECT 3.135 3.92 3.265 4.05 ;
 RECT 3.55 3.525 3.68 3.655 ;
 RECT 1.89 4.3 2.02 4.43 ;
 RECT 6.62 3.545 6.75 3.675 ;
 RECT 2.36 4.15 2.49 4.28 ;
 RECT 4.86 3.52 4.99 3.65 ;
 RECT 6.62 3.285 6.75 3.415 ;
 RECT 1.375 4.07 1.505 4.2 ;
 RECT 4.39 3.52 4.52 3.65 ;
 RECT 1.375 4.33 1.505 4.46 ;
 RECT 3.41 1.475 3.54 1.605 ;
 RECT 3.41 1.735 3.54 1.865 ;
 RECT 3.41 1.995 3.54 2.125 ;
 RECT 4 3.16 4.13 3.29 ;
 RECT 5.995 3.16 6.125 3.29 ;
 RECT 6.04 0.975 6.17 1.105 ;
 RECT 6.04 1.26 6.17 1.39 ;
 RECT 5.46 0.82 5.59 0.95 ;
 RECT 4.89 1.26 5.02 1.39 ;
 RECT 4.89 0.975 5.02 1.105 ;
 RECT 4.39 1.59 4.52 1.72 ;
 RECT 4.39 1.305 4.52 1.435 ;
 RECT 3.86 0.945 3.99 1.075 ;
 RECT 3.86 1.21 3.99 1.34 ;
 RECT 3.86 1.485 3.99 1.615 ;
 RECT 5.125 2.315 5.255 2.445 ;
 LAYER M1 ;
 RECT 4.885 1.095 5.025 1.185 ;
 RECT 4.885 1.325 5.025 1.46 ;
 RECT 4.885 0.905 5.025 0.955 ;
 RECT 3.855 0.875 3.995 0.955 ;
 RECT 3.855 1.095 3.995 1.685 ;
 RECT 3.855 0.955 5.025 1.095 ;
 RECT 4.885 1.185 6.175 1.325 ;
 RECT 6.035 0.9 6.175 1.185 ;
 RECT 6.035 1.325 6.175 1.46 ;
 RECT 4.385 1.235 4.525 1.65 ;
 RECT 6.02 1.79 6.16 2.395 ;
 RECT 4.385 1.65 6.16 1.79 ;
 RECT 5.98 2.395 6.25 2.65 ;
 RECT 2.355 4.045 2.495 4.41 ;
 RECT 3.545 3.36 3.685 4.41 ;
 RECT 2.355 4.41 3.685 4.55 ;
 RECT 3.93 3.1 4.2 3.22 ;
 RECT 3.545 3.22 4.2 3.36 ;
 END
END LSDNENCLX1

MACRO LSDNENCLX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 12.8 BY 5.76 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.02 2.17 5.38 2.55 ;
 END
 ANTENNAGATEAREA 0.31 ;
 END ENB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 12.8 2.96 ;
 RECT 4.385 2.96 4.525 3.72 ;
 RECT 3.075 2.96 3.215 3.705 ;
 RECT 6.65 2.96 6.79 3.745 ;
 RECT 7.29 2.96 7.43 3.69 ;
 RECT 9.635 2.96 9.775 3.69 ;
 RECT 10.95 2.96 11.09 3.69 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.065 3.89 3.385 4.28 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END D

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 12.8 5.2 ;
 RECT 1.885 4.21 2.025 5.04 ;
 RECT 1.375 4 1.515 5.04 ;
 END
 END VDDH

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 12.8 0.08 ;
 RECT 3.405 0.08 3.545 2.195 ;
 RECT 5.455 0.08 5.595 1.03 ;
 RECT 7.075 0.08 7.215 1.845 ;
 RECT 8.46 0.08 8.6 1.845 ;
 RECT 9.59 0.08 9.73 1.845 ;
 RECT 10.975 0.08 11.115 1.845 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 12.8 5.84 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.75 3.12 12.11 3.455 ;
 RECT 10.265 4.025 12 4.165 ;
 RECT 11.86 3.455 12 4.025 ;
 RECT 10.265 3.265 10.405 4.025 ;
 END
 ANTENNADIFFAREA 1.354 ;
 END Q

 OBS
 LAYER PO ;
 RECT 3.33 4.14 3.43 4.67 ;
 RECT 2.14 3.8 2.24 4.67 ;
 RECT 3.33 3.275 3.43 3.91 ;
 RECT 3.085 3.91 3.43 4.14 ;
 RECT 2.14 4.67 3.43 4.77 ;
 RECT 6.31 2.11 8.215 2.21 ;
 RECT 6.31 2.21 6.41 2.415 ;
 RECT 8.115 0.355 8.215 2.11 ;
 RECT 7.385 0.355 7.485 2.11 ;
 RECT 7.665 2.21 7.765 4.05 ;
 RECT 6.31 2.645 6.41 3.11 ;
 RECT 6.255 3.11 6.485 3.34 ;
 RECT 6.31 2.415 6.54 2.645 ;
 RECT 4.17 0.535 4.27 2.16 ;
 RECT 4.17 2.16 4.74 2.26 ;
 RECT 4.17 2.26 4.27 3.11 ;
 RECT 4.64 0.535 4.74 2.16 ;
 RECT 3.95 3.11 4.27 3.34 ;
 RECT 4.17 3.34 4.27 3.97 ;
 RECT 11.88 2.425 11.98 3.2 ;
 RECT 11.83 2.215 12.06 2.425 ;
 RECT 11.815 3.2 12.045 3.41 ;
 RECT 8.95 2.45 9.05 3.1 ;
 RECT 9.9 0.185 10 2.295 ;
 RECT 9.9 2.395 10 3.975 ;
 RECT 10.63 0.19 10.73 2.295 ;
 RECT 10.63 2.395 10.73 3.975 ;
 RECT 8.91 2.24 9.14 2.295 ;
 RECT 8.91 2.395 9.14 2.45 ;
 RECT 8.91 2.295 10.73 2.395 ;
 RECT 8.885 3.1 9.115 3.31 ;
 RECT 5.235 0.535 5.335 2.06 ;
 RECT 5.235 2.06 5.815 2.16 ;
 RECT 5.235 2.16 5.335 2.275 ;
 RECT 5.715 0.535 5.815 2.06 ;
 RECT 5.075 2.275 5.335 2.455 ;
 RECT 4.64 2.555 4.74 3.97 ;
 RECT 4.64 2.455 5.335 2.555 ;
 LAYER CO ;
 RECT 3.41 1.475 3.54 1.605 ;
 RECT 3.41 1.735 3.54 1.865 ;
 RECT 3.41 1.995 3.54 2.125 ;
 RECT 4 3.16 4.13 3.29 ;
 RECT 6.305 3.16 6.435 3.29 ;
 RECT 10.955 3.49 11.085 3.62 ;
 RECT 10.27 3.49 10.4 3.62 ;
 RECT 9.64 3.49 9.77 3.62 ;
 RECT 10.98 1.21 11.11 1.34 ;
 RECT 10.225 0.945 10.355 1.075 ;
 RECT 10.98 1.485 11.11 1.615 ;
 RECT 10.98 0.945 11.11 1.075 ;
 RECT 9.595 1.21 9.725 1.34 ;
 RECT 10.225 1.21 10.355 1.34 ;
 RECT 9.595 1.485 9.725 1.615 ;
 RECT 10.225 1.485 10.355 1.615 ;
 RECT 9.595 0.945 9.725 1.075 ;
 RECT 8.065 3.205 8.195 3.335 ;
 RECT 8.065 3.49 8.195 3.62 ;
 RECT 8.465 1.21 8.595 1.34 ;
 RECT 8.465 1.485 8.595 1.615 ;
 RECT 8.465 0.945 8.595 1.075 ;
 RECT 7.71 1.21 7.84 1.34 ;
 RECT 7.71 1.485 7.84 1.615 ;
 RECT 7.71 0.945 7.84 1.075 ;
 RECT 7.08 1.21 7.21 1.34 ;
 RECT 7.08 1.485 7.21 1.615 ;
 RECT 7.08 0.945 7.21 1.075 ;
 RECT 7.295 3.205 7.425 3.335 ;
 RECT 7.295 3.49 7.425 3.62 ;
 RECT 6.04 0.975 6.17 1.105 ;
 RECT 6.04 1.26 6.17 1.39 ;
 RECT 5.46 0.82 5.59 0.95 ;
 RECT 4.89 1.26 5.02 1.39 ;
 RECT 4.89 0.975 5.02 1.105 ;
 RECT 4.39 1.59 4.52 1.72 ;
 RECT 4.39 1.305 4.52 1.435 ;
 RECT 3.86 0.945 3.99 1.075 ;
 RECT 3.86 1.21 3.99 1.34 ;
 RECT 3.86 1.485 3.99 1.615 ;
 RECT 6.36 2.465 6.49 2.595 ;
 RECT 3.92 3.52 4.05 3.65 ;
 RECT 3.08 3.525 3.21 3.655 ;
 RECT 3.135 3.96 3.265 4.09 ;
 RECT 3.55 3.525 3.68 3.655 ;
 RECT 1.89 4.28 2.02 4.41 ;
 RECT 6.655 3.545 6.785 3.675 ;
 RECT 11.88 2.255 12.01 2.385 ;
 RECT 11.865 3.24 11.995 3.37 ;
 RECT 8.96 2.28 9.09 2.41 ;
 RECT 8.935 3.14 9.065 3.27 ;
 RECT 5.125 2.315 5.255 2.445 ;
 RECT 2.36 4.15 2.49 4.28 ;
 RECT 4.86 3.52 4.99 3.65 ;
 RECT 6.655 3.285 6.785 3.415 ;
 RECT 1.38 4.07 1.51 4.2 ;
 RECT 4.39 3.52 4.52 3.65 ;
 RECT 1.38 4.33 1.51 4.46 ;
 LAYER M1 ;
 RECT 4.885 1.095 5.025 1.185 ;
 RECT 4.885 1.325 5.025 1.46 ;
 RECT 4.885 0.665 5.025 0.955 ;
 RECT 3.855 0.485 3.995 0.955 ;
 RECT 3.855 1.095 3.995 2.12 ;
 RECT 3.855 0.955 5.025 1.095 ;
 RECT 4.885 1.185 6.175 1.325 ;
 RECT 6.035 0.665 6.175 1.185 ;
 RECT 6.035 1.325 6.175 1.46 ;
 RECT 2.355 4.095 2.495 4.42 ;
 RECT 3.545 3.36 3.685 4.42 ;
 RECT 3.93 3.1 4.2 3.22 ;
 RECT 3.545 3.22 4.2 3.36 ;
 RECT 2.355 4.42 3.685 4.56 ;
 RECT 4.03 3.655 4.17 3.88 ;
 RECT 3.85 3.515 4.17 3.655 ;
 RECT 4.855 3.34 4.995 3.88 ;
 RECT 6.235 3.1 6.505 3.2 ;
 RECT 6.235 3.34 6.505 3.36 ;
 RECT 4.855 3.2 6.505 3.34 ;
 RECT 4.03 3.88 4.995 4.02 ;
 RECT 4.385 1.235 4.525 1.65 ;
 RECT 6.33 1.79 6.47 2.395 ;
 RECT 4.385 1.65 6.47 1.79 ;
 RECT 6.29 2.395 6.56 2.655 ;
 RECT 10.22 0.855 10.36 2.235 ;
 RECT 11.83 2.215 12.06 2.235 ;
 RECT 11.83 2.375 12.06 2.425 ;
 RECT 10.22 2.235 12.06 2.375 ;
 RECT 7.705 0.855 7.845 2.235 ;
 RECT 7.705 2.24 9.14 2.375 ;
 RECT 8.91 2.375 9.14 2.45 ;
 RECT 7.705 2.235 9.115 2.24 ;
 RECT 8.06 3.275 8.2 3.825 ;
 RECT 8.885 3.1 9.115 3.135 ;
 RECT 8.885 3.275 9.115 3.31 ;
 RECT 8.06 3.135 9.115 3.275 ;
 END
END LSDNENCLX2

MACRO LSDNENCLX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 13.065 BY 5.76 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.285 2.17 5.645 2.55 ;
 END
 ANTENNAGATEAREA 0.31 ;
 END ENB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 13.065 2.96 ;
 RECT 11.215 2.96 11.355 3.69 ;
 RECT 6.955 2.96 7.095 4.1 ;
 RECT 4.65 2.96 4.79 3.72 ;
 RECT 9.9 2.96 10.04 3.69 ;
 RECT 7.555 2.96 7.695 3.69 ;
 RECT 3.34 2.96 3.48 3.75 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.33 3.89 3.65 4.28 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END D

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 13.065 5.2 ;
 RECT 1.31 3.605 1.45 5.04 ;
 RECT 1.77 3.665 1.91 5.04 ;
 END
 END VDDH

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 13.065 0.08 ;
 RECT 7.34 0.08 7.48 1.845 ;
 RECT 9.855 0.08 9.995 1.845 ;
 RECT 3.67 0.08 3.81 2.195 ;
 RECT 8.725 0.08 8.865 1.845 ;
 RECT 11.24 0.08 11.38 1.845 ;
 RECT 5.72 0.08 5.86 1.03 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 13.065 5.84 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.96 3.12 12.4 3.45 ;
 RECT 10.53 4.025 12.265 4.165 ;
 RECT 12.125 3.45 12.265 4.025 ;
 RECT 10.53 3.265 10.67 4.025 ;
 END
 ANTENNADIFFAREA 1.354 ;
 END Q

 OBS
 LAYER PO ;
 RECT 3.595 3.225 3.695 3.915 ;
 RECT 3.35 3.915 3.695 4.245 ;
 RECT 2.025 3.385 2.125 4.245 ;
 RECT 2.025 4.245 3.695 4.345 ;
 RECT 12.145 2.425 12.245 3.2 ;
 RECT 12.08 3.2 12.31 3.41 ;
 RECT 12.095 2.215 12.325 2.425 ;
 RECT 9.215 2.45 9.315 3.1 ;
 RECT 9.175 2.24 9.405 2.295 ;
 RECT 9.175 2.295 10.995 2.395 ;
 RECT 9.175 2.395 9.405 2.45 ;
 RECT 10.165 0.185 10.265 2.295 ;
 RECT 10.165 2.395 10.265 3.975 ;
 RECT 10.895 0.19 10.995 2.295 ;
 RECT 10.895 2.395 10.995 3.975 ;
 RECT 9.15 3.1 9.38 3.31 ;
 RECT 5.34 2.275 5.6 2.455 ;
 RECT 5.5 2.16 5.6 2.275 ;
 RECT 5.5 0.535 5.6 2.06 ;
 RECT 5.5 2.06 6.08 2.16 ;
 RECT 5.98 0.535 6.08 2.06 ;
 RECT 4.905 2.555 5.005 4.05 ;
 RECT 4.905 2.455 5.6 2.555 ;
 RECT 4.435 2.26 4.535 3.11 ;
 RECT 4.905 0.535 5.005 2.16 ;
 RECT 4.435 0.535 4.535 2.16 ;
 RECT 4.435 2.16 5.005 2.26 ;
 RECT 4.215 3.11 4.535 3.34 ;
 RECT 4.435 3.34 4.535 3.97 ;
 RECT 6.575 2.21 6.675 2.415 ;
 RECT 6.575 2.645 6.675 3.11 ;
 RECT 6.575 2.11 8.48 2.21 ;
 RECT 8.38 0.355 8.48 2.11 ;
 RECT 7.65 0.355 7.75 2.11 ;
 RECT 7.93 2.21 8.03 4.05 ;
 RECT 6.575 2.415 6.805 2.645 ;
 RECT 6.52 3.11 6.75 3.34 ;
 LAYER CO ;
 RECT 1.775 3.735 1.905 3.865 ;
 RECT 6.96 3.9 7.09 4.03 ;
 RECT 2.245 3.735 2.375 3.865 ;
 RECT 12.13 3.24 12.26 3.37 ;
 RECT 9.225 2.28 9.355 2.41 ;
 RECT 9.2 3.14 9.33 3.27 ;
 RECT 5.39 2.315 5.52 2.445 ;
 RECT 11.22 3.49 11.35 3.62 ;
 RECT 10.535 3.49 10.665 3.62 ;
 RECT 9.905 3.49 10.035 3.62 ;
 RECT 11.245 1.21 11.375 1.34 ;
 RECT 10.49 0.945 10.62 1.075 ;
 RECT 11.245 1.485 11.375 1.615 ;
 RECT 11.245 0.945 11.375 1.075 ;
 RECT 9.86 1.21 9.99 1.34 ;
 RECT 10.49 1.21 10.62 1.34 ;
 RECT 9.86 1.485 9.99 1.615 ;
 RECT 10.49 1.485 10.62 1.615 ;
 RECT 9.86 0.945 9.99 1.075 ;
 RECT 8.33 3.205 8.46 3.335 ;
 RECT 8.33 3.49 8.46 3.62 ;
 RECT 8.73 1.21 8.86 1.34 ;
 RECT 8.73 1.485 8.86 1.615 ;
 RECT 8.73 0.945 8.86 1.075 ;
 RECT 7.975 1.21 8.105 1.34 ;
 RECT 7.975 1.485 8.105 1.615 ;
 RECT 7.975 0.945 8.105 1.075 ;
 RECT 7.345 1.21 7.475 1.34 ;
 RECT 7.345 1.485 7.475 1.615 ;
 RECT 7.345 0.945 7.475 1.075 ;
 RECT 7.56 3.205 7.69 3.335 ;
 RECT 7.56 3.49 7.69 3.62 ;
 RECT 6.305 0.975 6.435 1.105 ;
 RECT 6.305 1.26 6.435 1.39 ;
 RECT 5.725 0.82 5.855 0.95 ;
 RECT 5.155 1.26 5.285 1.39 ;
 RECT 5.155 0.975 5.285 1.105 ;
 RECT 4.655 1.59 4.785 1.72 ;
 RECT 4.655 1.305 4.785 1.435 ;
 RECT 4.125 0.945 4.255 1.075 ;
 RECT 4.125 1.21 4.255 1.34 ;
 RECT 4.125 1.485 4.255 1.615 ;
 RECT 12.145 2.255 12.275 2.385 ;
 RECT 5.125 3.52 5.255 3.65 ;
 RECT 6.96 3.64 7.09 3.77 ;
 RECT 1.315 3.675 1.445 3.805 ;
 RECT 4.655 3.52 4.785 3.65 ;
 RECT 1.315 3.935 1.445 4.065 ;
 RECT 3.675 1.475 3.805 1.605 ;
 RECT 3.675 1.735 3.805 1.865 ;
 RECT 3.675 1.995 3.805 2.125 ;
 RECT 4.265 3.16 4.395 3.29 ;
 RECT 6.57 3.16 6.7 3.29 ;
 RECT 6.625 2.465 6.755 2.595 ;
 RECT 4.185 3.52 4.315 3.65 ;
 RECT 3.345 3.525 3.475 3.655 ;
 RECT 3.4 3.96 3.53 4.09 ;
 RECT 3.815 3.525 3.945 3.655 ;
 LAYER M1 ;
 RECT 4.65 1.235 4.79 1.65 ;
 RECT 6.595 1.79 6.735 2.395 ;
 RECT 4.65 1.65 6.735 1.79 ;
 RECT 6.555 2.395 6.825 2.65 ;
 RECT 8.325 3.275 8.465 3.825 ;
 RECT 9.15 3.1 9.38 3.135 ;
 RECT 9.15 3.275 9.38 3.31 ;
 RECT 8.325 3.135 9.38 3.275 ;
 RECT 7.97 0.855 8.11 2.235 ;
 RECT 7.97 2.24 9.405 2.375 ;
 RECT 7.97 2.235 9.38 2.24 ;
 RECT 9.175 2.375 9.405 2.45 ;
 RECT 10.485 0.855 10.625 2.235 ;
 RECT 12.095 2.215 12.325 2.235 ;
 RECT 12.095 2.375 12.325 2.425 ;
 RECT 10.485 2.235 12.325 2.375 ;
 RECT 5.15 1.095 5.29 1.185 ;
 RECT 5.15 1.325 5.29 1.46 ;
 RECT 4.12 0.485 4.26 0.955 ;
 RECT 4.12 1.095 4.26 2.12 ;
 RECT 5.15 0.665 5.29 0.955 ;
 RECT 4.12 0.955 5.29 1.095 ;
 RECT 5.15 1.185 6.44 1.325 ;
 RECT 6.3 0.665 6.44 1.185 ;
 RECT 6.3 1.325 6.44 1.46 ;
 RECT 2.24 3.685 2.38 4.465 ;
 RECT 3.81 3.36 3.95 4.465 ;
 RECT 4.195 3.105 4.465 3.22 ;
 RECT 3.81 3.22 4.465 3.36 ;
 RECT 2.24 4.465 3.95 4.605 ;
 RECT 4.295 3.655 4.435 3.88 ;
 RECT 4.115 3.515 4.435 3.655 ;
 RECT 5.12 3.34 5.26 3.88 ;
 RECT 6.5 3.1 6.77 3.2 ;
 RECT 6.5 3.34 6.77 3.36 ;
 RECT 5.12 3.2 6.77 3.34 ;
 RECT 4.295 3.88 5.26 4.02 ;
 END
END LSDNENCLX4

MACRO LSDNENCLX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 15.225 BY 5.76 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.205 2.17 5.565 2.55 ;
 END
 ANTENNAGATEAREA 0.31 ;
 END ENB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 15.225 2.96 ;
 RECT 13.47 2.96 13.61 3.69 ;
 RECT 4.57 2.96 4.71 3.72 ;
 RECT 10.92 2.96 11.06 3.69 ;
 RECT 7.475 2.96 7.615 3.69 ;
 RECT 3.26 2.96 3.4 3.75 ;
 RECT 12.235 2.96 12.375 3.69 ;
 RECT 6.88 2.96 7.02 3.745 ;
 RECT 9.01 2.96 9.15 3.69 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.25 3.89 3.57 4.28 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END D

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 15.225 5.2 ;
 RECT 1.69 3.94 1.83 5.04 ;
 RECT 1.28 3.785 1.42 5.04 ;
 END
 END VDDH

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 15.225 0.08 ;
 RECT 8.645 0.08 8.785 1.845 ;
 RECT 12.26 0.08 12.4 1.845 ;
 RECT 5.64 0.08 5.78 1.03 ;
 RECT 13.495 0.08 13.635 1.845 ;
 RECT 7.26 0.08 7.4 1.845 ;
 RECT 10.875 0.08 11.015 1.845 ;
 RECT 9.825 0.08 9.965 1.845 ;
 RECT 3.59 0.08 3.73 2.195 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 15.225 5.84 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.37 3.125 14.86 3.485 ;
 RECT 11.55 4.025 14.665 4.165 ;
 RECT 14.525 3.485 14.665 4.025 ;
 RECT 11.55 3.265 11.69 4.025 ;
 RECT 12.845 3.265 12.985 4.025 ;
 END
 ANTENNADIFFAREA 2.59 ;
 END Q

 OBS
 LAYER PO ;
 RECT 5.42 0.535 5.52 2.06 ;
 RECT 5.42 2.06 6 2.16 ;
 RECT 5.42 2.16 5.52 2.275 ;
 RECT 5.9 0.535 6 2.06 ;
 RECT 5.26 2.275 5.52 2.455 ;
 RECT 4.825 2.555 4.925 4.05 ;
 RECT 4.825 2.455 5.52 2.555 ;
 RECT 14.545 2.425 14.645 3.2 ;
 RECT 14.48 3.2 14.71 3.41 ;
 RECT 14.495 2.215 14.725 2.425 ;
 RECT 4.355 0.535 4.455 2.16 ;
 RECT 4.355 2.16 4.925 2.26 ;
 RECT 4.355 2.26 4.455 3.11 ;
 RECT 4.825 0.535 4.925 2.16 ;
 RECT 4.135 3.11 4.455 3.34 ;
 RECT 4.355 3.34 4.455 3.97 ;
 RECT 1.945 4.285 3.595 4.305 ;
 RECT 1.945 4.305 3.41 4.385 ;
 RECT 3.27 4.2 3.595 4.285 ;
 RECT 1.945 3.475 2.045 4.285 ;
 RECT 3.27 3.91 3.615 4.2 ;
 RECT 3.515 3.275 3.615 3.91 ;
 RECT 9.925 2.45 10.025 3.1 ;
 RECT 9.885 2.24 10.115 2.295 ;
 RECT 9.885 2.395 10.115 2.45 ;
 RECT 9.885 2.295 13.345 2.395 ;
 RECT 13.245 0.185 13.345 2.295 ;
 RECT 13.245 2.395 13.345 3.975 ;
 RECT 12.57 0.185 12.67 2.295 ;
 RECT 12.57 2.395 12.67 3.975 ;
 RECT 11.185 0.185 11.285 2.295 ;
 RECT 11.185 2.395 11.285 3.975 ;
 RECT 11.915 0.19 12.015 2.295 ;
 RECT 11.915 2.395 12.015 3.975 ;
 RECT 9.86 3.1 10.09 3.31 ;
 RECT 6.495 2.11 9.655 2.16 ;
 RECT 6.495 2.16 9.65 2.21 ;
 RECT 6.495 2.21 6.595 2.415 ;
 RECT 6.495 2.645 6.595 3.11 ;
 RECT 8.61 2.21 8.71 4.05 ;
 RECT 9.555 0.355 9.655 2.11 ;
 RECT 8.945 0.355 9.045 2.11 ;
 RECT 8.3 0.355 8.4 2.11 ;
 RECT 7.57 0.355 7.67 2.11 ;
 RECT 7.85 2.21 7.95 4.05 ;
 RECT 6.495 2.415 6.725 2.645 ;
 RECT 6.44 3.11 6.67 3.34 ;
 LAYER CO ;
 RECT 6.49 3.16 6.62 3.29 ;
 RECT 13.475 3.49 13.605 3.62 ;
 RECT 12.85 3.49 12.98 3.62 ;
 RECT 13.5 1.21 13.63 1.34 ;
 RECT 13.5 1.485 13.63 1.615 ;
 RECT 13.5 0.945 13.63 1.075 ;
 RECT 12.865 0.945 12.995 1.075 ;
 RECT 12.865 1.21 12.995 1.34 ;
 RECT 12.865 1.485 12.995 1.615 ;
 RECT 9.015 3.205 9.145 3.335 ;
 RECT 9.015 3.49 9.145 3.62 ;
 RECT 9.83 1.485 9.96 1.615 ;
 RECT 9.83 0.945 9.96 1.075 ;
 RECT 9.83 1.21 9.96 1.34 ;
 RECT 9.27 1.21 9.4 1.34 ;
 RECT 9.27 1.485 9.4 1.615 ;
 RECT 9.27 0.945 9.4 1.075 ;
 RECT 12.24 3.49 12.37 3.62 ;
 RECT 11.555 3.49 11.685 3.62 ;
 RECT 10.925 3.49 11.055 3.62 ;
 RECT 12.265 1.21 12.395 1.34 ;
 RECT 11.51 0.945 11.64 1.075 ;
 RECT 12.265 1.485 12.395 1.615 ;
 RECT 12.265 0.945 12.395 1.075 ;
 RECT 10.88 1.21 11.01 1.34 ;
 RECT 11.51 1.21 11.64 1.34 ;
 RECT 10.88 1.485 11.01 1.615 ;
 RECT 11.51 1.485 11.64 1.615 ;
 RECT 10.88 0.945 11.01 1.075 ;
 RECT 8.25 3.205 8.38 3.335 ;
 RECT 8.25 3.49 8.38 3.62 ;
 RECT 8.65 1.21 8.78 1.34 ;
 RECT 8.65 1.485 8.78 1.615 ;
 RECT 8.65 0.945 8.78 1.075 ;
 RECT 7.895 1.21 8.025 1.34 ;
 RECT 7.895 1.485 8.025 1.615 ;
 RECT 7.895 0.945 8.025 1.075 ;
 RECT 7.265 1.21 7.395 1.34 ;
 RECT 7.265 1.485 7.395 1.615 ;
 RECT 7.265 0.945 7.395 1.075 ;
 RECT 7.48 3.205 7.61 3.335 ;
 RECT 7.48 3.49 7.61 3.62 ;
 RECT 1.285 4.115 1.415 4.245 ;
 RECT 3.595 1.475 3.725 1.605 ;
 RECT 3.595 1.735 3.725 1.865 ;
 RECT 3.595 1.995 3.725 2.125 ;
 RECT 4.185 3.16 4.315 3.29 ;
 RECT 6.225 0.975 6.355 1.105 ;
 RECT 6.225 1.26 6.355 1.39 ;
 RECT 5.645 0.82 5.775 0.95 ;
 RECT 5.075 1.26 5.205 1.39 ;
 RECT 5.075 0.975 5.205 1.105 ;
 RECT 4.575 1.59 4.705 1.72 ;
 RECT 4.575 1.305 4.705 1.435 ;
 RECT 4.045 0.945 4.175 1.075 ;
 RECT 4.045 1.21 4.175 1.34 ;
 RECT 4.045 1.485 4.175 1.615 ;
 RECT 5.31 2.315 5.44 2.445 ;
 RECT 14.53 3.24 14.66 3.37 ;
 RECT 9.935 2.28 10.065 2.41 ;
 RECT 9.91 3.14 10.04 3.27 ;
 RECT 14.545 2.255 14.675 2.385 ;
 RECT 6.545 2.465 6.675 2.595 ;
 RECT 4.105 3.52 4.235 3.65 ;
 RECT 3.265 3.525 3.395 3.655 ;
 RECT 3.32 3.96 3.45 4.09 ;
 RECT 3.735 3.525 3.865 3.655 ;
 RECT 1.695 4.015 1.825 4.145 ;
 RECT 6.885 3.545 7.015 3.675 ;
 RECT 2.165 3.825 2.295 3.955 ;
 RECT 5.045 3.52 5.175 3.65 ;
 RECT 6.885 3.285 7.015 3.415 ;
 RECT 1.285 3.855 1.415 3.985 ;
 RECT 4.575 3.52 4.705 3.65 ;
 LAYER M1 ;
 RECT 5.07 1.095 5.21 1.185 ;
 RECT 5.07 1.325 5.21 1.46 ;
 RECT 5.07 0.665 5.21 0.955 ;
 RECT 4.04 0.485 4.18 0.955 ;
 RECT 4.04 1.095 4.18 2.12 ;
 RECT 4.04 0.955 5.21 1.095 ;
 RECT 5.07 1.185 6.36 1.325 ;
 RECT 6.22 0.665 6.36 1.185 ;
 RECT 6.22 1.325 6.36 1.46 ;
 RECT 9.265 0.855 9.405 2.235 ;
 RECT 7.89 0.855 8.03 2.235 ;
 RECT 9.885 2.375 10.115 2.45 ;
 RECT 7.89 2.235 10.115 2.375 ;
 RECT 8.245 3.155 8.385 3.855 ;
 RECT 8.245 3.855 10.045 3.995 ;
 RECT 9.905 3.31 10.045 3.855 ;
 RECT 9.86 3.1 10.09 3.31 ;
 RECT 12.86 0.855 13 2.235 ;
 RECT 11.505 0.855 11.645 2.235 ;
 RECT 14.38 2.145 14.82 2.235 ;
 RECT 14.38 2.375 14.82 2.5 ;
 RECT 11.505 2.235 14.82 2.375 ;
 RECT 4.57 1.235 4.71 1.65 ;
 RECT 6.515 1.79 6.655 2.395 ;
 RECT 4.57 1.65 6.655 1.79 ;
 RECT 6.475 2.395 6.745 2.655 ;
 RECT 2.16 3.775 2.3 4.505 ;
 RECT 3.73 3.36 3.87 4.505 ;
 RECT 4.115 3.1 4.385 3.22 ;
 RECT 3.73 3.22 4.385 3.36 ;
 RECT 2.16 4.505 3.87 4.645 ;
 RECT 4.215 3.655 4.355 3.88 ;
 RECT 4.035 3.515 4.355 3.655 ;
 RECT 5.04 3.34 5.18 3.88 ;
 RECT 6.42 3.105 6.69 3.2 ;
 RECT 6.42 3.34 6.69 3.36 ;
 RECT 5.04 3.2 6.69 3.34 ;
 RECT 4.215 3.88 5.18 4.02 ;
 END
END LSDNENCLX8

MACRO LSDNENX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.36 BY 5.76 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.67 3.955 4.04 4.29 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.36 2.96 ;
 RECT 0.325 2.96 0.465 3.745 ;
 RECT 1.61 3.515 2.245 3.655 ;
 RECT 0.835 2.96 0.975 3.75 ;
 RECT 3.86 2.96 4 3.735 ;
 RECT 2.105 2.96 2.245 3.515 ;
 END
 END VSS

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.825 3.89 1.145 4.19 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END ENB

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 7.36 5.2 ;
 RECT 5.835 3.855 5.975 5.04 ;
 RECT 5.425 3.945 5.565 5.04 ;
 END
 END VDDH

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.36 0.08 ;
 RECT 0.74 1.48 1.06 1.62 ;
 RECT 0.5 0.08 0.64 1.115 ;
 RECT 2.145 0.08 2.285 1.675 ;
 RECT 0.74 1.62 0.88 1.955 ;
 RECT 0.92 0.08 1.06 1.48 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 7.36 5.84 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.675 1.87 2.755 2.01 ;
 RECT 2.615 2.395 2.93 2.66 ;
 RECT 1.675 1.13 1.815 1.87 ;
 RECT 2.615 2.01 2.755 2.395 ;
 RECT 2.615 1.09 2.755 1.87 ;
 END
 ANTENNADIFFAREA 0.764 ;
 END Q

 OBS
 LAYER PO ;
 RECT 2.4 0.795 2.5 3.95 ;
 RECT 2.4 3.95 2.63 4.16 ;
 RECT 1.09 2.34 1.19 3.91 ;
 RECT 0.845 3.91 1.19 4.14 ;
 RECT 1.09 4.14 1.19 4.21 ;
 RECT 0.995 1.35 1.095 2.24 ;
 RECT 0.995 2.24 1.19 2.34 ;
 RECT 5.2 3.32 5.3 4.545 ;
 RECT 3.645 3.315 3.745 3.975 ;
 RECT 5.2 3.315 5.31 3.32 ;
 RECT 3.645 3.975 3.93 4.205 ;
 RECT 3.645 4.205 3.745 4.295 ;
 RECT 3.645 3.215 5.31 3.315 ;
 RECT 1.93 2.585 2.03 3.11 ;
 RECT 1.685 2.35 2.03 2.355 ;
 RECT 1.67 2.355 2.03 2.585 ;
 RECT 1.93 0.785 2.03 2.35 ;
 RECT 1.71 3.11 2.03 3.34 ;
 RECT 1.93 3.34 2.03 4.045 ;
 RECT 2.68 2.645 2.78 3.11 ;
 RECT 2.68 2.415 2.91 2.645 ;
 RECT 2.68 3.11 2.91 3.34 ;
 LAYER CO ;
 RECT 3.73 4.025 3.86 4.155 ;
 RECT 1.68 1.48 1.81 1.61 ;
 RECT 1.31 3.525 1.44 3.655 ;
 RECT 1.215 1.755 1.345 1.885 ;
 RECT 0.745 1.755 0.875 1.885 ;
 RECT 5.84 3.925 5.97 4.055 ;
 RECT 2.62 1.21 2.75 1.34 ;
 RECT 0.84 3.525 0.97 3.655 ;
 RECT 5.84 4.185 5.97 4.315 ;
 RECT 2.62 3.52 2.75 3.65 ;
 RECT 0.895 3.96 1.025 4.09 ;
 RECT 1.68 3.52 1.81 3.65 ;
 RECT 2.62 1.485 2.75 1.615 ;
 RECT 1.68 1.2 1.81 1.33 ;
 RECT 0.33 3.545 0.46 3.675 ;
 RECT 0.33 3.285 0.46 3.415 ;
 RECT 1.68 1.75 1.81 1.88 ;
 RECT 2.45 3.99 2.58 4.12 ;
 RECT 3.39 3.51 3.52 3.64 ;
 RECT 2.15 1.48 2.28 1.61 ;
 RECT 2.15 1.2 2.28 1.33 ;
 RECT 5.43 4.1 5.56 4.23 ;
 RECT 4.945 4.1 5.075 4.23 ;
 RECT 1.72 2.405 1.85 2.535 ;
 RECT 2.73 2.465 2.86 2.595 ;
 RECT 3.865 3.515 3.995 3.645 ;
 RECT 0.505 0.395 0.635 0.525 ;
 RECT 0.505 0.655 0.635 0.785 ;
 RECT 0.505 0.915 0.635 1.045 ;
 RECT 1.76 3.16 1.89 3.29 ;
 RECT 2.73 3.16 2.86 3.29 ;
 LAYER M1 ;
 RECT 3.385 4.125 3.525 4.55 ;
 RECT 2.4 3.95 2.63 3.985 ;
 RECT 2.4 4.125 2.63 4.16 ;
 RECT 3.385 3.4 3.525 3.985 ;
 RECT 2.395 3.985 3.525 4.125 ;
 RECT 3.385 4.55 5.08 4.69 ;
 RECT 4.94 4.03 5.08 4.55 ;
 RECT 1.21 1.515 1.35 2.38 ;
 RECT 1.65 2.335 1.92 2.38 ;
 RECT 1.65 2.52 1.92 2.605 ;
 RECT 1.21 2.38 1.92 2.52 ;
 RECT 1.305 3.36 1.445 3.73 ;
 RECT 1.69 3.1 1.96 3.22 ;
 RECT 1.305 3.22 1.96 3.36 ;
 RECT 2.615 3.1 2.93 3.36 ;
 RECT 2.615 3.36 2.755 3.77 ;
 END
END LSDNENX1

MACRO LSDNENX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 5.76 ;
 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 4.8 5.2 ;
 RECT 3.345 3.795 3.485 5.04 ;
 RECT 2.93 3.735 3.07 5.04 ;
 END
 END VDDH

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 1.435 0.08 1.575 1.02 ;
 RECT 0.415 0.08 0.555 1.295 ;
 RECT 1.965 0.08 2.105 1.405 ;
 RECT 2.95 0.08 3.09 0.82 ;
 RECT 3.92 0.08 4.06 0.885 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 4.8 5.84 ;
 END
 END VDDL

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 3.375 2.635 3.65 2.8 ;
 RECT 0.84 2.96 0.98 3.715 ;
 RECT 0.51 2.96 0.65 2.985 ;
 RECT 0.51 2.735 0.65 2.8 ;
 RECT 1.43 2.245 1.57 2.8 ;
 END
 END VSS

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.24 1.42 1.615 1.76 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END ENB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.805 3.855 1.17 4.21 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.445 1.455 2.885 1.76 ;
 RECT 2.375 1.915 2.665 2.055 ;
 RECT 2.445 0.98 3.57 1.12 ;
 RECT 2.445 1.76 2.585 1.915 ;
 RECT 3.43 1.12 3.57 1.355 ;
 RECT 3.43 0.28 3.57 0.98 ;
 RECT 2.445 1.12 2.585 1.455 ;
 RECT 2.445 0.285 2.585 0.98 ;
 END
 ANTENNADIFFAREA 1.11 ;
 END Q

 OBS
 LAYER PO ;
 RECT 1.095 4.425 2.815 4.525 ;
 RECT 1.095 4.085 1.195 4.425 ;
 RECT 2.715 3.565 2.815 4.425 ;
 RECT 1.095 3.265 1.195 3.875 ;
 RECT 0.94 3.875 1.195 4.085 ;
 RECT 3.205 1.98 3.305 2.73 ;
 RECT 3.7 0.09 3.8 1.88 ;
 RECT 3.7 1.98 3.8 2.73 ;
 RECT 3.205 1.72 3.435 1.88 ;
 RECT 3.205 0.09 3.305 1.72 ;
 RECT 3.205 1.88 3.8 1.98 ;
 RECT 2.04 1.545 2.32 1.6 ;
 RECT 2.04 1.7 2.32 1.755 ;
 RECT 1.69 1.6 2.32 1.7 ;
 RECT 1.69 1.7 1.79 3.88 ;
 RECT 2.22 0.19 2.32 1.545 ;
 RECT 2.715 0.19 2.815 2.715 ;
 RECT 2.22 1.755 2.32 2.72 ;
 RECT 1.38 3.88 1.835 4.09 ;
 RECT 2.22 0.09 2.815 0.19 ;
 RECT 1.21 0.205 1.31 1.55 ;
 RECT 1.21 1.76 1.31 2.695 ;
 RECT 1.21 1.55 1.47 1.76 ;
 LAYER CO ;
 RECT 3.445 2.64 3.575 2.77 ;
 RECT 2.45 1.92 2.58 2.05 ;
 RECT 2.95 2.485 3.08 2.615 ;
 RECT 2.935 3.785 3.065 3.915 ;
 RECT 1.32 3.51 1.45 3.64 ;
 RECT 2.46 4.095 2.59 4.225 ;
 RECT 3.255 1.76 3.385 1.89 ;
 RECT 2.09 1.585 2.22 1.715 ;
 RECT 0.99 3.915 1.12 4.045 ;
 RECT 1.29 1.59 1.42 1.72 ;
 RECT 1.43 3.92 1.56 4.05 ;
 RECT 0.845 3.515 0.975 3.645 ;
 RECT 2.935 4.095 3.065 4.225 ;
 RECT 3.935 2.36 4.065 2.49 ;
 RECT 1.965 2.485 2.095 2.615 ;
 RECT 3.925 0.625 4.055 0.755 ;
 RECT 3.925 0.35 4.055 0.48 ;
 RECT 3.435 1.155 3.565 1.285 ;
 RECT 3.435 0.895 3.565 1.025 ;
 RECT 3.435 0.625 3.565 0.755 ;
 RECT 3.435 0.35 3.565 0.48 ;
 RECT 2.955 0.625 3.085 0.755 ;
 RECT 2.955 0.35 3.085 0.48 ;
 RECT 2.45 1.155 2.58 1.285 ;
 RECT 2.45 0.895 2.58 1.025 ;
 RECT 2.45 0.625 2.58 0.755 ;
 RECT 2.45 0.35 2.58 0.48 ;
 RECT 1.97 1.155 2.1 1.285 ;
 RECT 1.97 0.895 2.1 1.025 ;
 RECT 1.435 2.315 1.565 2.445 ;
 RECT 0.96 2.315 1.09 2.445 ;
 RECT 1.44 0.52 1.57 0.65 ;
 RECT 1.44 0.83 1.57 0.96 ;
 RECT 0.96 0.52 1.09 0.65 ;
 RECT 0.96 0.83 1.09 0.96 ;
 RECT 0.42 1.09 0.55 1.22 ;
 RECT 3.35 3.855 3.48 3.985 ;
 RECT 0.515 2.795 0.645 2.925 ;
 RECT 3.35 4.115 3.48 4.245 ;
 RECT 0.42 0.83 0.55 0.96 ;
 RECT 1.97 0.35 2.1 0.48 ;
 RECT 1.97 0.625 2.1 0.755 ;
 RECT 2.46 3.785 2.59 3.915 ;
 LAYER M1 ;
 RECT 1.895 2.48 4.135 2.495 ;
 RECT 1.895 2.495 3.225 2.62 ;
 RECT 3.085 2.355 4.135 2.48 ;
 RECT 2.45 4.19 2.595 4.27 ;
 RECT 2.455 3.725 2.595 4.19 ;
 RECT 1.315 4.09 1.455 4.27 ;
 RECT 1.315 4.27 2.595 4.41 ;
 RECT 1.315 3.44 1.455 3.88 ;
 RECT 1.315 3.88 1.61 4.09 ;
 RECT 1.93 1.755 2.235 1.825 ;
 RECT 1.93 1.545 2.27 1.755 ;
 RECT 2.805 2.15 2.945 2.2 ;
 RECT 1.935 2.2 2.945 2.34 ;
 RECT 1.935 2.105 2.075 2.2 ;
 RECT 0.955 1.965 2.075 2.105 ;
 RECT 0.955 0.44 1.095 1.965 ;
 RECT 0.955 2.105 1.095 2.515 ;
 RECT 3.205 1.72 3.435 2.01 ;
 RECT 2.805 2.01 3.435 2.15 ;
 END
END LSDNENX2

MACRO LSDNENX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.68 BY 5.76 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.9 1.42 2.275 1.76 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END ENB

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.615 1.03 6.71 1.17 ;
 RECT 3.55 1.96 3.82 2.1 ;
 RECT 4.535 1.96 4.805 2.1 ;
 RECT 3.615 1.48 4.055 1.785 ;
 RECT 3.615 0.4 3.755 1.03 ;
 RECT 6.57 0.335 6.71 1.03 ;
 RECT 4.6 0.37 4.74 1.03 ;
 RECT 5.595 0.305 5.735 1.03 ;
 RECT 3.615 1.17 3.755 1.48 ;
 RECT 3.615 1.785 3.755 1.96 ;
 RECT 4.6 1.17 4.74 1.96 ;
 END
 ANTENNADIFFAREA 1.998 ;
 END Q

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 7.68 5.2 ;
 RECT 3.56 3.605 3.7 5.04 ;
 RECT 3.975 3.69 4.115 5.04 ;
 END
 END VDDH

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.805 3.855 1.17 4.21 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.68 0.08 ;
 RECT 4.12 0.08 4.26 0.88 ;
 RECT 7.06 0.08 7.2 0.885 ;
 RECT 2.095 0.08 2.235 1.02 ;
 RECT 3.135 0.08 3.275 1.405 ;
 RECT 6.085 0.08 6.225 0.885 ;
 RECT 5.095 0.08 5.235 0.88 ;
 RECT 1.165 0.08 1.305 1.35 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 7.68 5.84 ;
 END
 END VDDL

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.68 2.96 ;
 RECT 6.515 2.57 6.79 2.8 ;
 RECT 5.54 2.585 5.815 2.8 ;
 RECT 0.84 2.96 0.98 3.715 ;
 RECT 2.09 2.245 2.23 2.8 ;
 RECT 0.51 2.96 0.65 2.985 ;
 RECT 0.51 2.735 0.65 2.8 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 2.66 1.7 2.76 3.915 ;
 RECT 1.38 3.88 1.61 3.915 ;
 RECT 1.38 4.015 1.61 4.09 ;
 RECT 3.39 0.19 3.49 1.6 ;
 RECT 2.66 1.6 3.49 1.7 ;
 RECT 3.39 1.7 3.49 2.72 ;
 RECT 4.87 0.19 4.97 2.715 ;
 RECT 4.385 0.19 4.485 2.715 ;
 RECT 3.885 0.19 3.985 2.715 ;
 RECT 1.38 3.915 2.76 4.015 ;
 RECT 3.39 0.09 4.97 0.19 ;
 RECT 5.37 0.09 5.47 1.71 ;
 RECT 5.37 1.71 5.665 1.87 ;
 RECT 6.845 0.09 6.945 1.87 ;
 RECT 6.845 1.97 6.945 2.73 ;
 RECT 6.35 0.09 6.45 1.87 ;
 RECT 6.35 1.97 6.45 2.73 ;
 RECT 5.37 1.97 5.47 2.73 ;
 RECT 5.865 0.09 5.965 1.87 ;
 RECT 5.865 1.97 5.965 2.73 ;
 RECT 5.37 1.87 6.945 1.97 ;
 RECT 1.87 0.205 1.97 1.55 ;
 RECT 1.87 1.55 2.13 1.76 ;
 RECT 1.87 1.76 1.97 2.695 ;
 RECT 1.095 4.085 1.195 4.27 ;
 RECT 3.345 3.46 3.445 4.27 ;
 RECT 1.095 3.265 1.195 3.875 ;
 RECT 0.94 3.875 1.195 4.085 ;
 RECT 1.095 4.27 3.445 4.37 ;
 LAYER CO ;
 RECT 1.43 3.92 1.56 4.05 ;
 RECT 5.485 1.75 5.615 1.88 ;
 RECT 7.065 0.675 7.195 0.805 ;
 RECT 6.575 0.705 6.705 0.835 ;
 RECT 6.575 0.435 6.705 0.565 ;
 RECT 6.575 0.965 6.705 1.095 ;
 RECT 5.1 0.675 5.23 0.805 ;
 RECT 4.605 0.495 4.735 0.625 ;
 RECT 4.605 0.765 4.735 0.895 ;
 RECT 4.605 1.025 4.735 1.155 ;
 RECT 3.98 3.75 4.11 3.88 ;
 RECT 3.09 3.99 3.22 4.12 ;
 RECT 1.17 0.835 1.3 0.965 ;
 RECT 5.61 2.625 5.74 2.755 ;
 RECT 1.32 3.51 1.45 3.64 ;
 RECT 3.565 3.68 3.695 3.81 ;
 RECT 3.62 1.965 3.75 2.095 ;
 RECT 2.1 0.83 2.23 0.96 ;
 RECT 3.14 0.45 3.27 0.58 ;
 RECT 3.565 3.99 3.695 4.12 ;
 RECT 3.62 0.755 3.75 0.885 ;
 RECT 0.845 3.515 0.975 3.645 ;
 RECT 4.12 2.525 4.25 2.655 ;
 RECT 4.125 0.675 4.255 0.805 ;
 RECT 5.6 0.68 5.73 0.81 ;
 RECT 3.14 0.72 3.27 0.85 ;
 RECT 1.17 1.095 1.3 1.225 ;
 RECT 3.98 4.01 4.11 4.14 ;
 RECT 1.62 0.52 1.75 0.65 ;
 RECT 2.095 2.32 2.225 2.45 ;
 RECT 3.62 1.015 3.75 1.145 ;
 RECT 0.515 2.795 0.645 2.925 ;
 RECT 3.14 0.98 3.27 1.11 ;
 RECT 3.62 0.485 3.75 0.615 ;
 RECT 2.1 0.52 2.23 0.65 ;
 RECT 1.62 2.315 1.75 2.445 ;
 RECT 5.6 0.41 5.73 0.54 ;
 RECT 5.6 0.94 5.73 1.07 ;
 RECT 3.135 2.525 3.265 2.655 ;
 RECT 1.62 0.83 1.75 0.96 ;
 RECT 6.09 0.675 6.22 0.805 ;
 RECT 0.99 3.915 1.12 4.045 ;
 RECT 1.95 1.59 2.08 1.72 ;
 RECT 6.585 2.625 6.715 2.755 ;
 RECT 7.095 2.195 7.225 2.325 ;
 RECT 6.1 2.195 6.23 2.325 ;
 RECT 5.1 2.525 5.23 2.655 ;
 RECT 4.605 1.965 4.735 2.095 ;
 LAYER M1 ;
 RECT 3.065 2.52 5.4 2.66 ;
 RECT 5.26 2.33 5.4 2.52 ;
 RECT 5.26 2.19 7.295 2.33 ;
 RECT 1.315 4.09 1.455 4.215 ;
 RECT 3.085 3.405 3.225 4.23 ;
 RECT 1.31 4.215 1.455 4.23 ;
 RECT 1.315 3.44 1.455 3.88 ;
 RECT 1.315 3.88 1.61 4.09 ;
 RECT 1.31 4.23 3.225 4.37 ;
 RECT 3.105 2.05 3.245 2.24 ;
 RECT 1.615 1.91 3.245 2.05 ;
 RECT 1.615 0.44 1.755 1.91 ;
 RECT 1.615 2.05 1.755 2.515 ;
 RECT 4.975 1.885 5.115 2.24 ;
 RECT 3.105 2.24 5.115 2.38 ;
 RECT 4.975 1.745 5.665 1.885 ;
 RECT 5.435 1.71 5.665 1.745 ;
 RECT 5.435 1.885 5.665 1.92 ;
 END
END LSDNENX4

MACRO LSDNENX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.52 BY 5.76 ;
 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 11.52 5.2 ;
 RECT 3 4.005 3.14 5.04 ;
 RECT 3.41 4.025 3.55 5.04 ;
 END
 END VDDH

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.52 0.08 ;
 RECT 3.31 0.08 3.45 0.875 ;
 RECT 8.01 0.08 8.15 0.875 ;
 RECT 4.25 0.08 4.39 0.875 ;
 RECT 5.19 0.08 5.33 0.875 ;
 RECT 10.95 0.08 11.09 1.35 ;
 RECT 10.12 0.08 10.26 1.055 ;
 RECT 6.13 0.08 6.27 0.875 ;
 RECT 2.37 0.08 2.51 0.875 ;
 RECT 7.07 0.08 7.21 0.875 ;
 RECT 8.95 0.08 9.09 0.875 ;
 RECT 1.43 0.08 1.57 0.875 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 11.52 5.84 ;
 END
 END VDDL

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.52 2.96 ;
 RECT 0.965 2.96 1.105 3.785 ;
 RECT 10.845 2.38 10.985 2.8 ;
 RECT 10.12 1.81 10.26 2.8 ;
 RECT 5.66 1.94 5.8 2.8 ;
 RECT 0.35 2.96 0.49 3.765 ;
 RECT 6.6 1.915 6.74 2.8 ;
 RECT 7.54 1.915 7.68 2.8 ;
 RECT 8.48 1.915 8.62 2.8 ;
 END
 END VSS

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.93 1.25 10.3 1.49 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END ENB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.84 3.935 1.295 4.28 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.725 1.48 2.04 1.825 ;
 RECT 1.9 1.825 2.04 2.215 ;
 RECT 1.9 1.02 8.62 1.16 ;
 RECT 1.9 1.16 2.04 1.48 ;
 RECT 1.9 0.345 2.04 1.02 ;
 RECT 6.6 0.345 6.74 1.02 ;
 RECT 4.72 1.16 4.86 2.215 ;
 RECT 2.84 0.345 2.98 1.02 ;
 RECT 7.54 0.345 7.68 1.02 ;
 RECT 3.78 0.345 3.92 1.02 ;
 RECT 8.48 0.345 8.62 1.02 ;
 RECT 4.72 0.345 4.86 1.02 ;
 RECT 2.84 1.16 2.98 2.215 ;
 RECT 5.66 0.345 5.8 1.02 ;
 RECT 3.78 1.16 3.92 2.215 ;
 END
 ANTENNADIFFAREA 3.96 ;
 END Q

 OBS
 LAYER PO ;
 RECT 6.855 0.175 6.955 2.495 ;
 RECT 8.265 0.175 8.365 2.495 ;
 RECT 6.385 0.175 6.485 2.495 ;
 RECT 7.795 0.175 7.895 2.495 ;
 RECT 5.915 0.175 6.015 2.495 ;
 RECT 7.325 0.175 7.425 2.495 ;
 RECT 5.445 0.175 5.545 2.495 ;
 RECT 8.735 0.175 8.835 2.495 ;
 RECT 9.25 2.37 9.48 2.495 ;
 RECT 5.445 2.495 9.48 2.595 ;
 RECT 1.22 4.145 1.32 4.63 ;
 RECT 2.785 3.805 2.885 4.63 ;
 RECT 1.22 3.345 1.32 3.935 ;
 RECT 1.065 3.935 1.32 4.145 ;
 RECT 1.22 4.63 2.885 4.73 ;
 RECT 9.905 0.325 10.005 1.27 ;
 RECT 9.905 1.27 10.16 1.48 ;
 RECT 9.905 1.48 10.005 2.435 ;
 RECT 1.835 2.635 1.935 3.155 ;
 RECT 4.505 0.175 4.605 2.535 ;
 RECT 2.155 0.175 2.255 2.535 ;
 RECT 4.035 0.175 4.135 2.535 ;
 RECT 1.685 0.175 1.785 2.535 ;
 RECT 3.565 0.175 3.665 2.535 ;
 RECT 3.095 0.175 3.195 2.535 ;
 RECT 4.975 0.175 5.075 2.535 ;
 RECT 2.625 0.175 2.725 2.535 ;
 RECT 1.685 2.535 5.075 2.635 ;
 RECT 1.78 3.155 2.01 3.365 ;
 LAYER CO ;
 RECT 10.955 1.15 11.085 1.28 ;
 RECT 10.85 2.73 10.98 2.86 ;
 RECT 10.85 2.47 10.98 2.6 ;
 RECT 3.415 4.355 3.545 4.485 ;
 RECT 3.415 4.095 3.545 4.225 ;
 RECT 10.955 0.89 11.085 1.02 ;
 RECT 8.955 0.415 9.085 0.545 ;
 RECT 8.955 0.675 9.085 0.805 ;
 RECT 8.955 2.015 9.085 2.145 ;
 RECT 8.485 0.675 8.615 0.805 ;
 RECT 1.905 0.675 2.035 0.805 ;
 RECT 1.905 0.415 2.035 0.545 ;
 RECT 1.435 2.015 1.565 2.145 ;
 RECT 1.435 0.415 1.565 0.545 ;
 RECT 1.435 0.675 1.565 0.805 ;
 RECT 2.535 4.355 2.665 4.485 ;
 RECT 0.97 3.585 1.1 3.715 ;
 RECT 1.44 3.595 1.57 3.725 ;
 RECT 3.005 4.315 3.135 4.445 ;
 RECT 3.005 4.055 3.135 4.185 ;
 RECT 9.655 2.015 9.785 2.145 ;
 RECT 9.655 0.595 9.785 0.725 ;
 RECT 9.655 0.855 9.785 0.985 ;
 RECT 10.125 0.595 10.255 0.725 ;
 RECT 10.125 2.015 10.255 2.145 ;
 RECT 10.125 0.855 10.255 0.985 ;
 RECT 0.355 3.48 0.485 3.61 ;
 RECT 0.355 3.22 0.485 3.35 ;
 RECT 9.3 2.41 9.43 2.54 ;
 RECT 1.115 3.975 1.245 4.105 ;
 RECT 9.98 1.31 10.11 1.44 ;
 RECT 1.83 3.195 1.96 3.325 ;
 RECT 7.075 0.415 7.205 0.545 ;
 RECT 8.485 0.415 8.615 0.545 ;
 RECT 8.015 0.415 8.145 0.545 ;
 RECT 7.545 0.675 7.675 0.805 ;
 RECT 7.545 2.015 7.675 2.145 ;
 RECT 8.015 2.015 8.145 2.145 ;
 RECT 7.545 0.415 7.675 0.545 ;
 RECT 7.075 2.015 7.205 2.145 ;
 RECT 8.015 0.675 8.145 0.805 ;
 RECT 8.485 2.015 8.615 2.145 ;
 RECT 7.075 0.675 7.205 0.805 ;
 RECT 6.605 0.415 6.735 0.545 ;
 RECT 5.665 0.675 5.795 0.805 ;
 RECT 6.135 2.015 6.265 2.145 ;
 RECT 6.135 0.675 6.265 0.805 ;
 RECT 6.605 0.675 6.735 0.805 ;
 RECT 6.135 0.415 6.265 0.545 ;
 RECT 5.665 2.015 5.795 2.145 ;
 RECT 5.665 0.415 5.795 0.545 ;
 RECT 6.605 2.015 6.735 2.145 ;
 RECT 5.195 0.415 5.325 0.545 ;
 RECT 4.255 0.675 4.385 0.805 ;
 RECT 4.725 2.015 4.855 2.145 ;
 RECT 4.725 0.675 4.855 0.805 ;
 RECT 5.195 0.675 5.325 0.805 ;
 RECT 4.725 0.415 4.855 0.545 ;
 RECT 4.255 2.015 4.385 2.145 ;
 RECT 4.255 0.415 4.385 0.545 ;
 RECT 5.195 2.015 5.325 2.145 ;
 RECT 3.785 0.415 3.915 0.545 ;
 RECT 2.845 0.675 2.975 0.805 ;
 RECT 3.315 2.015 3.445 2.145 ;
 RECT 3.315 0.675 3.445 0.805 ;
 RECT 3.785 0.675 3.915 0.805 ;
 RECT 3.315 0.415 3.445 0.545 ;
 RECT 2.845 2.015 2.975 2.145 ;
 RECT 2.845 0.415 2.975 0.545 ;
 RECT 3.785 2.015 3.915 2.145 ;
 RECT 2.375 2.015 2.505 2.145 ;
 RECT 1.905 2.015 2.035 2.145 ;
 RECT 2.375 0.675 2.505 0.805 ;
 RECT 2.535 4.095 2.665 4.225 ;
 RECT 2.375 0.415 2.505 0.545 ;
 LAYER M1 ;
 RECT 8.01 1.775 8.15 2.215 ;
 RECT 7.07 1.775 7.21 2.215 ;
 RECT 6.13 1.775 6.27 2.215 ;
 RECT 4.25 1.945 4.39 2.48 ;
 RECT 3.31 1.945 3.45 2.48 ;
 RECT 2.37 1.945 2.51 2.48 ;
 RECT 1.43 1.945 1.57 2.48 ;
 RECT 1.43 2.48 5.33 2.62 ;
 RECT 5.19 1.775 5.33 2.48 ;
 RECT 8.95 1.775 9.09 2.215 ;
 RECT 5.19 1.635 9.09 1.775 ;
 RECT 9.65 0.525 9.79 2.415 ;
 RECT 9.25 2.37 9.48 2.415 ;
 RECT 9.25 2.555 9.48 2.58 ;
 RECT 9.25 2.415 9.79 2.555 ;
 RECT 1.435 3.365 1.575 4.215 ;
 RECT 2.53 4.045 2.67 4.215 ;
 RECT 2.53 4.355 2.67 4.535 ;
 RECT 1.78 3.155 2.01 3.225 ;
 RECT 1.435 3.225 2.01 3.365 ;
 RECT 1.435 4.215 2.67 4.355 ;
 END
END LSDNENX8

MACRO LSDNX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.08 BY 5.76 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.3 1.795 5.6 2.03 ;
 RECT 5.3 1.47 5.6 1.655 ;
 RECT 4.675 1.655 5.6 1.795 ;
 RECT 4.675 0.53 4.815 1.655 ;
 END
 ANTENNADIFFAREA 0.63 ;
 END Q

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 6.08 5.2 ;
 RECT 1.46 3.965 1.6 5.04 ;
 RECT 1.97 4.015 2.11 5.04 ;
 END
 END VDDH

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.995 4.04 4.295 4.31 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.08 2.96 ;
 RECT 4.185 2.96 4.325 3.75 ;
 RECT 3.205 2.96 3.345 3.745 ;
 RECT 5.145 2.96 5.285 3.725 ;
 END
 END VSS

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.08 0.08 ;
 RECT 4.185 0.08 4.325 1.175 ;
 RECT 3.67 0.08 3.81 1.34 ;
 RECT 5.145 0.08 5.285 1 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 6.08 5.84 ;
 END
 END VDDL

 OBS
 LAYER PO ;
 RECT 3.97 4.29 4.07 4.63 ;
 RECT 2.225 3.815 2.325 4.63 ;
 RECT 3.97 3.365 4.07 4.06 ;
 RECT 3.97 4.06 4.27 4.29 ;
 RECT 2.225 4.63 4.07 4.73 ;
 RECT 4.93 0.145 5.03 2.99 ;
 RECT 4.45 0.17 4.55 2.99 ;
 RECT 4.45 3.09 4.55 3.935 ;
 RECT 3.56 3.09 3.785 3.335 ;
 RECT 4.93 3.09 5.03 3.935 ;
 RECT 3.56 2.99 5.03 3.09 ;
 RECT 5.455 2.03 5.555 3.51 ;
 RECT 5.455 3.51 5.685 3.74 ;
 RECT 5.325 1.79 5.555 2.03 ;
 LAYER CO ;
 RECT 4.095 4.11 4.225 4.24 ;
 RECT 4.19 3.525 4.32 3.655 ;
 RECT 2.445 4.27 2.575 4.4 ;
 RECT 4.68 1.195 4.81 1.325 ;
 RECT 1.465 4.055 1.595 4.185 ;
 RECT 4.68 3.525 4.81 3.655 ;
 RECT 3.675 0.88 3.805 1.01 ;
 RECT 5.505 3.56 5.635 3.69 ;
 RECT 4.19 0.435 4.32 0.565 ;
 RECT 3.72 3.585 3.85 3.715 ;
 RECT 3.675 0.62 3.805 0.75 ;
 RECT 1.975 4.165 2.105 4.295 ;
 RECT 3.21 3.285 3.34 3.415 ;
 RECT 4.68 3.265 4.81 3.395 ;
 RECT 4.19 3.525 4.32 3.655 ;
 RECT 4.19 0.975 4.32 1.105 ;
 RECT 1.465 4.315 1.595 4.445 ;
 RECT 4.19 0.715 4.32 0.845 ;
 RECT 3.61 3.155 3.74 3.285 ;
 RECT 5.15 3.265 5.28 3.395 ;
 RECT 5.15 3.525 5.28 3.655 ;
 RECT 5.15 0.715 5.28 0.845 ;
 RECT 5.15 0.435 5.28 0.565 ;
 RECT 4.68 0.935 4.81 1.065 ;
 RECT 4.68 0.655 4.81 0.785 ;
 RECT 3.675 1.14 3.805 1.27 ;
 RECT 5.375 1.85 5.505 1.98 ;
 RECT 3.21 3.545 3.34 3.675 ;
 LAYER M1 ;
 RECT 4.675 3.165 4.815 3.865 ;
 RECT 4.675 3.865 5.685 4.005 ;
 RECT 5.455 3.51 5.685 3.865 ;
 RECT 2.44 4.15 2.58 4.265 ;
 RECT 2.44 4.405 2.58 4.515 ;
 RECT 3.715 3.355 3.855 4.265 ;
 RECT 3.555 3.105 3.855 3.355 ;
 RECT 2.44 4.265 3.855 4.405 ;
 END
END LSDNX2

MACRO LSDNX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.04 BY 5.76 ;
 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 7.04 5.2 ;
 RECT 1.465 3.975 1.605 5.04 ;
 RECT 1.975 3.985 2.115 5.04 ;
 END
 END VDDH

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.04 2.96 ;
 RECT 4.185 2.96 4.325 3.79 ;
 RECT 5.14 2.96 5.28 3.72 ;
 RECT 6.09 2.96 6.23 3.74 ;
 RECT 3.205 2.96 3.345 3.74 ;
 END
 END VSS

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.04 0.08 ;
 RECT 6.09 0.08 6.23 1.91 ;
 RECT 4.195 0.08 4.335 2.225 ;
 RECT 5.14 0.08 5.28 2.125 ;
 RECT 3.67 0.08 3.81 1.975 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 7.04 5.84 ;
 END
 END VDDL

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.995 3.935 4.295 4.205 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.37 2.56 6.67 2.565 ;
 RECT 6.265 2.105 6.665 2.295 ;
 RECT 5.62 1.72 5.76 2.295 ;
 RECT 4.67 1.7 4.81 2.295 ;
 RECT 4.67 2.295 6.67 2.435 ;
 RECT 6.265 2.435 6.67 2.56 ;
 END
 ANTENNADIFFAREA 1.15 ;
 END Q

 OBS
 LAYER PO ;
 RECT 3.97 4.185 4.07 4.6 ;
 RECT 2.23 3.72 2.33 4.6 ;
 RECT 3.97 3.36 4.07 3.955 ;
 RECT 3.97 3.955 4.27 4.185 ;
 RECT 2.23 4.6 4.07 4.7 ;
 RECT 4.45 1.11 4.55 2.545 ;
 RECT 4.45 2.545 5.975 2.645 ;
 RECT 4.45 2.645 4.55 3.08 ;
 RECT 4.45 3.18 4.55 3.93 ;
 RECT 3.56 3.18 3.785 3.375 ;
 RECT 4.925 1.125 5.025 2.545 ;
 RECT 4.925 2.645 5.025 3.93 ;
 RECT 5.875 1.125 5.975 2.545 ;
 RECT 5.875 2.645 5.975 3.93 ;
 RECT 5.395 1.125 5.495 2.545 ;
 RECT 5.395 2.645 5.495 3.93 ;
 RECT 3.56 3.08 4.55 3.18 ;
 RECT 6.42 2.545 6.52 3.115 ;
 RECT 6.42 3.115 6.645 3.345 ;
 RECT 6.42 2.315 6.645 2.545 ;
 LAYER CO ;
 RECT 5.625 1.805 5.755 1.935 ;
 RECT 6.47 3.165 6.6 3.295 ;
 RECT 1.47 4.045 1.6 4.175 ;
 RECT 2.45 4.28 2.58 4.41 ;
 RECT 3.675 1.255 3.805 1.385 ;
 RECT 3.675 1.515 3.805 1.645 ;
 RECT 1.98 4.19 2.11 4.32 ;
 RECT 3.675 1.775 3.805 1.905 ;
 RECT 4.095 4.005 4.225 4.135 ;
 RECT 3.21 3.28 3.34 3.41 ;
 RECT 4.2 1.41 4.33 1.54 ;
 RECT 4.675 2.105 4.805 2.235 ;
 RECT 1.47 4.305 1.6 4.435 ;
 RECT 6.095 1.685 6.225 1.815 ;
 RECT 4.675 1.805 4.805 1.935 ;
 RECT 3.61 3.195 3.74 3.325 ;
 RECT 5.145 3.52 5.275 3.65 ;
 RECT 5.615 3.34 5.745 3.47 ;
 RECT 3.21 3.54 3.34 3.67 ;
 RECT 6.095 3.52 6.225 3.65 ;
 RECT 4.2 1.985 4.33 2.115 ;
 RECT 6.095 1.41 6.225 1.54 ;
 RECT 3.72 3.58 3.85 3.71 ;
 RECT 4.19 3.57 4.32 3.7 ;
 RECT 5.625 2.105 5.755 2.235 ;
 RECT 4.67 3.34 4.8 3.47 ;
 RECT 6.47 2.365 6.6 2.495 ;
 RECT 5.145 1.925 5.275 2.055 ;
 RECT 5.145 1.41 5.275 1.54 ;
 LAYER M1 ;
 RECT 5.61 3.27 5.75 3.945 ;
 RECT 4.665 3.27 4.805 3.945 ;
 RECT 6.37 3.365 6.51 3.945 ;
 RECT 4.66 3.945 6.51 4.085 ;
 RECT 6.37 3.1 6.67 3.365 ;
 RECT 2.445 4.08 2.585 4.275 ;
 RECT 2.445 4.415 2.585 4.47 ;
 RECT 3.715 3.395 3.855 4.275 ;
 RECT 3.555 3.145 3.855 3.395 ;
 RECT 2.445 4.275 3.855 4.415 ;
 END
END LSDNX4

MACRO LSDNX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.24 BY 5.76 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.215 1.475 9.62 1.795 ;
 RECT 8.54 0.81 8.68 1.795 ;
 RECT 7.585 0.81 7.725 1.795 ;
 RECT 6.615 0.81 6.755 1.795 ;
 RECT 5.65 0.81 5.79 1.795 ;
 RECT 5.65 1.795 9.62 1.935 ;
 END
 ANTENNADIFFAREA 2.28 ;
 END Q

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.24 0.08 ;
 RECT 4.01 0.08 4.15 1.215 ;
 RECT 5.17 0.08 5.31 1.255 ;
 RECT 9.01 0.08 9.15 1.24 ;
 RECT 8.055 0.08 8.195 1.435 ;
 RECT 7.085 0.08 7.225 1.435 ;
 RECT 6.12 0.08 6.26 1.435 ;
 RECT 2.145 0.08 2.285 1.35 ;
 RECT 2.67 0.08 2.81 1.535 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 10.24 5.84 ;
 END
 END VDDL

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.28 2.8 10.24 2.96 ;
 RECT 4.005 2.96 4.145 3.82 ;
 RECT 9.01 2.96 9.15 3.95 ;
 RECT 8.055 2.96 8.195 3.95 ;
 RECT 7.085 2.96 7.225 3.945 ;
 RECT 2.67 2.96 2.81 3.71 ;
 RECT 1.585 2.96 1.725 3.4 ;
 RECT 5.13 3.555 5.27 3.935 ;
 RECT 6.12 3.555 6.26 3.95 ;
 RECT 5.13 3.415 6.26 3.555 ;
 RECT 6.12 2.96 6.26 3.415 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.47 3.87 2.77 4.14 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END D

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 10.24 5.2 ;
 RECT 2.66 4.28 2.8 5.04 ;
 RECT 1.44 3.96 1.58 5.04 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 2.445 3.89 2.745 4.12 ;
 RECT 2.445 4.12 2.545 4.69 ;
 RECT 2.445 3.24 2.545 3.89 ;
 RECT 3.785 1.995 3.885 3.11 ;
 RECT 3.205 3.11 3.885 3.21 ;
 RECT 3.785 3.21 3.885 4.125 ;
 RECT 4.265 0.41 4.365 1.895 ;
 RECT 4.265 1.995 4.365 4.125 ;
 RECT 4.895 0.405 4.995 1.895 ;
 RECT 4.895 1.995 4.995 4.135 ;
 RECT 3.205 1.895 4.995 1.995 ;
 RECT 3.205 1.765 3.43 1.895 ;
 RECT 3.785 0.405 3.885 1.895 ;
 RECT 3.205 3.21 3.43 3.34 ;
 RECT 9.37 1.915 9.47 3.115 ;
 RECT 9.37 3.115 9.595 3.345 ;
 RECT 9.37 1.685 9.595 1.915 ;
 RECT 2.09 2.74 2.19 3.02 ;
 RECT 2.925 0.405 3.025 2.64 ;
 RECT 2.925 2.74 3.025 4 ;
 RECT 2.09 2.64 3.025 2.74 ;
 RECT 2.035 3.02 2.26 3.33 ;
 RECT 8.325 0.41 8.425 4.035 ;
 RECT 5.435 1.99 5.535 3.05 ;
 RECT 5.435 3.28 5.535 4.035 ;
 RECT 5.435 0.41 5.535 1.76 ;
 RECT 5.235 1.76 5.535 1.99 ;
 RECT 5.905 0.41 6.005 4.035 ;
 RECT 6.4 0.41 6.5 4.035 ;
 RECT 6.87 0.41 6.97 4.035 ;
 RECT 7.37 0.41 7.47 4.035 ;
 RECT 7.84 0.41 7.94 4.035 ;
 RECT 7.84 0.31 8.425 0.41 ;
 RECT 8.795 0.41 8.895 4.035 ;
 RECT 5.305 3.05 5.535 3.28 ;
 RECT 5.435 4.035 6.005 4.135 ;
 RECT 5.905 0.31 6.5 0.41 ;
 RECT 6.4 4.035 6.97 4.135 ;
 RECT 6.87 0.31 7.47 0.41 ;
 RECT 7.37 4.035 7.94 4.135 ;
 RECT 8.325 4.035 8.895 4.135 ;
 LAYER CO ;
 RECT 3.15 0.89 3.28 1.02 ;
 RECT 4.015 0.72 4.145 0.85 ;
 RECT 9.015 3.715 9.145 3.845 ;
 RECT 4.6 3.635 4.73 3.765 ;
 RECT 3.53 1.235 3.66 1.365 ;
 RECT 2.085 3.15 2.215 3.28 ;
 RECT 5.355 3.11 5.485 3.24 ;
 RECT 2.195 3.46 2.325 3.59 ;
 RECT 7.59 3.635 7.72 3.765 ;
 RECT 7.09 0.72 7.22 0.85 ;
 RECT 2.57 3.94 2.7 4.07 ;
 RECT 5.655 0.895 5.785 1.025 ;
 RECT 2.15 0.63 2.28 0.76 ;
 RECT 2.195 4.34 2.325 4.47 ;
 RECT 8.545 0.895 8.675 1.025 ;
 RECT 9.42 1.735 9.55 1.865 ;
 RECT 1.59 3.2 1.72 3.33 ;
 RECT 4.01 3.585 4.14 3.715 ;
 RECT 9.42 3.165 9.55 3.295 ;
 RECT 6.125 3.715 6.255 3.845 ;
 RECT 2.15 0.89 2.28 1.02 ;
 RECT 2.665 4.34 2.795 4.47 ;
 RECT 2.15 1.15 2.28 1.28 ;
 RECT 5.175 1 5.305 1.13 ;
 RECT 3.255 1.815 3.385 1.945 ;
 RECT 1.59 2.935 1.72 3.065 ;
 RECT 8.06 3.715 8.19 3.845 ;
 RECT 3.255 3.16 3.385 3.29 ;
 RECT 7.59 0.895 7.72 1.025 ;
 RECT 9.015 0.985 9.145 1.115 ;
 RECT 2.675 1.22 2.805 1.35 ;
 RECT 9.015 0.72 9.145 0.85 ;
 RECT 3.15 3.53 3.28 3.66 ;
 RECT 5.175 0.72 5.305 0.85 ;
 RECT 6.62 0.895 6.75 1.025 ;
 RECT 3.15 1.34 3.28 1.47 ;
 RECT 1.445 4.29 1.575 4.42 ;
 RECT 1.445 4.03 1.575 4.16 ;
 RECT 4.6 1.28 4.73 1.41 ;
 RECT 8.545 1.28 8.675 1.41 ;
 RECT 5.655 3.765 5.785 3.895 ;
 RECT 3.53 0.72 3.66 0.85 ;
 RECT 2.675 3.465 2.805 3.595 ;
 RECT 8.06 1.235 8.19 1.365 ;
 RECT 5.655 1.28 5.785 1.41 ;
 RECT 6.125 1.235 6.255 1.365 ;
 RECT 8.545 3.635 8.675 3.765 ;
 RECT 6.62 1.28 6.75 1.41 ;
 RECT 6.62 3.635 6.75 3.765 ;
 RECT 5.135 3.715 5.265 3.845 ;
 RECT 5.285 1.81 5.415 1.94 ;
 RECT 7.09 3.715 7.22 3.845 ;
 RECT 7.59 1.28 7.72 1.41 ;
 RECT 7.09 1.235 7.22 1.365 ;
 RECT 4.6 0.895 4.73 1.025 ;
 RECT 8.06 0.72 8.19 0.85 ;
 RECT 2.675 0.645 2.805 0.775 ;
 RECT 6.125 0.72 6.255 0.85 ;
 RECT 4.015 0.98 4.145 1.11 ;
 RECT 3.525 3.715 3.655 3.845 ;
 LAYER M1 ;
 RECT 3.525 1.465 5.155 1.605 ;
 RECT 4.595 0.81 4.735 1.465 ;
 RECT 5.015 1.605 5.155 1.805 ;
 RECT 3.525 0.65 3.665 1.465 ;
 RECT 5.015 1.805 5.49 1.945 ;
 RECT 8.54 3.565 8.68 4.16 ;
 RECT 7.585 3.565 7.725 4.16 ;
 RECT 6.615 3.565 6.755 4.16 ;
 RECT 5.65 3.695 5.79 4.16 ;
 RECT 5.65 4.16 9.46 4.3 ;
 RECT 9.32 3.365 9.46 4.16 ;
 RECT 9.32 3.105 9.62 3.365 ;
 RECT 2.19 3.35 2.33 4.53 ;
 RECT 2.03 3.1 2.33 3.35 ;
 RECT 3.145 3.14 3.455 3.36 ;
 RECT 3.155 3.1 3.455 3.14 ;
 RECT 3.145 3.36 3.285 3.875 ;
 RECT 3.145 1.745 3.455 2.01 ;
 RECT 3.155 2.01 3.455 2.015 ;
 RECT 3.145 0.785 3.285 1.745 ;
 RECT 4.595 3.255 4.735 4.095 ;
 RECT 3.52 4.095 4.735 4.235 ;
 RECT 3.52 3.615 3.66 4.095 ;
 RECT 5.305 3.1 5.535 3.115 ;
 RECT 5.305 3.255 5.535 3.27 ;
 RECT 4.595 3.115 5.535 3.255 ;
 END
END LSDNX8

MACRO LSUPENCLX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 5.76 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 1.685 3.395 1.945 3.535 ;
 RECT 1.325 2.085 1.6 2.225 ;
 RECT 2.46 2.96 2.88 3.645 ;
 RECT 2.285 2.02 2.425 2.8 ;
 RECT 3.185 2.1 3.325 2.8 ;
 RECT 3.185 2.96 3.325 3.475 ;
 RECT 1.75 3.535 1.89 3.58 ;
 RECT 1.75 2.96 1.89 3.395 ;
 RECT 1.425 2.225 1.565 2.8 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 3.72 1.96 3.745 ;
 RECT 2.05 3.11 2.32 3.25 ;
 RECT 1.555 3.885 1.96 4.04 ;
 RECT 1.555 3.745 2.255 3.885 ;
 RECT 2.115 3.25 2.255 3.745 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 4.8 5.2 ;
 RECT 2.07 4.26 2.49 4.665 ;
 RECT 2.215 4.665 2.355 5.04 ;
 RECT 1.745 4.3 1.885 5.04 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.6 1.475 2.905 1.81 ;
 RECT 2.765 0.545 2.905 1.475 ;
 RECT 3.655 2.4 4.14 2.62 ;
 RECT 2.765 1.82 3.795 1.96 ;
 RECT 2.765 1.96 2.905 2.29 ;
 RECT 2.765 1.81 2.905 1.82 ;
 RECT 3.655 1.96 3.795 2.4 ;
 END
 ANTENNADIFFAREA 0.73 ;
 END Q

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.4 1.38 3.73 1.68 ;
 END
 ANTENNAGATEAREA 0.16 ;
 END ENB

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 0.47 0.08 0.61 1.275 ;
 RECT 3.655 0.08 3.795 1.02 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 4.8 5.84 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 1 2.535 1.1 3.06 ;
 RECT 1.15 1.84 1.25 2.435 ;
 RECT 1 2.435 1.25 2.535 ;
 RECT 0.93 3.06 1.16 3.29 ;
 RECT 1.53 3.17 1.63 3.785 ;
 RECT 1.53 3.785 1.83 4.015 ;
 RECT 1.53 4.015 1.63 4.73 ;
 RECT 1.15 0.215 1.25 1.29 ;
 RECT 2.55 0.215 2.65 1.595 ;
 RECT 2.2 1.595 2.65 1.825 ;
 RECT 2.55 1.825 2.65 2.685 ;
 RECT 1.15 0.115 2.65 0.215 ;
 RECT 1.65 2.4 2.145 2.5 ;
 RECT 2.045 2.5 2.145 3.065 ;
 RECT 2.045 3.065 2.3 3.295 ;
 RECT 1.65 1.84 1.75 2.4 ;
 RECT 1.455 1.165 1.75 1.395 ;
 RECT 1.65 0.395 1.75 1.165 ;
 RECT 3.975 2.615 4.075 3.155 ;
 RECT 3.91 3.155 4.14 3.385 ;
 RECT 3.91 2.405 4.14 2.615 ;
 RECT 3.44 1.64 3.54 3.795 ;
 RECT 3.44 0.145 3.54 1.43 ;
 RECT 3.44 1.43 3.67 1.64 ;
 LAYER CO ;
 RECT 1.505 1.215 1.635 1.345 ;
 RECT 2.295 1.125 2.425 1.255 ;
 RECT 0.9 0.835 1.03 0.965 ;
 RECT 1.28 3.4 1.41 3.53 ;
 RECT 2.77 2.09 2.9 2.22 ;
 RECT 0.98 3.11 1.11 3.24 ;
 RECT 0.475 0.565 0.605 0.695 ;
 RECT 1.75 4.37 1.88 4.5 ;
 RECT 1.87 0.815 2 0.945 ;
 RECT 2.465 3.185 2.595 3.315 ;
 RECT 0.9 2.09 1.03 2.22 ;
 RECT 2.225 4.3 2.355 4.43 ;
 RECT 2.25 1.645 2.38 1.775 ;
 RECT 2.77 1.19 2.9 1.32 ;
 RECT 2.465 3.445 2.595 3.575 ;
 RECT 1.4 2.09 1.53 2.22 ;
 RECT 2.745 3.445 2.875 3.575 ;
 RECT 1.65 3.835 1.78 3.965 ;
 RECT 2.295 0.815 2.425 0.945 ;
 RECT 2.12 3.115 2.25 3.245 ;
 RECT 2.77 0.93 2.9 1.06 ;
 RECT 2.77 0.665 2.9 0.795 ;
 RECT 3.19 0.56 3.32 0.69 ;
 RECT 0.475 1.085 0.605 1.215 ;
 RECT 3.96 3.205 4.09 3.335 ;
 RECT 3.66 2.09 3.79 2.22 ;
 RECT 3.19 2.16 3.32 2.29 ;
 RECT 3.66 3.295 3.79 3.425 ;
 RECT 3.19 3.295 3.32 3.425 ;
 RECT 3.66 0.82 3.79 0.95 ;
 RECT 3.66 0.51 3.79 0.64 ;
 RECT 3.19 0.82 3.32 0.95 ;
 RECT 3.19 0.82 3.32 0.95 ;
 RECT 1.28 4.36 1.41 4.49 ;
 RECT 0.475 0.825 0.605 0.955 ;
 RECT 1.87 2.09 2 2.22 ;
 RECT 2.29 2.09 2.42 2.22 ;
 RECT 2.745 3.185 2.875 3.315 ;
 RECT 1.4 0.83 1.53 0.96 ;
 RECT 1.755 3.4 1.885 3.53 ;
 RECT 3.96 2.445 4.09 2.575 ;
 RECT 3.49 1.47 3.62 1.6 ;
 LAYER M1 ;
 RECT 1.395 0.38 1.535 1.02 ;
 RECT 2.29 0.38 2.43 1.385 ;
 RECT 3.185 0.38 3.325 1.02 ;
 RECT 1.395 0.24 3.325 0.38 ;
 RECT 0.895 0.76 1.035 1.45 ;
 RECT 0.895 1.59 1.035 2.29 ;
 RECT 1.5 1.165 1.64 1.45 ;
 RECT 0.895 1.45 1.64 1.59 ;
 RECT 1.275 3.245 1.415 4.56 ;
 RECT 0.93 3.105 1.415 3.245 ;
 RECT 3.6 3.1 4.195 3.51 ;
 RECT 1.865 0.745 2.005 1.64 ;
 RECT 1.865 1.78 2.005 2.29 ;
 RECT 1.865 1.64 2.46 1.78 ;
 RECT 2.2 1.6 2.46 1.64 ;
 RECT 2.2 1.78 2.46 1.83 ;
 END
END LSUPENCLX1

MACRO LSUPENCLX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 5.76 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 1.685 3.395 1.945 3.535 ;
 RECT 1.325 2.085 1.6 2.225 ;
 RECT 2.46 2.96 2.88 3.645 ;
 RECT 2.285 2.16 2.425 2.8 ;
 RECT 3.245 2.16 3.385 2.8 ;
 RECT 3.63 2.1 3.77 2.8 ;
 RECT 1.75 3.535 1.89 3.58 ;
 RECT 1.75 2.96 1.89 3.395 ;
 RECT 1.425 2.225 1.565 2.8 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 3.72 1.96 3.745 ;
 RECT 2.05 3.11 2.32 3.25 ;
 RECT 1.555 3.885 1.96 4.04 ;
 RECT 1.555 3.745 2.255 3.885 ;
 RECT 2.115 3.25 2.255 3.745 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END D

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 4.8 5.2 ;
 RECT 2.07 4.26 2.49 4.665 ;
 RECT 2.215 4.665 2.355 5.04 ;
 RECT 1.745 4.3 1.885 5.04 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.6 1.475 2.905 1.81 ;
 RECT 2.765 0.545 2.905 1.475 ;
 RECT 2.765 1.82 4.24 1.96 ;
 RECT 2.765 1.96 2.905 2.415 ;
 RECT 2.765 1.81 2.905 1.82 ;
 RECT 4.1 1.96 4.24 2.315 ;
 END
 ANTENNADIFFAREA 0.62 ;
 END Q

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.865 1.38 4.195 1.68 ;
 END
 ANTENNAGATEAREA 0.14 ;
 END ENB

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 0.47 0.08 0.61 1.275 ;
 RECT 4.1 0.08 4.24 1.02 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 4.8 5.84 ;
 END
 END VDDH

 OBS
 LAYER PO ;
 RECT 1.455 1.365 1.75 1.595 ;
 RECT 1.65 0.395 1.75 1.365 ;
 RECT 1 2.535 1.1 3.06 ;
 RECT 1.15 1.84 1.25 2.435 ;
 RECT 1 2.435 1.25 2.535 ;
 RECT 0.93 3.06 1.16 3.29 ;
 RECT 1.53 3.17 1.63 3.785 ;
 RECT 1.53 3.785 1.83 4.015 ;
 RECT 1.53 4.015 1.63 4.73 ;
 RECT 3.02 0.215 3.12 2.715 ;
 RECT 1.15 0.215 1.25 1.3 ;
 RECT 1.15 0.115 3.12 0.215 ;
 RECT 2.55 0.215 2.65 1.595 ;
 RECT 2.2 1.595 2.65 1.825 ;
 RECT 2.55 1.825 2.65 2.685 ;
 RECT 1.65 2.4 2.145 2.5 ;
 RECT 2.045 2.5 2.145 3.065 ;
 RECT 2.045 3.065 2.3 3.295 ;
 RECT 1.65 1.84 1.75 2.4 ;
 RECT 3.885 1.64 3.985 2.545 ;
 RECT 3.885 0.09 3.985 1.43 ;
 RECT 3.885 1.43 4.115 1.64 ;
 LAYER CO ;
 RECT 1.505 1.415 1.635 1.545 ;
 RECT 2.295 1.125 2.425 1.255 ;
 RECT 0.9 0.835 1.03 0.965 ;
 RECT 1.28 3.4 1.41 3.53 ;
 RECT 2.77 2.21 2.9 2.34 ;
 RECT 0.98 3.11 1.11 3.24 ;
 RECT 0.475 0.565 0.605 0.695 ;
 RECT 1.75 4.37 1.88 4.5 ;
 RECT 1.87 0.815 2 0.945 ;
 RECT 2.465 3.185 2.595 3.315 ;
 RECT 0.9 2.09 1.03 2.22 ;
 RECT 2.225 4.3 2.355 4.43 ;
 RECT 2.25 1.645 2.38 1.775 ;
 RECT 2.77 1.19 2.9 1.32 ;
 RECT 2.465 3.445 2.595 3.575 ;
 RECT 1.4 2.09 1.53 2.22 ;
 RECT 2.745 3.445 2.875 3.575 ;
 RECT 1.65 3.835 1.78 3.965 ;
 RECT 2.295 0.815 2.425 0.945 ;
 RECT 2.12 3.115 2.25 3.245 ;
 RECT 3.25 2.23 3.38 2.36 ;
 RECT 3.245 1.125 3.375 1.255 ;
 RECT 3.245 0.815 3.375 0.945 ;
 RECT 2.77 0.93 2.9 1.06 ;
 RECT 2.77 0.665 2.9 0.795 ;
 RECT 3.635 0.56 3.765 0.69 ;
 RECT 0.475 1.085 0.605 1.215 ;
 RECT 4.105 2.09 4.235 2.22 ;
 RECT 3.635 2.16 3.765 2.29 ;
 RECT 4.105 0.82 4.235 0.95 ;
 RECT 4.105 0.51 4.235 0.64 ;
 RECT 3.635 0.82 3.765 0.95 ;
 RECT 3.635 0.82 3.765 0.95 ;
 RECT 1.28 4.36 1.41 4.49 ;
 RECT 0.475 0.825 0.605 0.955 ;
 RECT 1.87 2.09 2 2.22 ;
 RECT 2.29 2.23 2.42 2.36 ;
 RECT 2.745 3.185 2.875 3.315 ;
 RECT 1.4 0.83 1.53 0.96 ;
 RECT 1.755 3.4 1.885 3.53 ;
 RECT 3.935 1.47 4.065 1.6 ;
 LAYER M1 ;
 RECT 1.395 0.38 1.535 1.02 ;
 RECT 2.29 0.38 2.43 1.385 ;
 RECT 3.63 0.38 3.77 1.02 ;
 RECT 3.24 0.38 3.38 1.385 ;
 RECT 1.395 0.24 3.77 0.38 ;
 RECT 1.275 3.245 1.415 4.56 ;
 RECT 0.93 3.105 1.415 3.245 ;
 RECT 0.895 0.76 1.035 1.45 ;
 RECT 0.895 1.59 1.035 2.29 ;
 RECT 1.44 1.31 1.725 1.45 ;
 RECT 1.44 1.59 1.725 1.62 ;
 RECT 0.895 1.45 1.725 1.59 ;
 RECT 1.865 0.745 2.005 1.64 ;
 RECT 1.865 1.78 2.005 2.29 ;
 RECT 1.865 1.64 2.46 1.78 ;
 RECT 2.2 1.6 2.46 1.64 ;
 RECT 2.2 1.78 2.46 1.83 ;
 END
END LSUPENCLX2

MACRO AODFFARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.64 BY 5.76 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.64 2.96 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.44 1.48 2.91 1.75 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.395 0.495 1.72 0.78 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.56 4.68 7.8 4.92 ;
 RECT 5.71 4.985 5.85 5.4 ;
 RECT 4.875 4.845 5.85 4.985 ;
 RECT 4.805 5.35 5.085 5.49 ;
 RECT 7.65 4.92 7.79 5.4 ;
 RECT 7.65 3.11 8.06 3.25 ;
 RECT 7.65 3.25 7.79 4.68 ;
 RECT 4.875 4.985 5.015 5.35 ;
 RECT 5.71 5.4 7.79 5.54 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.64 0.08 ;
 RECT 5.895 0.08 6.13 0.55 ;
 RECT 2.55 0.08 2.69 1.055 ;
 RECT 0.745 0.08 0.885 0.775 ;
 RECT 3.295 0.08 3.435 0.39 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 8.64 5.84 ;
 RECT 4.165 5.1 4.305 5.68 ;
 RECT 5.27 5.17 5.41 5.68 ;
 RECT 1.47 4.89 1.61 5.68 ;
 RECT 0.685 4.96 0.825 5.68 ;
 RECT 2.96 5.1 3.1 5.68 ;
 RECT 2.59 4.955 2.73 5.68 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.03 3.72 2.36 3.96 ;
 RECT 2.03 3.96 2.17 5.07 ;
 RECT 2.03 3.475 2.17 3.72 ;
 END
 ANTENNADIFFAREA 0.584 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.52 4.04 3.96 4.28 ;
 RECT 3.52 4.28 3.66 5.22 ;
 RECT 3.52 3.485 3.66 4.04 ;
 END
 ANTENNADIFFAREA 0.616 ;
 END QN

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.295 1.73 1.72 2.115 ;
 RECT 1.58 1.585 1.72 1.73 ;
 RECT 6.635 2.46 6.885 2.52 ;
 RECT 3.225 2.34 3.475 2.52 ;
 RECT 2.55 1.98 2.69 2.52 ;
 RECT 1.58 2.115 1.72 2.52 ;
 RECT 1.1 2.52 6.885 2.66 ;
 END
 END VDDG

 OBS
 LAYER PO ;
 RECT 3.15 1.52 3.75 1.62 ;
 RECT 3.585 1.62 3.685 2.68 ;
 RECT 6.265 1.61 6.365 2.68 ;
 RECT 3.15 1.44 3.395 1.52 ;
 RECT 3.15 1.62 3.395 1.69 ;
 RECT 4.515 0.705 4.615 1.165 ;
 RECT 3.65 0.585 3.75 1.165 ;
 RECT 4.515 0.47 4.8 0.705 ;
 RECT 3.585 2.68 6.365 2.78 ;
 RECT 3.65 1.165 4.615 1.265 ;
 RECT 2.3 2.98 2.4 4.395 ;
 RECT 2.3 4.495 2.4 5.455 ;
 RECT 1.715 4.395 2.4 4.495 ;
 RECT 1.715 4.345 1.925 4.395 ;
 RECT 1.715 4.495 1.925 4.58 ;
 RECT 1.81 2.98 1.91 4.345 ;
 RECT 1.81 4.58 1.91 5.455 ;
 RECT 3.305 4.41 3.875 4.49 ;
 RECT 3.305 4.49 4.24 4.51 ;
 RECT 3.775 4.51 4.24 4.72 ;
 RECT 3.775 4.72 3.875 5.635 ;
 RECT 3.305 2.98 3.405 4.41 ;
 RECT 3.305 4.51 3.405 5.635 ;
 RECT 3.775 2.98 3.875 4.41 ;
 RECT 7.135 2.67 7.235 3.085 ;
 RECT 5.62 3.185 5.72 4.195 ;
 RECT 5.62 3.085 7.235 3.185 ;
 RECT 5.96 3.06 6.18 3.085 ;
 RECT 5.96 3.185 6.18 3.3 ;
 RECT 7.015 2.43 7.235 2.67 ;
 RECT 1.445 0.585 2.435 0.685 ;
 RECT 2.335 0.685 2.435 2.465 ;
 RECT 1.445 0.515 1.69 0.585 ;
 RECT 1.445 0.685 1.69 0.765 ;
 RECT 7.015 1.32 8.32 1.42 ;
 RECT 8.22 1.42 8.32 3.76 ;
 RECT 7.24 3.76 8.32 3.86 ;
 RECT 7.24 3.86 7.46 4 ;
 RECT 7.015 1.205 7.235 1.32 ;
 RECT 7.015 1.42 7.235 1.445 ;
 RECT 7.82 2.415 8.04 3.305 ;
 RECT 5.405 0.695 5.505 1.61 ;
 RECT 5.44 1.71 5.54 2.345 ;
 RECT 5.405 1.61 5.54 1.71 ;
 RECT 5.285 0.465 5.525 0.695 ;
 RECT 6.41 4.54 6.51 5.075 ;
 RECT 6.355 5.075 6.585 5.305 ;
 RECT 5.94 3.485 6.04 4.38 ;
 RECT 5.94 4.59 6.04 5.125 ;
 RECT 5.825 4.38 6.06 4.59 ;
 RECT 4.47 1.595 4.57 2.35 ;
 RECT 3.93 1.445 4.175 1.495 ;
 RECT 3.93 1.595 4.175 1.69 ;
 RECT 3.93 1.495 4.57 1.595 ;
 RECT 2.81 0.655 2.91 1.495 ;
 RECT 2.615 1.495 2.91 1.745 ;
 RECT 2.81 1.745 2.91 2.37 ;
 RECT 5.13 3.07 5.23 3.82 ;
 RECT 4.985 3.82 5.23 4.06 ;
 RECT 5.13 4.06 5.23 5.12 ;
 RECT 6.57 1.61 6.835 1.74 ;
 RECT 6.735 1.74 6.835 2.31 ;
 RECT 6.545 0.635 6.645 1.51 ;
 RECT 6.545 1.51 6.835 1.61 ;
 RECT 5.005 0.65 5.105 1.215 ;
 RECT 4.965 1.45 5.065 2.345 ;
 RECT 4.965 1.215 5.195 1.45 ;
 RECT 4.53 3.07 4.63 4.45 ;
 RECT 4.83 4.55 4.93 5.3 ;
 RECT 4.53 4.45 4.93 4.55 ;
 RECT 4.83 5.3 5.06 5.54 ;
 RECT 0.905 2.475 1.325 3.315 ;
 RECT 6.455 4.225 7.09 4.325 ;
 RECT 6.455 3.465 6.555 4.225 ;
 RECT 7.49 2.5 7.59 3.365 ;
 RECT 5.545 4.45 5.645 5.505 ;
 RECT 5.545 5.505 7.09 5.605 ;
 RECT 6.99 4.325 7.09 5.505 ;
 RECT 7.42 2.26 7.64 2.5 ;
 RECT 6.455 3.365 7.59 3.465 ;
 RECT 5.705 0.285 5.805 1.24 ;
 RECT 3.97 0.185 5.805 0.285 ;
 RECT 3.97 0.285 4.07 0.51 ;
 RECT 3.93 0.51 4.175 0.755 ;
 RECT 3.65 1.265 3.75 1.52 ;
 LAYER CO ;
 RECT 2.035 4.075 2.165 4.205 ;
 RECT 4.58 4.77 4.71 4.9 ;
 RECT 6.16 3.765 6.29 3.895 ;
 RECT 5.88 4.42 6.01 4.55 ;
 RECT 2.035 3.55 2.165 3.68 ;
 RECT 4.06 4.54 4.19 4.67 ;
 RECT 0.69 5.015 0.82 5.145 ;
 RECT 0.69 5.275 0.82 5.405 ;
 RECT 0.75 0.59 0.88 0.72 ;
 RECT 0.75 0.33 0.88 0.46 ;
 RECT 5.015 1.26 5.145 1.39 ;
 RECT 6.96 0.88 7.09 1.01 ;
 RECT 6.955 1.84 7.085 1.97 ;
 RECT 3.3 0.21 3.43 0.34 ;
 RECT 6.685 2.465 6.815 2.595 ;
 RECT 5.03 3.875 5.16 4.005 ;
 RECT 3.525 5.025 3.655 5.155 ;
 RECT 6.74 4.77 6.87 4.9 ;
 RECT 6.74 3.825 6.87 3.955 ;
 RECT 4.715 1.925 4.845 2.055 ;
 RECT 4.735 0.88 4.865 1.01 ;
 RECT 4.22 1.94 4.35 2.07 ;
 RECT 4.265 0.88 4.395 1.01 ;
 RECT 3.985 1.49 4.115 1.62 ;
 RECT 3.87 0.905 4 1.035 ;
 RECT 2.675 1.55 2.805 1.68 ;
 RECT 3.985 0.555 4.115 0.685 ;
 RECT 5.275 5.24 5.405 5.37 ;
 RECT 1.56 3.84 1.69 3.97 ;
 RECT 2.035 3.81 2.165 3.94 ;
 RECT 1.56 3.32 1.69 3.45 ;
 RECT 7.865 2.465 7.995 2.595 ;
 RECT 7.465 2.31 7.595 2.44 ;
 RECT 7.06 2.48 7.19 2.61 ;
 RECT 5.34 0.515 5.47 0.645 ;
 RECT 5.945 0.41 6.075 0.54 ;
 RECT 6.625 1.55 6.755 1.68 ;
 RECT 6.405 5.125 6.535 5.255 ;
 RECT 3.525 3.555 3.655 3.685 ;
 RECT 6 3.115 6.13 3.245 ;
 RECT 3.295 2.345 3.425 2.475 ;
 RECT 2.965 5.155 3.095 5.285 ;
 RECT 3.055 3.745 3.185 3.875 ;
 RECT 3.055 4.035 3.185 4.165 ;
 RECT 3.055 3.45 3.185 3.58 ;
 RECT 1.15 3.125 1.28 3.255 ;
 RECT 1.15 2.525 1.28 2.655 ;
 RECT 3.805 1.825 3.935 1.955 ;
 RECT 4.62 0.525 4.75 0.655 ;
 RECT 2.035 4.89 2.165 5.02 ;
 RECT 3.525 3.845 3.655 3.975 ;
 RECT 4.88 5.355 5.01 5.485 ;
 RECT 3.525 4.105 3.655 4.235 ;
 RECT 5.665 1.63 5.795 1.76 ;
 RECT 5.185 1.95 5.315 2.08 ;
 RECT 3.21 1.495 3.34 1.625 ;
 RECT 6.015 1.95 6.145 2.08 ;
 RECT 2.595 5.01 2.725 5.14 ;
 RECT 2.535 3.84 2.665 3.97 ;
 RECT 2.535 3.58 2.665 3.71 ;
 RECT 2.535 3.32 2.665 3.45 ;
 RECT 5.37 3.63 5.5 3.76 ;
 RECT 6.16 4.77 6.29 4.9 ;
 RECT 4.73 3.81 4.86 3.94 ;
 RECT 1.56 3.58 1.69 3.71 ;
 RECT 3.03 1.995 3.16 2.125 ;
 RECT 3.16 0.875 3.29 1.005 ;
 RECT 2.555 2.05 2.685 2.18 ;
 RECT 2.555 0.875 2.685 1.005 ;
 RECT 2.085 0.875 2.215 1.005 ;
 RECT 2.085 2.115 2.215 2.245 ;
 RECT 1.505 0.57 1.635 0.7 ;
 RECT 1.475 4.96 1.605 5.09 ;
 RECT 4.11 3.45 4.24 3.58 ;
 RECT 4.17 5.155 4.3 5.285 ;
 RECT 1.755 4.4 1.885 4.53 ;
 RECT 7.285 3.81 7.415 3.94 ;
 RECT 7.06 1.26 7.19 1.39 ;
 RECT 7.865 3.115 7.995 3.245 ;
 RECT 1.585 2.175 1.715 2.305 ;
 RECT 1.585 1.915 1.715 2.045 ;
 RECT 1.585 1.655 1.715 1.785 ;
 LAYER M1 ;
 RECT 5.115 1.945 6.215 2.085 ;
 RECT 6.95 1.015 7.09 1.255 ;
 RECT 6.95 1.395 7.09 2.035 ;
 RECT 4.965 1.255 7.26 1.395 ;
 RECT 6.89 0.875 7.16 1.015 ;
 RECT 1.555 3.26 1.695 4.04 ;
 RECT 2.53 3.26 2.67 4.04 ;
 RECT 3.05 3.26 3.19 4.235 ;
 RECT 4.105 3.26 4.245 3.655 ;
 RECT 5.365 3.26 5.505 3.815 ;
 RECT 1.085 3.12 5.505 3.26 ;
 RECT 5.935 3.11 6.585 3.25 ;
 RECT 6.445 3.25 6.585 5.12 ;
 RECT 6.335 5.12 6.6 5.26 ;
 RECT 4.55 0.52 5.195 0.66 ;
 RECT 5.055 0.66 5.195 0.97 ;
 RECT 5.055 0.97 6.69 1.11 ;
 RECT 6.55 0.505 7.6 0.645 ;
 RECT 7.46 0.645 7.6 2.51 ;
 RECT 6.55 0.645 6.69 0.97 ;
 RECT 4.725 3.74 4.865 4.235 ;
 RECT 4.575 4.375 4.715 4.815 ;
 RECT 3.885 4.815 4.715 4.955 ;
 RECT 3.24 4.81 3.38 5.385 ;
 RECT 2.31 4.67 3.38 4.81 ;
 RECT 3.24 5.385 4.025 5.525 ;
 RECT 3.885 4.955 4.025 5.385 ;
 RECT 1.75 4.32 1.89 5.395 ;
 RECT 2.31 4.81 2.45 5.395 ;
 RECT 1.75 5.395 2.45 5.535 ;
 RECT 4.575 4.235 6.015 4.375 ;
 RECT 5.875 4.375 6.015 4.6 ;
 RECT 5.335 0.445 5.475 0.69 ;
 RECT 6.27 0.36 6.41 0.69 ;
 RECT 5.335 0.69 6.41 0.83 ;
 RECT 7.86 0.36 8 2.66 ;
 RECT 6.27 0.22 8 0.36 ;
 RECT 1.86 1.01 2 1.195 ;
 RECT 1.86 1.335 2 2.11 ;
 RECT 1.86 2.25 2 2.255 ;
 RECT 1.86 2.11 2.285 2.25 ;
 RECT 1.86 0.87 2.285 1.01 ;
 RECT 2.83 0.67 2.97 1.195 ;
 RECT 1.86 1.195 2.97 1.335 ;
 RECT 4.26 0.36 4.4 1.935 ;
 RECT 2.83 0.53 3.715 0.67 ;
 RECT 3.575 0.22 4.4 0.36 ;
 RECT 3.575 0.36 3.715 0.53 ;
 RECT 4.15 1.935 4.42 2.075 ;
 RECT 3.07 1.63 3.21 1.99 ;
 RECT 3.07 1.475 3.415 1.63 ;
 RECT 3.155 0.825 3.295 1.475 ;
 RECT 2.96 1.99 3.21 2.13 ;
 RECT 4.555 1.625 6.81 1.765 ;
 RECT 4.555 0.975 4.87 1.115 ;
 RECT 4.73 0.805 4.87 0.975 ;
 RECT 4.71 1.765 4.85 1.92 ;
 RECT 6.57 1.545 6.81 1.625 ;
 RECT 4.555 1.115 4.695 1.625 ;
 RECT 4.64 1.92 4.92 2.06 ;
 RECT 6.735 3.775 6.875 3.805 ;
 RECT 6.735 3.945 6.875 4.95 ;
 RECT 6.735 3.805 7.485 3.945 ;
 RECT 4.385 3.55 4.525 3.85 ;
 RECT 4.23 3.99 4.37 4.535 ;
 RECT 3.99 4.535 4.37 4.675 ;
 RECT 4.23 3.85 4.525 3.99 ;
 RECT 4.385 3.41 5.165 3.55 ;
 RECT 5.025 3.955 6.295 4.095 ;
 RECT 6.155 3.71 6.295 3.955 ;
 RECT 6.155 4.095 6.295 4.965 ;
 RECT 5.025 3.55 5.165 3.955 ;
 RECT 3.865 0.5 4.12 0.965 ;
 RECT 3.865 1.96 4.005 2.225 ;
 RECT 3.865 0.965 4.005 1.44 ;
 RECT 3.865 1.67 4.005 1.82 ;
 RECT 3.865 1.44 4.12 1.67 ;
 RECT 3.735 1.82 4.005 1.96 ;
 RECT 3.865 2.32 6.495 2.365 ;
 RECT 3.865 2.225 7.195 2.32 ;
 RECT 7.055 2.32 7.195 2.66 ;
 RECT 6.355 2.18 7.195 2.225 ;
 END
END AODFFARX2

MACRO AODFFNARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.32 BY 5.76 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.32 2.96 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.94 1.475 2.36 1.76 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.77 0.445 1.15 0.825 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.24 4.36 7.48 4.6 ;
 RECT 5.39 4.985 5.53 5.4 ;
 RECT 4.555 4.845 5.53 4.985 ;
 RECT 4.485 5.35 4.76 5.49 ;
 RECT 7.33 4.6 7.47 5.4 ;
 RECT 7.33 3.11 7.74 3.25 ;
 RECT 7.33 3.25 7.47 4.36 ;
 RECT 4.555 4.985 4.695 5.35 ;
 RECT 5.39 5.4 7.47 5.54 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.32 0.08 ;
 RECT 5.575 0.08 5.81 0.55 ;
 RECT 1.98 0.08 2.12 1.055 ;
 RECT 0.365 0.08 0.505 0.775 ;
 RECT 2.725 0.08 2.865 0.39 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 8.32 5.84 ;
 RECT 3.845 5.1 3.985 5.68 ;
 RECT 4.95 5.17 5.09 5.68 ;
 RECT 2.255 4.89 2.395 5.68 ;
 RECT 1.47 4.96 1.61 5.68 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.76 4.04 3 4.28 ;
 RECT 2.815 4.28 2.955 5.07 ;
 RECT 2.815 3.475 2.955 4.04 ;
 END
 ANTENNADIFFAREA 0.471 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.2 3.71 3.64 3.955 ;
 RECT 3.2 3.955 3.34 5.22 ;
 RECT 3.2 3.485 3.34 3.71 ;
 END
 ANTENNADIFFAREA 0.512 ;
 END QN

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.32 3.12 5.185 3.26 ;
 RECT 1.93 4.02 2.07 4.22 ;
 RECT 1.615 3.635 2.07 4.02 ;
 RECT 5.045 3.26 5.185 3.815 ;
 RECT 2.34 3.26 2.48 3.675 ;
 RECT 3.785 3.26 3.925 3.655 ;
 RECT 1.93 3.26 2.07 3.635 ;
 END
 END VDDG

 OBS
 LAYER PO ;
 RECT 6.815 2.67 6.915 3.085 ;
 RECT 5.3 3.185 5.4 4.195 ;
 RECT 5.64 3.06 5.86 3.085 ;
 RECT 5.64 3.185 5.86 3.3 ;
 RECT 5.3 3.085 6.915 3.185 ;
 RECT 6.695 2.43 6.915 2.67 ;
 RECT 4.81 3.07 4.91 3.82 ;
 RECT 4.665 3.82 4.91 4.06 ;
 RECT 4.81 4.06 4.91 5.12 ;
 RECT 1.1 2.475 1.58 3.315 ;
 RECT 6.135 3.465 6.235 4.26 ;
 RECT 7.17 2.5 7.27 3.365 ;
 RECT 5.225 4.45 5.325 5.505 ;
 RECT 5.225 5.505 6.77 5.605 ;
 RECT 6.67 4.36 6.77 5.505 ;
 RECT 6.135 4.26 6.77 4.36 ;
 RECT 7.1 2.26 7.32 2.5 ;
 RECT 6.135 3.365 7.27 3.465 ;
 RECT 7.9 1.42 8 3.76 ;
 RECT 6.695 1.205 6.915 1.32 ;
 RECT 6.695 1.42 6.915 1.445 ;
 RECT 6.695 1.32 8 1.42 ;
 RECT 6.92 3.86 7.14 4 ;
 RECT 6.92 3.76 8 3.86 ;
 RECT 3.5 2.68 6.045 2.78 ;
 RECT 3.5 2.035 3.6 2.68 ;
 RECT 5.945 1.61 6.045 2.68 ;
 RECT 3.5 1.79 3.745 2.035 ;
 RECT 6.09 4.54 6.19 5.075 ;
 RECT 6.035 5.075 6.265 5.305 ;
 RECT 3.55 0.565 3.795 0.71 ;
 RECT 4.195 0.705 4.295 1.255 ;
 RECT 4.195 0.565 4.48 0.705 ;
 RECT 3.54 0.47 4.48 0.565 ;
 RECT 3.54 0.465 4.475 0.47 ;
 RECT 5.385 0.285 5.485 1.24 ;
 RECT 4.15 1.59 4.25 2.35 ;
 RECT 3.08 0.185 5.485 0.285 ;
 RECT 3.08 0.285 3.18 1.49 ;
 RECT 2.58 1.49 4.25 1.59 ;
 RECT 3.015 1.59 3.115 2.365 ;
 RECT 2.58 1.44 2.825 1.49 ;
 RECT 2.58 1.59 2.825 1.69 ;
 RECT 3.455 2.98 3.555 4.49 ;
 RECT 3.455 4.72 3.555 5.635 ;
 RECT 3.455 4.49 3.92 4.72 ;
 RECT 4.21 3.07 4.31 4.45 ;
 RECT 4.51 4.55 4.61 5.3 ;
 RECT 4.21 4.45 4.61 4.55 ;
 RECT 4.51 5.3 4.74 5.54 ;
 RECT 5.62 3.485 5.72 4.38 ;
 RECT 5.62 4.59 5.72 5.125 ;
 RECT 5.505 4.38 5.74 4.59 ;
 RECT 5.085 0.695 5.185 1.61 ;
 RECT 5.12 1.71 5.22 2.345 ;
 RECT 5.085 1.61 5.22 1.71 ;
 RECT 4.965 0.465 5.205 0.695 ;
 RECT 2.595 2.98 2.695 4.495 ;
 RECT 2.595 4.73 2.695 5.455 ;
 RECT 2.5 4.495 2.71 4.73 ;
 RECT 1.765 0.685 1.865 2.465 ;
 RECT 0.84 0.515 1.085 0.585 ;
 RECT 0.84 0.685 1.085 0.765 ;
 RECT 0.84 0.585 1.865 0.685 ;
 RECT 2.24 0.655 2.34 1.495 ;
 RECT 2.045 1.495 2.34 1.745 ;
 RECT 2.24 1.745 2.34 2.37 ;
 RECT 6.25 1.61 6.515 1.74 ;
 RECT 6.415 1.74 6.515 2.31 ;
 RECT 6.225 0.635 6.325 1.51 ;
 RECT 6.225 1.51 6.515 1.61 ;
 RECT 4.685 0.65 4.785 1.215 ;
 RECT 4.645 1.45 4.745 2.345 ;
 RECT 4.645 1.215 4.875 1.45 ;
 RECT 7.5 2.415 7.72 3.305 ;
 LAYER CO ;
 RECT 6.085 5.125 6.215 5.255 ;
 RECT 3.205 3.555 3.335 3.685 ;
 RECT 5.68 3.115 5.81 3.245 ;
 RECT 4.71 3.875 4.84 4.005 ;
 RECT 3.205 5.025 3.335 5.155 ;
 RECT 6.42 4.77 6.55 4.9 ;
 RECT 6.42 3.825 6.55 3.955 ;
 RECT 5.05 3.63 5.18 3.76 ;
 RECT 5.84 4.77 5.97 4.9 ;
 RECT 5.02 0.515 5.15 0.645 ;
 RECT 1.405 3.125 1.535 3.255 ;
 RECT 4.955 5.24 5.085 5.37 ;
 RECT 2.82 3.81 2.95 3.94 ;
 RECT 2.345 3.235 2.475 3.365 ;
 RECT 6.965 3.81 7.095 3.94 ;
 RECT 6.74 1.26 6.87 1.39 ;
 RECT 7.545 3.115 7.675 3.245 ;
 RECT 2.46 1.995 2.59 2.125 ;
 RECT 2.59 0.875 2.72 1.005 ;
 RECT 1.985 2.05 2.115 2.18 ;
 RECT 1.985 0.875 2.115 1.005 ;
 RECT 1.515 0.875 1.645 1.005 ;
 RECT 1.515 2.115 1.645 2.245 ;
 RECT 0.89 0.575 1.02 0.705 ;
 RECT 2.105 1.55 2.235 1.68 ;
 RECT 3.235 1.785 3.365 1.915 ;
 RECT 4.865 1.95 4.995 2.08 ;
 RECT 2.345 3.495 2.475 3.625 ;
 RECT 6.305 1.55 6.435 1.68 ;
 RECT 4.695 1.26 4.825 1.39 ;
 RECT 6.64 0.88 6.77 1.01 ;
 RECT 6.635 1.84 6.765 1.97 ;
 RECT 2.73 0.21 2.86 0.34 ;
 RECT 6.365 2.465 6.495 2.595 ;
 RECT 5.695 1.95 5.825 2.08 ;
 RECT 3.605 0.51 3.735 0.64 ;
 RECT 3.79 3.45 3.92 3.58 ;
 RECT 3.85 5.155 3.98 5.285 ;
 RECT 2.54 4.55 2.67 4.68 ;
 RECT 0.37 0.59 0.5 0.72 ;
 RECT 0.37 0.33 0.5 0.46 ;
 RECT 1.935 4.025 2.065 4.155 ;
 RECT 1.935 3.765 2.065 3.895 ;
 RECT 1.935 3.505 2.065 3.635 ;
 RECT 7.545 2.465 7.675 2.595 ;
 RECT 7.145 2.31 7.275 2.44 ;
 RECT 6.74 2.48 6.87 2.61 ;
 RECT 2.82 4.89 2.95 5.02 ;
 RECT 3.205 3.845 3.335 3.975 ;
 RECT 5.345 1.63 5.475 1.76 ;
 RECT 1.405 2.525 1.535 2.655 ;
 RECT 1.475 5.015 1.605 5.145 ;
 RECT 1.475 5.275 1.605 5.405 ;
 RECT 3.3 0.905 3.43 1.035 ;
 RECT 2.82 4.075 2.95 4.205 ;
 RECT 4.26 4.77 4.39 4.9 ;
 RECT 5.84 3.765 5.97 3.895 ;
 RECT 5.56 4.42 5.69 4.55 ;
 RECT 2.82 3.55 2.95 3.68 ;
 RECT 3.74 4.54 3.87 4.67 ;
 RECT 2.26 4.96 2.39 5.09 ;
 RECT 4.3 0.525 4.43 0.655 ;
 RECT 4.56 5.355 4.69 5.485 ;
 RECT 2.64 1.495 2.77 1.625 ;
 RECT 2.725 2.345 2.855 2.475 ;
 RECT 4.395 1.925 4.525 2.055 ;
 RECT 4.415 0.88 4.545 1.01 ;
 RECT 3.9 1.94 4.03 2.07 ;
 RECT 3.945 0.88 4.075 1.01 ;
 RECT 3.555 1.835 3.685 1.965 ;
 RECT 4.41 3.81 4.54 3.94 ;
 RECT 5.625 0.41 5.755 0.54 ;
 LAYER M1 ;
 RECT 4.795 1.945 5.895 2.085 ;
 RECT 4.23 0.52 4.875 0.66 ;
 RECT 4.735 0.66 4.875 0.97 ;
 RECT 7.14 0.645 7.28 2.51 ;
 RECT 6.23 0.505 7.28 0.645 ;
 RECT 4.735 0.97 6.37 1.11 ;
 RECT 6.23 0.645 6.37 0.97 ;
 RECT 5.015 0.445 5.155 0.69 ;
 RECT 5.95 0.22 7.68 0.36 ;
 RECT 7.54 0.36 7.68 2.66 ;
 RECT 5.95 0.36 6.09 0.69 ;
 RECT 5.015 0.69 6.09 0.83 ;
 RECT 6.63 1.015 6.77 1.255 ;
 RECT 6.63 1.395 6.77 2.035 ;
 RECT 4.645 1.255 6.94 1.395 ;
 RECT 6.57 0.875 6.84 1.015 ;
 RECT 4.405 3.74 4.545 4.235 ;
 RECT 4.255 4.375 4.395 4.815 ;
 RECT 3.565 4.815 4.395 4.955 ;
 RECT 2.535 4.5 2.675 5.4 ;
 RECT 2.535 5.4 3.705 5.54 ;
 RECT 3.565 4.955 3.705 5.4 ;
 RECT 4.255 4.235 5.695 4.375 ;
 RECT 5.555 4.375 5.695 4.6 ;
 RECT 5.615 3.11 6.265 3.25 ;
 RECT 6.125 3.25 6.265 5.12 ;
 RECT 6.015 5.12 6.28 5.26 ;
 RECT 6.415 3.775 6.555 3.805 ;
 RECT 6.415 3.945 6.555 4.95 ;
 RECT 6.415 3.805 7.165 3.945 ;
 RECT 4.065 3.55 4.205 3.85 ;
 RECT 3.91 3.99 4.05 4.535 ;
 RECT 3.67 4.535 4.05 4.675 ;
 RECT 3.91 3.85 4.205 3.99 ;
 RECT 4.065 3.41 4.845 3.55 ;
 RECT 4.705 3.55 4.845 3.955 ;
 RECT 4.705 3.955 5.975 4.095 ;
 RECT 5.835 3.71 5.975 3.955 ;
 RECT 5.835 4.095 5.975 4.965 ;
 RECT 3.295 1.035 3.435 1.78 ;
 RECT 3.6 0.5 3.74 0.505 ;
 RECT 3.6 0.645 3.74 0.895 ;
 RECT 3.23 0.895 3.74 1.005 ;
 RECT 3.23 1.005 3.73 1.035 ;
 RECT 3.51 1.92 3.69 2.015 ;
 RECT 3.165 1.78 3.69 1.92 ;
 RECT 3.53 0.505 3.785 0.645 ;
 RECT 2.26 0.67 2.4 1.195 ;
 RECT 1.29 1.195 2.4 1.335 ;
 RECT 1.29 1.01 1.43 1.195 ;
 RECT 1.29 1.335 1.43 2.11 ;
 RECT 1.29 2.25 1.43 2.255 ;
 RECT 1.29 2.11 1.715 2.25 ;
 RECT 1.29 0.87 1.715 1.01 ;
 RECT 3.94 0.36 4.08 1.935 ;
 RECT 2.26 0.53 3.26 0.67 ;
 RECT 3.12 0.22 4.08 0.36 ;
 RECT 3.12 0.36 3.26 0.53 ;
 RECT 3.83 1.935 4.1 2.075 ;
 RECT 4.235 1.625 6.49 1.765 ;
 RECT 4.235 0.975 4.55 1.115 ;
 RECT 4.41 0.805 4.55 0.975 ;
 RECT 4.39 1.765 4.53 1.92 ;
 RECT 6.25 1.545 6.49 1.625 ;
 RECT 4.235 1.115 4.375 1.625 ;
 RECT 4.32 1.92 4.6 2.06 ;
 RECT 1.345 2.52 6.565 2.66 ;
 RECT 1.98 1.98 2.12 2.52 ;
 RECT 6.315 2.46 6.565 2.52 ;
 RECT 2.655 2.34 2.905 2.52 ;
 RECT 3.205 2.225 6.875 2.32 ;
 RECT 6.735 2.32 6.875 2.66 ;
 RECT 6.035 2.18 6.875 2.225 ;
 RECT 3.205 2.32 6.175 2.365 ;
 RECT 2.39 1.99 3.025 2.06 ;
 RECT 2.5 1.63 2.64 1.99 ;
 RECT 2.39 2.06 3.345 2.13 ;
 RECT 2.5 1.475 2.845 1.63 ;
 RECT 2.585 0.825 2.725 1.475 ;
 RECT 3.205 2.2 3.345 2.225 ;
 RECT 2.885 2.13 3.345 2.2 ;
 END
END AODFFNARX1

MACRO AODFFNARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.64 BY 5.76 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.64 2.96 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.36 1.475 2.68 1.755 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.1 0.51 1.4 0.775 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.56 4.37 7.8 4.6 ;
 RECT 5.71 4.985 5.85 5.4 ;
 RECT 4.875 4.845 5.85 4.985 ;
 RECT 4.805 5.35 5.08 5.49 ;
 RECT 7.65 4.6 7.79 5.4 ;
 RECT 7.65 3.11 8.06 3.25 ;
 RECT 7.65 3.25 7.79 4.37 ;
 RECT 4.875 4.985 5.015 5.35 ;
 RECT 5.71 5.4 7.79 5.54 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.64 0.08 ;
 RECT 5.895 0.08 6.13 0.55 ;
 RECT 2.3 0.08 2.44 1.055 ;
 RECT 0.43 0.08 0.57 0.775 ;
 RECT 3.045 0.08 3.185 0.39 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 8.64 5.84 ;
 RECT 1.16 4.96 1.565 5.68 ;
 RECT 4.165 5.1 4.305 5.68 ;
 RECT 5.27 5.17 5.41 5.68 ;
 RECT 1.83 4.89 1.97 5.68 ;
 RECT 2.95 5.1 3.09 5.68 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.39 3.4 2.68 3.65 ;
 RECT 2.39 3.65 2.53 5.07 ;
 END
 ANTENNADIFFAREA 0.576 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.52 3.72 3.965 3.965 ;
 RECT 3.52 3.965 3.66 5.22 ;
 RECT 3.52 3.485 3.66 3.72 ;
 END
 ANTENNADIFFAREA 0.586 ;
 END QN

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.295 3.635 1.72 4.02 ;
 RECT 1.52 4.02 1.66 4.22 ;
 RECT 1.38 3.12 5.505 3.26 ;
 RECT 5.365 3.26 5.505 3.815 ;
 RECT 1.915 3.26 2.055 4.04 ;
 RECT 4.105 3.26 4.245 3.655 ;
 RECT 2.95 3.26 3.09 4.145 ;
 RECT 1.52 3.26 1.66 3.635 ;
 END
 END VDDG

 OBS
 LAYER PO ;
 RECT 5.405 0.695 5.505 1.61 ;
 RECT 5.44 1.71 5.54 2.345 ;
 RECT 5.405 1.61 5.54 1.71 ;
 RECT 5.285 0.465 5.525 0.695 ;
 RECT 1.115 0.515 1.36 0.58 ;
 RECT 1.115 0.68 1.36 0.765 ;
 RECT 2.085 0.68 2.185 2.465 ;
 RECT 1.115 0.58 2.185 0.68 ;
 RECT 2.175 2.98 2.275 4.345 ;
 RECT 2.175 4.58 2.275 5.455 ;
 RECT 2.075 4.345 2.285 4.41 ;
 RECT 2.075 4.41 2.745 4.51 ;
 RECT 2.075 4.51 2.285 4.58 ;
 RECT 2.645 2.98 2.745 4.41 ;
 RECT 2.645 4.51 2.745 5.455 ;
 RECT 3.3 4.485 3.875 4.49 ;
 RECT 3.3 4.49 4.24 4.585 ;
 RECT 3.775 4.585 4.24 4.72 ;
 RECT 3.775 4.72 3.875 5.635 ;
 RECT 3.3 2.98 3.4 4.485 ;
 RECT 3.3 4.585 3.4 5.635 ;
 RECT 3.775 2.98 3.875 4.485 ;
 RECT 3.82 2.68 6.365 2.78 ;
 RECT 3.82 2.035 3.92 2.68 ;
 RECT 6.265 1.61 6.365 2.68 ;
 RECT 3.82 1.79 4.065 2.035 ;
 RECT 2.56 0.655 2.66 1.495 ;
 RECT 2.365 1.495 2.66 1.745 ;
 RECT 2.56 1.745 2.66 2.37 ;
 RECT 3.87 0.565 4.115 0.71 ;
 RECT 4.515 0.705 4.615 1.255 ;
 RECT 4.515 0.565 4.8 0.705 ;
 RECT 3.83 0.47 4.8 0.565 ;
 RECT 3.83 0.465 4.795 0.47 ;
 RECT 3.4 0.285 3.5 1.49 ;
 RECT 5.705 0.285 5.805 1.24 ;
 RECT 3.4 0.185 5.805 0.285 ;
 RECT 2.9 1.44 3.145 1.49 ;
 RECT 2.9 1.59 3.145 1.69 ;
 RECT 2.9 1.49 4.57 1.59 ;
 RECT 3.335 1.59 3.435 2.405 ;
 RECT 4.47 1.59 4.57 2.35 ;
 RECT 7.82 2.415 8.04 3.305 ;
 RECT 6.41 4.54 6.51 5.075 ;
 RECT 6.355 5.075 6.585 5.305 ;
 RECT 6.57 1.61 6.835 1.74 ;
 RECT 6.735 1.74 6.835 2.31 ;
 RECT 6.545 0.635 6.645 1.51 ;
 RECT 6.545 1.51 6.835 1.61 ;
 RECT 5.005 0.65 5.105 1.215 ;
 RECT 4.965 1.45 5.065 2.345 ;
 RECT 4.965 1.215 5.195 1.45 ;
 RECT 7.015 1.32 8.32 1.42 ;
 RECT 8.22 1.42 8.32 3.76 ;
 RECT 7.24 3.76 8.32 3.86 ;
 RECT 7.24 3.86 7.46 4 ;
 RECT 7.015 1.205 7.235 1.32 ;
 RECT 7.015 1.42 7.235 1.445 ;
 RECT 5.13 3.07 5.23 3.82 ;
 RECT 4.985 3.82 5.23 4.06 ;
 RECT 5.13 4.06 5.23 5.12 ;
 RECT 4.53 3.07 4.63 4.45 ;
 RECT 4.83 4.55 4.93 5.3 ;
 RECT 4.53 4.45 4.93 4.55 ;
 RECT 4.83 5.3 5.06 5.54 ;
 RECT 5.94 3.485 6.04 4.38 ;
 RECT 5.94 4.59 6.04 5.125 ;
 RECT 5.825 4.38 6.06 4.59 ;
 RECT 1.14 2.475 1.62 3.315 ;
 RECT 6.455 4.26 7.09 4.36 ;
 RECT 6.455 3.465 6.555 4.26 ;
 RECT 7.49 2.5 7.59 3.365 ;
 RECT 5.545 4.45 5.645 5.505 ;
 RECT 5.545 5.505 7.09 5.605 ;
 RECT 6.99 4.36 7.09 5.505 ;
 RECT 7.42 2.26 7.64 2.5 ;
 RECT 6.455 3.365 7.59 3.465 ;
 RECT 7.135 2.67 7.235 3.085 ;
 RECT 5.62 3.185 5.72 4.195 ;
 RECT 5.62 3.085 7.235 3.185 ;
 RECT 5.96 3.06 6.18 3.085 ;
 RECT 5.96 3.185 6.18 3.3 ;
 RECT 7.015 2.43 7.235 2.67 ;
 LAYER CO ;
 RECT 1.92 3.58 2.05 3.71 ;
 RECT 2.395 4.075 2.525 4.205 ;
 RECT 4.58 4.77 4.71 4.9 ;
 RECT 1.445 3.125 1.575 3.255 ;
 RECT 1.445 2.525 1.575 2.655 ;
 RECT 2.395 3.55 2.525 3.68 ;
 RECT 4.06 4.54 4.19 4.67 ;
 RECT 1.835 4.96 1.965 5.09 ;
 RECT 4.11 3.45 4.24 3.58 ;
 RECT 4.17 5.155 4.3 5.285 ;
 RECT 2.115 4.4 2.245 4.53 ;
 RECT 5.275 5.24 5.405 5.37 ;
 RECT 1.92 3.84 2.05 3.97 ;
 RECT 2.395 3.81 2.525 3.94 ;
 RECT 0.435 0.59 0.565 0.72 ;
 RECT 0.435 0.33 0.565 0.46 ;
 RECT 1.525 4.025 1.655 4.155 ;
 RECT 1.525 3.765 1.655 3.895 ;
 RECT 1.525 3.505 1.655 3.635 ;
 RECT 4.88 5.355 5.01 5.485 ;
 RECT 6.405 5.125 6.535 5.255 ;
 RECT 3.525 3.555 3.655 3.685 ;
 RECT 5.945 0.41 6.075 0.54 ;
 RECT 6.625 1.55 6.755 1.68 ;
 RECT 5.015 1.26 5.145 1.39 ;
 RECT 6.96 0.88 7.09 1.01 ;
 RECT 6.955 1.84 7.085 1.97 ;
 RECT 3.05 0.21 3.18 0.34 ;
 RECT 6.685 2.465 6.815 2.595 ;
 RECT 6.015 1.95 6.145 2.08 ;
 RECT 4.22 1.94 4.35 2.07 ;
 RECT 4.265 0.88 4.395 1.01 ;
 RECT 1.835 2.115 1.965 2.245 ;
 RECT 1.43 5.275 1.56 5.405 ;
 RECT 7.285 3.81 7.415 3.94 ;
 RECT 7.06 1.26 7.19 1.39 ;
 RECT 7.865 3.115 7.995 3.245 ;
 RECT 7.865 2.465 7.995 2.595 ;
 RECT 7.06 2.48 7.19 2.61 ;
 RECT 2.395 4.89 2.525 5.02 ;
 RECT 3.525 3.845 3.655 3.975 ;
 RECT 5.665 1.63 5.795 1.76 ;
 RECT 5.185 1.95 5.315 2.08 ;
 RECT 6 3.115 6.13 3.245 ;
 RECT 5.03 3.875 5.16 4.005 ;
 RECT 3.525 5.025 3.655 5.155 ;
 RECT 6.74 4.77 6.87 4.9 ;
 RECT 6.74 3.825 6.87 3.955 ;
 RECT 5.37 3.63 5.5 3.76 ;
 RECT 1.165 5.015 1.295 5.145 ;
 RECT 1.165 5.275 1.295 5.405 ;
 RECT 2.955 3.88 3.085 4.01 ;
 RECT 2.955 5.155 3.085 5.285 ;
 RECT 2.955 3.45 3.085 3.58 ;
 RECT 3.925 0.51 4.055 0.64 ;
 RECT 1.43 5.015 1.56 5.145 ;
 RECT 1.92 3.32 2.05 3.45 ;
 RECT 5.34 0.515 5.47 0.645 ;
 RECT 2.96 1.495 3.09 1.625 ;
 RECT 3.045 2.345 3.175 2.475 ;
 RECT 4.715 1.925 4.845 2.055 ;
 RECT 4.735 0.88 4.865 1.01 ;
 RECT 6.16 4.77 6.29 4.9 ;
 RECT 4.73 3.81 4.86 3.94 ;
 RECT 3.875 1.835 4.005 1.965 ;
 RECT 3.62 0.905 3.75 1.035 ;
 RECT 2.78 1.995 2.91 2.125 ;
 RECT 2.91 0.875 3.04 1.005 ;
 RECT 2.305 2.105 2.435 2.235 ;
 RECT 2.305 0.875 2.435 1.005 ;
 RECT 1.835 0.875 1.965 1.005 ;
 RECT 6.16 3.765 6.29 3.895 ;
 RECT 5.88 4.42 6.01 4.55 ;
 RECT 1.175 0.57 1.305 0.7 ;
 RECT 2.425 1.55 2.555 1.68 ;
 RECT 3.555 1.785 3.685 1.915 ;
 RECT 4.62 0.525 4.75 0.655 ;
 RECT 7.465 2.31 7.595 2.44 ;
 LAYER M1 ;
 RECT 5.935 3.11 6.585 3.25 ;
 RECT 6.445 3.25 6.585 5.12 ;
 RECT 6.335 5.12 6.6 5.26 ;
 RECT 2.11 4.32 2.25 5.21 ;
 RECT 3.23 4.735 3.37 5.4 ;
 RECT 2.67 4.595 3.37 4.735 ;
 RECT 2.67 4.735 2.81 5.21 ;
 RECT 2.11 5.21 2.81 5.35 ;
 RECT 4.725 3.74 4.865 4.235 ;
 RECT 4.575 4.375 4.715 4.815 ;
 RECT 3.885 4.815 4.715 4.955 ;
 RECT 3.23 5.4 4.025 5.54 ;
 RECT 3.885 4.955 4.025 5.4 ;
 RECT 4.575 4.235 6.015 4.375 ;
 RECT 5.875 4.375 6.015 4.6 ;
 RECT 5.335 0.445 5.475 0.69 ;
 RECT 7.86 0.36 8 2.66 ;
 RECT 6.27 0.22 8 0.36 ;
 RECT 6.27 0.36 6.41 0.69 ;
 RECT 5.335 0.69 6.41 0.83 ;
 RECT 5.115 1.945 6.215 2.085 ;
 RECT 4.55 0.52 5.195 0.66 ;
 RECT 5.055 0.66 5.195 0.97 ;
 RECT 7.46 0.645 7.6 2.51 ;
 RECT 6.55 0.505 7.6 0.645 ;
 RECT 5.055 0.97 6.69 1.11 ;
 RECT 6.55 0.645 6.69 0.97 ;
 RECT 6.95 1.015 7.09 1.255 ;
 RECT 6.95 1.395 7.09 2.035 ;
 RECT 6.89 0.875 7.16 1.015 ;
 RECT 4.965 1.255 7.26 1.395 ;
 RECT 1.61 1.01 1.75 1.195 ;
 RECT 1.61 1.335 1.75 2.11 ;
 RECT 1.61 2.25 1.75 2.255 ;
 RECT 1.61 2.11 2.035 2.25 ;
 RECT 1.61 0.87 2.035 1.01 ;
 RECT 1.61 1.195 2.72 1.335 ;
 RECT 2.58 0.67 2.72 1.195 ;
 RECT 4.26 0.36 4.4 1.935 ;
 RECT 2.58 0.53 3.58 0.67 ;
 RECT 3.44 0.22 4.4 0.36 ;
 RECT 3.44 0.36 3.58 0.53 ;
 RECT 4.15 1.935 4.42 2.075 ;
 RECT 4.68 1.625 6.81 1.765 ;
 RECT 4.73 0.805 4.87 0.975 ;
 RECT 4.68 0.975 4.87 1.115 ;
 RECT 4.71 1.765 4.85 1.92 ;
 RECT 6.57 1.545 6.81 1.625 ;
 RECT 4.64 1.92 4.92 2.06 ;
 RECT 4.68 1.115 4.82 1.625 ;
 RECT 6.735 3.775 6.875 3.805 ;
 RECT 6.735 3.945 6.875 4.95 ;
 RECT 6.735 3.805 7.485 3.945 ;
 RECT 4.385 3.55 4.525 3.85 ;
 RECT 4.23 3.99 4.37 4.535 ;
 RECT 3.99 4.535 4.37 4.675 ;
 RECT 4.23 3.85 4.525 3.99 ;
 RECT 4.385 3.41 5.165 3.55 ;
 RECT 5.025 3.55 5.165 3.955 ;
 RECT 5.025 3.955 6.295 4.095 ;
 RECT 6.155 3.71 6.295 3.955 ;
 RECT 6.155 4.095 6.295 4.965 ;
 RECT 3.615 1.035 3.755 1.78 ;
 RECT 3.92 0.5 4.06 0.505 ;
 RECT 3.92 0.645 4.06 0.895 ;
 RECT 3.83 1.92 4.01 2.015 ;
 RECT 3.485 1.78 4.01 1.92 ;
 RECT 3.85 0.505 4.105 0.645 ;
 RECT 3.55 0.895 4.06 1.035 ;
 RECT 1.365 2.52 6.885 2.66 ;
 RECT 2.3 2.055 2.44 2.52 ;
 RECT 6.635 2.46 6.885 2.52 ;
 RECT 2.975 2.34 3.225 2.52 ;
 RECT 3.525 2.225 7.195 2.32 ;
 RECT 7.055 2.32 7.195 2.66 ;
 RECT 6.355 2.18 7.195 2.225 ;
 RECT 3.525 2.32 6.495 2.365 ;
 RECT 2.73 1.99 3.345 2.06 ;
 RECT 2.82 1.63 2.96 1.99 ;
 RECT 2.73 2.06 3.665 2.13 ;
 RECT 2.82 1.475 3.165 1.63 ;
 RECT 2.905 0.825 3.045 1.475 ;
 RECT 3.525 2.2 3.665 2.225 ;
 RECT 3.205 2.13 3.665 2.2 ;
 END
END AODFFNARX2

MACRO AOINVX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 5.76 ;
 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.825 1.68 2.52 1.84 ;
 RECT 2.265 1.84 2.52 2.12 ;
 RECT 2.265 1.65 2.52 1.68 ;
 END
 END VDDG

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.705 0.84 2.04 1.08 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END INP

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 2.31 0.08 2.45 0.765 ;
 RECT 1.9 0.08 2.04 0.53 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 3.84 5.84 ;
 RECT 2.31 4.975 2.45 5.68 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.845 2.96 ;
 END
 END VDD

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 1.48 1.565 1.72 ;
 RECT 1.425 1.72 1.565 1.89 ;
 RECT 1.425 0.26 1.565 1.48 ;
 END
 ANTENNADIFFAREA 0.213 ;
 END ZN

 OBS
 LAYER PO ;
 RECT 1.68 0.1 1.78 2.185 ;
 RECT 1.725 0.845 1.955 1.075 ;
 LAYER CO ;
 RECT 2.315 5.31 2.445 5.44 ;
 RECT 2.315 5.035 2.445 5.165 ;
 RECT 1.905 0.33 2.035 0.46 ;
 RECT 1.905 1.695 2.035 1.825 ;
 RECT 1.775 0.895 1.905 1.025 ;
 RECT 1.43 1.685 1.56 1.815 ;
 RECT 1.43 0.33 1.56 0.46 ;
 RECT 2.315 0.305 2.445 0.435 ;
 RECT 2.315 0.565 2.445 0.695 ;
 RECT 2.315 1.69 2.445 1.82 ;
 RECT 2.315 1.95 2.445 2.08 ;
 END
END AOINVX1

MACRO AOINVX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 5.76 ;
 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.825 1.68 2.46 1.76 ;
 RECT 2.255 1.84 2.585 2.15 ;
 RECT 1.825 1.76 2.585 1.84 ;
 RECT 2.31 1.62 2.45 1.68 ;
 END
 END VDDG

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.74 0.84 2.04 1.13 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END INP

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 2.31 0.08 2.45 0.765 ;
 RECT 1.9 0.08 2.04 0.53 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 3.84 5.84 ;
 RECT 2.31 4.975 2.45 5.68 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 END
 END VDD

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 1.48 1.565 1.72 ;
 RECT 1.425 1.72 1.565 1.89 ;
 RECT 1.425 0.26 1.565 1.48 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END ZN

 OBS
 LAYER PO ;
 RECT 1.68 0.1 1.78 2.745 ;
 RECT 1.775 0.89 2.005 1.12 ;
 LAYER CO ;
 RECT 2.315 5.31 2.445 5.44 ;
 RECT 2.315 5.035 2.445 5.165 ;
 RECT 1.905 0.33 2.035 0.46 ;
 RECT 1.905 1.695 2.035 1.825 ;
 RECT 1.825 0.94 1.955 1.07 ;
 RECT 1.43 1.685 1.56 1.815 ;
 RECT 1.43 0.33 1.56 0.46 ;
 RECT 2.315 0.305 2.445 0.435 ;
 RECT 2.315 0.565 2.445 0.695 ;
 RECT 2.315 1.69 2.445 1.82 ;
 RECT 2.315 1.95 2.445 2.08 ;
 END
END AOINVX2

MACRO AOINVX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 5.76 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.475 1.37 1.72 1.72 ;
 RECT 0.305 1.23 1.855 1.37 ;
 END
 ANTENNAGATEAREA 0.644 ;
 END INP

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.995 1.135 2.385 1.43 ;
 RECT 0.115 0.94 2.135 1.08 ;
 RECT 1.055 0.625 1.195 0.94 ;
 RECT 1.995 1.08 2.135 1.135 ;
 RECT 1.995 0.64 2.135 0.94 ;
 RECT 1.995 2 2.135 2.04 ;
 RECT 1.005 1.86 2.135 2 ;
 RECT 0.115 0.64 0.255 0.94 ;
 RECT 1.005 1.855 1.145 1.86 ;
 RECT 0.115 1.715 1.145 1.855 ;
 RECT 0.115 1.855 0.255 2.31 ;
 RECT 1.995 1.43 2.135 1.585 ;
 RECT 1.975 1.585 2.135 1.86 ;
 END
 ANTENNADIFFAREA 1.562 ;
 END ZN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 2.605 0.08 2.745 0.805 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 1.525 0.08 1.665 0.77 ;
 RECT 0.585 0.08 0.725 0.77 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 3.2 5.84 ;
 RECT 2.605 4.955 2.745 5.68 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 2.595 1.93 2.755 1.975 ;
 RECT 2.455 1.975 2.97 2.425 ;
 RECT 0.51 2.425 2.97 2.585 ;
 END
 END VDDG

 OBS
 LAYER PO ;
 RECT 0.84 0.275 0.94 1.185 ;
 RECT 0.84 1.415 0.94 2.79 ;
 RECT 0.755 1.185 0.985 1.415 ;
 RECT 1.78 0.275 1.88 1.185 ;
 RECT 1.625 1.185 1.88 1.415 ;
 RECT 1.78 1.415 1.88 2.79 ;
 RECT 1.31 0.275 1.41 1.185 ;
 RECT 1.31 1.415 1.41 2.79 ;
 RECT 1.2 1.185 1.43 1.415 ;
 RECT 0.37 0.275 0.47 1.185 ;
 RECT 0.37 1.415 0.47 2.79 ;
 RECT 0.305 1.185 0.535 1.415 ;
 LAYER CO ;
 RECT 2.61 0.625 2.74 0.755 ;
 RECT 2.61 2.025 2.74 2.155 ;
 RECT 2.61 2.295 2.74 2.425 ;
 RECT 2.61 0.355 2.74 0.485 ;
 RECT 0.59 0.59 0.72 0.72 ;
 RECT 0.59 2.43 0.72 2.56 ;
 RECT 0.355 1.235 0.485 1.365 ;
 RECT 0.805 1.235 0.935 1.365 ;
 RECT 0.12 2.13 0.25 2.26 ;
 RECT 1.53 2.44 1.66 2.57 ;
 RECT 1.675 1.235 1.805 1.365 ;
 RECT 2 1.86 2.13 1.99 ;
 RECT 1.06 1.865 1.19 1.995 ;
 RECT 1.25 1.235 1.38 1.365 ;
 RECT 0.12 1.86 0.25 1.99 ;
 RECT 2 0.69 2.13 0.82 ;
 RECT 0.12 0.69 0.25 0.82 ;
 RECT 1.06 0.675 1.19 0.805 ;
 RECT 1.53 0.59 1.66 0.72 ;
 RECT 2.61 5.005 2.74 5.135 ;
 RECT 2.61 5.275 2.74 5.405 ;
 END
END AOINVX4

MACRO BUSKP
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.595 1.45 1.735 1.82 ;
 RECT 0.51 1.15 0.93 1.31 ;
 RECT 1.97 0.32 2.11 1.31 ;
 RECT 0.51 1.31 2.11 1.45 ;
 END
 ANTENNADIFFAREA 0.214 ;
 END INP

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 2.65 0.08 2.79 0.825 ;
 RECT 0.69 0.08 0.83 0.55 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 0.7 1.59 0.84 2.8 ;
 RECT 2.625 2.12 2.765 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.47 0.15 0.57 1.22 ;
 RECT 0.47 1.22 0.755 1.45 ;
 RECT 0.47 1.45 0.57 2.43 ;
 RECT 0.945 0.825 1.175 0.925 ;
 RECT 0.945 0.725 1.85 0.825 ;
 RECT 1.5 0.15 1.85 0.725 ;
 RECT 1.375 0.825 1.475 1.99 ;
 RECT 0.945 0.14 1.295 0.725 ;
 RECT 1.075 0.925 1.175 1.99 ;
 LAYER CO ;
 RECT 0.575 1.27 0.705 1.4 ;
 RECT 0.995 0.745 1.125 0.875 ;
 RECT 2.63 2.43 2.76 2.56 ;
 RECT 2.655 0.37 2.785 0.5 ;
 RECT 2.655 0.64 2.785 0.77 ;
 RECT 2.63 2.17 2.76 2.3 ;
 RECT 1.975 0.37 2.105 0.5 ;
 RECT 0.695 0.37 0.825 0.5 ;
 RECT 0.22 0.37 0.35 0.5 ;
 RECT 1.6 1.64 1.73 1.77 ;
 RECT 0.705 2.065 0.835 2.195 ;
 RECT 0.705 1.64 0.835 1.77 ;
 RECT 0.22 1.64 0.35 1.77 ;
 RECT 0.22 2.065 0.35 2.195 ;
 LAYER M1 ;
 RECT 0.215 0.32 0.355 2.245 ;
 RECT 0.305 0.74 1.175 0.88 ;
 END
END BUSKP

MACRO CLOAD1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.24 BY 2.88 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.34 1.125 0.815 1.465 ;
 END
 ANTENNAGATEAREA 0.161 ;
 END INP

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.24 2.96 ;
 RECT 0.49 1.605 0.63 2.8 ;
 RECT 0.99 1.615 1.13 2.8 ;
 RECT 1.58 1.905 1.72 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.24 0.08 ;
 RECT 1.58 0.08 1.72 0.84 ;
 RECT 0.99 0.08 1.13 0.845 ;
 RECT 0.49 0.08 0.63 0.845 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.765 0.26 0.865 2.745 ;
 RECT 0.585 1.125 0.815 1.355 ;
 LAYER CO ;
 RECT 1.585 0.64 1.715 0.77 ;
 RECT 1.585 0.37 1.715 0.5 ;
 RECT 1.585 2.245 1.715 2.375 ;
 RECT 1.585 1.975 1.715 2.105 ;
 RECT 0.995 1.945 1.125 2.075 ;
 RECT 0.995 2.255 1.125 2.385 ;
 RECT 0.495 0.645 0.625 0.775 ;
 RECT 0.635 1.175 0.765 1.305 ;
 RECT 0.995 1.685 1.125 1.815 ;
 RECT 0.495 2.255 0.625 2.385 ;
 RECT 0.495 1.945 0.625 2.075 ;
 RECT 0.495 1.675 0.625 1.805 ;
 RECT 0.995 0.645 1.125 0.775 ;
 END
END CLOAD1

MACRO DCAP
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 1.92 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 1.92 0.08 ;
 RECT 1.37 0.08 1.51 0.755 ;
 RECT 0.38 0.08 0.52 0.5 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 1.92 2.96 ;
 RECT 0.385 2.17 0.525 2.8 ;
 RECT 1.37 1.835 1.51 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.64 1.63 0.74 2.785 ;
 RECT 0.37 1.4 0.6 1.53 ;
 RECT 0.37 1.53 0.74 1.63 ;
 RECT 0.64 0.09 0.74 1.095 ;
 RECT 0.81 1.195 1.04 1.325 ;
 RECT 0.64 1.095 1.04 1.195 ;
 LAYER CO ;
 RECT 0.42 1.45 0.55 1.58 ;
 RECT 0.86 1.145 0.99 1.275 ;
 RECT 1.375 1.885 1.505 2.015 ;
 RECT 1.375 0.315 1.505 0.445 ;
 RECT 1.375 2.175 1.505 2.305 ;
 RECT 0.86 2.215 0.99 2.345 ;
 RECT 0.39 2.22 0.52 2.35 ;
 RECT 1.375 0.575 1.505 0.705 ;
 RECT 0.865 0.39 0.995 0.52 ;
 RECT 0.385 0.32 0.515 0.45 ;
 LAYER M1 ;
 RECT 0.855 1.095 0.995 2.395 ;
 RECT 0.415 0.785 0.555 1.64 ;
 RECT 0.86 0.34 1 0.645 ;
 RECT 0.415 0.645 1 0.785 ;
 END
END DCAP

MACRO DHFILLHLH2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 0.64 BY 5.76 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 0.64 2.96 ;
 RECT 0.265 2.96 0.405 3.67 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 0.64 0.08 ;
 RECT 0.265 0.08 0.405 0.785 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 0.64 5.84 ;
 RECT 0.265 4.975 0.405 5.68 ;
 END
 END VDD

 OBS
 LAYER CO ;
 RECT 0.27 0.585 0.4 0.715 ;
 RECT 0.27 0.305 0.4 0.435 ;
 RECT 0.27 3.185 0.4 3.315 ;
 RECT 0.27 3.465 0.4 3.595 ;
 RECT 0.27 5.045 0.4 5.175 ;
 RECT 0.27 5.325 0.4 5.455 ;
 END
END DHFILLHLH2

MACRO DHFILLHLHLS11
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 5.76 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 1.82 2.96 2.24 3.645 ;
 END
 END VSS

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 3.52 5.2 ;
 RECT 1.43 4.26 1.85 4.665 ;
 RECT 1.575 4.665 1.715 5.04 ;
 END
 END VDDL

 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 1.73 0.08 1.87 1.025 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 3.52 5.84 ;
 END
 END VDDH

 OBS
 LAYER CO ;
 RECT 2.105 3.185 2.235 3.315 ;
 RECT 2.105 3.445 2.235 3.575 ;
 RECT 1.735 0.565 1.865 0.695 ;
 RECT 1.735 0.825 1.865 0.955 ;
 RECT 1.585 4.3 1.715 4.43 ;
 RECT 1.825 3.185 1.955 3.315 ;
 RECT 1.825 3.445 1.955 3.575 ;
 END
END DHFILLHLHLS11

MACRO DHFILLLHL2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 0.64 BY 5.76 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 0.64 2.96 ;
 RECT 0.255 2.96 0.395 3.125 ;
 RECT 0.255 2.565 0.395 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 0.64 0.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 0.64 5.84 ;
 END
 END VSS

 OBS
 LAYER CO ;
 RECT 0.26 2.625 0.39 2.755 ;
 RECT 0.26 2.895 0.39 3.025 ;
 END
END DHFILLLHL2

MACRO HEAD2X16
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.52 BY 5.76 ;
 PIN SLEEP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.38 0.345 0.805 0.78 ;
 END
 ANTENNAGATEAREA 0.072 ;
 END SLEEP

 PIN SLEEPOUT
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.425 0.98 2.915 1.18 ;
 RECT 2.425 0.81 2.915 0.84 ;
 RECT 7.77 0.98 7.91 2.295 ;
 RECT 7.77 0.315 7.91 0.84 ;
 RECT 8.71 0.98 8.85 2.295 ;
 RECT 8.71 0.315 8.85 0.84 ;
 RECT 6.83 0.98 6.97 2.295 ;
 RECT 6.83 0.315 6.97 0.84 ;
 RECT 3.07 0.98 3.21 2.295 ;
 RECT 3.07 0.315 3.21 0.84 ;
 RECT 2.13 0.98 2.27 2.29 ;
 RECT 2.13 0.84 8.855 0.98 ;
 RECT 2.13 0.315 2.27 0.84 ;
 RECT 4.01 0.98 4.15 2.295 ;
 RECT 4.01 0.315 4.15 0.84 ;
 RECT 4.95 0.98 5.09 2.295 ;
 RECT 4.95 0.315 5.09 0.84 ;
 RECT 5.89 0.98 6.03 2.29 ;
 RECT 5.89 0.315 6.03 0.84 ;
 END
 ANTENNADIFFAREA 4.72 ;
 END SLEEPOUT

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.52 2.96 ;
 RECT 1.185 2.96 1.325 4.01 ;
 RECT 2.125 2.96 2.265 3.95 ;
 RECT 3.065 2.96 3.205 3.95 ;
 RECT 4.005 2.96 4.145 3.95 ;
 RECT 4.945 2.96 5.085 3.95 ;
 RECT 6.825 2.96 6.965 3.95 ;
 RECT 5.885 2.96 6.025 3.95 ;
 RECT 8.705 2.96 8.845 3.95 ;
 RECT 7.765 2.96 7.905 3.95 ;
 END
 END VDD

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0.615 4.275 9.785 4.475 ;
 RECT 1.62 3.33 1.985 3.725 ;
 RECT 0.615 3.485 0.815 4.275 ;
 RECT 2.595 3.335 2.735 4.275 ;
 RECT 3.535 3.335 3.675 4.275 ;
 RECT 4.475 3.335 4.615 4.275 ;
 RECT 5.415 3.335 5.555 4.275 ;
 RECT 7.295 3.335 7.435 4.275 ;
 RECT 8.235 3.335 8.375 4.275 ;
 RECT 6.355 3.335 6.495 4.275 ;
 RECT 9.585 3.73 9.785 4.275 ;
 RECT 9.41 3.415 9.78 3.42 ;
 RECT 9.41 3.42 9.785 3.73 ;
 RECT 1.695 3.965 1.895 4.275 ;
 RECT 1.62 3.725 1.895 3.965 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.52 0.08 ;
 RECT 9.185 0.08 9.325 0.67 ;
 RECT 2.6 0.08 2.74 0.67 ;
 RECT 3.54 0.08 3.68 0.67 ;
 RECT 7.3 0.08 7.44 0.67 ;
 RECT 8.24 0.08 8.38 0.67 ;
 RECT 10.915 0.08 11.115 1.01 ;
 RECT 4.48 0.08 4.62 0.67 ;
 RECT 6.36 0.08 6.5 0.67 ;
 RECT 5.42 0.08 5.56 0.67 ;
 RECT 1.66 0.08 1.8 0.67 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 11.52 5.84 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.595 1.025 0.695 3 ;
 RECT 7.55 2.99 7.65 3 ;
 RECT 7.55 3.1 7.65 4.48 ;
 RECT 5.2 3.1 5.3 4.48 ;
 RECT 8.49 3.1 8.59 4.48 ;
 RECT 5.67 2.99 5.77 3 ;
 RECT 5.67 3.1 5.77 4.48 ;
 RECT 6.14 2.99 6.24 3 ;
 RECT 6.14 3.1 6.24 4.48 ;
 RECT 8.02 2.99 8.12 3 ;
 RECT 8.02 3.1 8.12 4.48 ;
 RECT 6.61 3.1 6.71 4.48 ;
 RECT 7.08 3.1 7.18 4.48 ;
 RECT 4.73 3.1 4.83 4.48 ;
 RECT 4.26 3.1 4.36 4.48 ;
 RECT 3.32 3.1 3.42 4.48 ;
 RECT 3.79 3.1 3.89 4.48 ;
 RECT 2.38 3.1 2.48 4.48 ;
 RECT 2.85 3.1 2.95 4.48 ;
 RECT 1.44 3.1 1.54 4.48 ;
 RECT 1.91 3.1 2.01 4.48 ;
 RECT 0.595 3.1 0.695 3.105 ;
 RECT 1.025 0.87 1.255 0.925 ;
 RECT 1.025 1.025 1.255 1.08 ;
 RECT 0.595 0.925 1.255 1.025 ;
 RECT 0.595 3 8.59 3.1 ;
 RECT 1.915 1.105 2.015 1.36 ;
 RECT 1.915 1.46 2.015 2.81 ;
 RECT 8.965 0.095 9.065 1.36 ;
 RECT 8.965 1.46 9.065 2.81 ;
 RECT 6.615 0.095 6.715 1.36 ;
 RECT 6.615 1.46 6.715 2.81 ;
 RECT 8.495 0.095 8.595 1.36 ;
 RECT 8.495 1.46 8.595 2.81 ;
 RECT 8.025 0.095 8.125 1.36 ;
 RECT 8.025 1.46 8.125 2.81 ;
 RECT 7.555 0.095 7.655 1.36 ;
 RECT 7.555 1.46 7.655 2.81 ;
 RECT 7.085 0.095 7.185 1.36 ;
 RECT 7.085 1.46 7.185 2.81 ;
 RECT 6.145 0.095 6.245 1.36 ;
 RECT 6.145 1.46 6.245 2.81 ;
 RECT 5.675 0.095 5.775 1.36 ;
 RECT 5.675 1.46 5.775 2.81 ;
 RECT 5.205 0.095 5.305 1.36 ;
 RECT 5.205 1.46 5.305 2.81 ;
 RECT 4.735 0.095 4.835 1.36 ;
 RECT 4.735 1.46 4.835 2.81 ;
 RECT 4.265 0.095 4.365 1.36 ;
 RECT 4.265 1.46 4.365 2.81 ;
 RECT 3.795 0.095 3.895 1.36 ;
 RECT 3.795 1.46 3.895 2.81 ;
 RECT 2.385 0.095 2.485 1.36 ;
 RECT 2.385 1.46 2.485 2.81 ;
 RECT 3.325 0.095 3.425 1.36 ;
 RECT 3.325 1.46 3.425 2.81 ;
 RECT 2.855 0.095 2.955 1.36 ;
 RECT 2.855 1.46 2.955 2.81 ;
 RECT 1.915 0.095 2.015 0.895 ;
 RECT 1.75 0.895 2.015 1.105 ;
 RECT 1.91 1.36 9.065 1.46 ;
 RECT 1.445 0.095 1.545 0.59 ;
 RECT 0.515 0.59 1.545 0.69 ;
 RECT 1.445 0.69 1.545 2.81 ;
 RECT 0.52 0.485 0.75 0.59 ;
 RECT 0.52 0.69 0.75 0.695 ;
 RECT 9.6 2.655 9.7 3.445 ;
 RECT 9.6 3.655 9.7 3.71 ;
 RECT 9.54 2.445 9.77 2.655 ;
 RECT 9.535 3.445 9.765 3.655 ;
 LAYER CO ;
 RECT 3.075 2.115 3.205 2.245 ;
 RECT 3.545 2.315 3.675 2.445 ;
 RECT 1.665 0.405 1.795 0.535 ;
 RECT 1.665 2.315 1.795 2.445 ;
 RECT 2.605 2.315 2.735 2.445 ;
 RECT 3.545 0.405 3.675 0.535 ;
 RECT 2.13 3.385 2.26 3.515 ;
 RECT 1.19 3.645 1.32 3.775 ;
 RECT 10.95 0.685 11.08 0.815 ;
 RECT 10.95 0.425 11.08 0.555 ;
 RECT 0.65 3.91 0.78 4.04 ;
 RECT 0.65 3.65 0.78 3.78 ;
 RECT 6.835 2.04 6.965 2.17 ;
 RECT 5.895 0.43 6.025 0.56 ;
 RECT 9.19 2.315 9.32 2.445 ;
 RECT 9.19 0.405 9.32 0.535 ;
 RECT 5.895 2.11 6.025 2.24 ;
 RECT 7.305 0.405 7.435 0.535 ;
 RECT 8.245 0.405 8.375 0.535 ;
 RECT 8.715 2.115 8.845 2.245 ;
 RECT 8.715 0.405 8.845 0.535 ;
 RECT 6.835 0.445 6.965 0.575 ;
 RECT 8.245 2.315 8.375 2.445 ;
 RECT 7.305 2.315 7.435 2.445 ;
 RECT 7.775 2.115 7.905 2.245 ;
 RECT 7.775 0.405 7.905 0.535 ;
 RECT 6.365 0.405 6.495 0.535 ;
 RECT 6.365 2.315 6.495 2.445 ;
 RECT 6.36 3.385 6.49 3.515 ;
 RECT 6.36 3.645 6.49 3.775 ;
 RECT 7.77 3.385 7.9 3.515 ;
 RECT 7.3 3.645 7.43 3.775 ;
 RECT 7.77 3.645 7.9 3.775 ;
 RECT 5.89 3.385 6.02 3.515 ;
 RECT 9.59 2.485 9.72 2.615 ;
 RECT 1.075 0.91 1.205 1.04 ;
 RECT 1.8 0.935 1.93 1.065 ;
 RECT 0.57 0.525 0.7 0.655 ;
 RECT 9.585 3.485 9.715 3.615 ;
 RECT 5.42 3.385 5.55 3.515 ;
 RECT 8.24 3.385 8.37 3.515 ;
 RECT 6.83 3.385 6.96 3.515 ;
 RECT 8.71 3.385 8.84 3.515 ;
 RECT 5.42 3.645 5.55 3.775 ;
 RECT 8.24 3.645 8.37 3.775 ;
 RECT 6.83 3.645 6.96 3.775 ;
 RECT 8.71 3.645 8.84 3.775 ;
 RECT 5.89 3.645 6.02 3.775 ;
 RECT 7.3 3.385 7.43 3.515 ;
 RECT 4.48 3.385 4.61 3.515 ;
 RECT 4.95 3.385 5.08 3.515 ;
 RECT 4.48 3.645 4.61 3.775 ;
 RECT 4.95 3.645 5.08 3.775 ;
 RECT 3.54 3.385 3.67 3.515 ;
 RECT 4.01 3.385 4.14 3.515 ;
 RECT 3.54 3.645 3.67 3.775 ;
 RECT 4.01 3.645 4.14 3.775 ;
 RECT 2.6 3.385 2.73 3.515 ;
 RECT 3.07 3.385 3.2 3.515 ;
 RECT 2.6 3.645 2.73 3.775 ;
 RECT 3.07 3.645 3.2 3.775 ;
 RECT 5.425 2.315 5.555 2.445 ;
 RECT 5.425 0.405 5.555 0.535 ;
 RECT 4.485 0.405 4.615 0.535 ;
 RECT 4.955 2.115 5.085 2.245 ;
 RECT 4.955 0.405 5.085 0.535 ;
 RECT 4.485 2.315 4.615 2.445 ;
 RECT 4.015 2.115 4.145 2.245 ;
 RECT 4.015 0.405 4.145 0.535 ;
 RECT 3.075 0.405 3.205 0.535 ;
 RECT 2.605 0.405 2.735 0.535 ;
 RECT 2.135 2.11 2.265 2.24 ;
 RECT 1.19 2.32 1.32 2.45 ;
 RECT 2.135 0.405 2.265 0.535 ;
 RECT 1.66 3.385 1.79 3.515 ;
 RECT 1.66 3.645 1.79 3.775 ;
 RECT 2.13 3.645 2.26 3.775 ;
 RECT 1.19 0.335 1.32 0.465 ;
 RECT 1.19 3.385 1.32 3.515 ;
 LAYER M1 ;
 RECT 8.24 2.26 8.38 2.52 ;
 RECT 7.3 2.26 7.44 2.52 ;
 RECT 6.36 2.265 6.5 2.52 ;
 RECT 5.42 2.26 5.56 2.52 ;
 RECT 4.48 2.26 4.62 2.52 ;
 RECT 3.54 2.26 3.68 2.52 ;
 RECT 2.6 2.265 2.74 2.52 ;
 RECT 1.66 2.265 1.8 2.52 ;
 RECT 9.185 2.26 9.325 2.52 ;
 RECT 9.49 2.34 9.835 2.52 ;
 RECT 1.655 2.52 9.835 2.66 ;
 RECT 0.97 0.81 1.325 0.87 ;
 RECT 0.97 1.01 1.325 1.145 ;
 RECT 1.185 0.24 1.325 0.81 ;
 RECT 1.185 1.145 1.325 2.555 ;
 RECT 0.97 0.87 1.985 1.01 ;
 RECT 1.63 0.835 1.985 0.87 ;
 RECT 1.63 1.01 1.985 1.19 ;
 END
END HEAD2X16

MACRO HEAD2X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 5.76 ;
 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0.785 4.345 3.045 4.545 ;
 RECT 1.865 4.035 2.065 4.345 ;
 RECT 1.79 3.795 2.065 4.035 ;
 RECT 0.785 3.555 0.985 4.345 ;
 RECT 3.915 3.72 4.22 3.755 ;
 RECT 3.915 3.51 4.22 3.52 ;
 RECT 2.865 3.52 4.22 3.525 ;
 RECT 2.845 3.72 3.045 4.345 ;
 RECT 2.845 3.525 4.22 3.72 ;
 RECT 1.79 3.4 2.155 3.795 ;
 END
 END VDDG

 PIN SLEEP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.365 0.345 0.91 0.78 ;
 END
 ANTENNAGATEAREA 0.072 ;
 END SLEEP

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 1.355 2.96 1.495 4.01 ;
 RECT 2.295 2.96 2.435 3.95 ;
 END
 END VDD

 PIN SLEEPOUT
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.295 1.59 2.435 2.29 ;
 RECT 2.295 0.22 2.435 1.035 ;
 RECT 3.235 1.59 3.375 2.295 ;
 RECT 2.295 1.035 3.19 1.45 ;
 RECT 2.295 1.45 3.375 1.59 ;
 END
 ANTENNADIFFAREA 0.598 ;
 END SLEEPOUT

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 3.695 0.08 3.895 1.01 ;
 RECT 2.765 0.08 2.905 0.595 ;
 RECT 1.825 0.08 1.965 0.635 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 4.8 5.84 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 2.08 1.105 2.18 1.78 ;
 RECT 2.08 1.88 2.18 2.81 ;
 RECT 3.49 1.88 3.59 2.81 ;
 RECT 3.02 1.88 3.12 2.81 ;
 RECT 2.55 0.09 2.65 1.78 ;
 RECT 2.55 1.88 2.65 2.81 ;
 RECT 2.08 0.09 2.18 0.895 ;
 RECT 1.92 0.895 2.18 1.105 ;
 RECT 2.08 1.78 3.59 1.88 ;
 RECT 0.765 1.025 0.865 3.015 ;
 RECT 2.08 3.115 2.18 4.55 ;
 RECT 1.61 3.115 1.71 4.55 ;
 RECT 1.195 0.87 1.425 0.925 ;
 RECT 1.195 1.025 1.425 1.08 ;
 RECT 0.765 0.925 1.425 1.025 ;
 RECT 0.765 3.015 2.18 3.115 ;
 RECT 3.925 3.515 4.16 3.725 ;
 RECT 4.06 2.66 4.16 3.515 ;
 RECT 4.06 2.45 4.29 2.66 ;
 RECT 1.61 0.09 1.71 0.58 ;
 RECT 1.61 0.68 1.71 2.835 ;
 RECT 0.52 0.485 0.75 0.58 ;
 RECT 0.52 0.68 0.75 0.695 ;
 RECT 0.52 0.58 1.71 0.68 ;
 LAYER CO ;
 RECT 1.83 3.715 1.96 3.845 ;
 RECT 3.71 2.315 3.84 2.445 ;
 RECT 2.3 3.455 2.43 3.585 ;
 RECT 1.83 2.315 1.96 2.445 ;
 RECT 3.24 2.115 3.37 2.245 ;
 RECT 2.3 0.385 2.43 0.515 ;
 RECT 1.83 0.385 1.96 0.515 ;
 RECT 1.36 3.715 1.49 3.845 ;
 RECT 1.36 2.32 1.49 2.45 ;
 RECT 2.3 2.11 2.43 2.24 ;
 RECT 1.36 3.455 1.49 3.585 ;
 RECT 2.3 3.715 2.43 3.845 ;
 RECT 1.83 3.455 1.96 3.585 ;
 RECT 2.77 2.315 2.9 2.445 ;
 RECT 2.77 0.385 2.9 0.515 ;
 RECT 1.36 0.315 1.49 0.445 ;
 RECT 3.73 0.425 3.86 0.555 ;
 RECT 0.82 3.98 0.95 4.11 ;
 RECT 0.82 3.72 0.95 3.85 ;
 RECT 3.73 0.685 3.86 0.815 ;
 RECT 1.97 0.935 2.1 1.065 ;
 RECT 1.245 0.91 1.375 1.04 ;
 RECT 3.975 3.555 4.105 3.685 ;
 RECT 4.11 2.49 4.24 2.62 ;
 RECT 0.57 0.525 0.7 0.655 ;
 LAYER M1 ;
 RECT 1.14 0.81 1.495 0.87 ;
 RECT 1.14 1.01 1.495 1.145 ;
 RECT 1.355 0.24 1.495 0.81 ;
 RECT 1.355 1.145 1.495 2.555 ;
 RECT 1.8 0.835 2.155 0.87 ;
 RECT 1.8 1.01 2.155 1.19 ;
 RECT 1.14 0.87 2.155 1.01 ;
 RECT 2.765 2.265 2.905 2.52 ;
 RECT 1.825 2.265 1.965 2.52 ;
 RECT 3.705 2.26 3.845 2.52 ;
 RECT 4.03 2.365 4.32 2.52 ;
 RECT 1.825 2.52 4.32 2.66 ;
 END
END HEAD2X2

MACRO HEAD2X32
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 19.52 BY 5.76 ;
 PIN SLEEP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.38 0.345 0.805 0.78 ;
 END
 ANTENNAGATEAREA 0.072 ;
 END SLEEP

 PIN SLEEPOUT
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.425 0.98 2.915 1.18 ;
 RECT 2.425 0.81 2.915 0.84 ;
 RECT 11.535 0.98 11.675 2.295 ;
 RECT 11.535 0.315 11.675 0.84 ;
 RECT 16.235 0.98 16.375 2.295 ;
 RECT 16.235 0.315 16.375 0.84 ;
 RECT 14.355 0.98 14.495 2.295 ;
 RECT 14.355 0.315 14.495 0.84 ;
 RECT 12.475 0.98 12.615 2.295 ;
 RECT 12.475 0.315 12.615 0.84 ;
 RECT 3.07 0.98 3.21 2.295 ;
 RECT 3.07 0.315 3.21 0.84 ;
 RECT 2.13 0.84 16.375 0.98 ;
 RECT 2.13 0.98 2.27 2.29 ;
 RECT 2.13 0.315 2.27 0.84 ;
 RECT 4.01 0.98 4.15 2.295 ;
 RECT 4.01 0.315 4.15 0.84 ;
 RECT 4.95 0.98 5.09 2.295 ;
 RECT 4.95 0.315 5.09 0.84 ;
 RECT 5.89 0.98 6.03 2.29 ;
 RECT 5.89 0.315 6.03 0.84 ;
 RECT 7.77 0.98 7.91 2.295 ;
 RECT 7.77 0.315 7.91 0.84 ;
 RECT 8.71 0.98 8.85 2.295 ;
 RECT 8.71 0.315 8.85 0.84 ;
 RECT 6.83 0.98 6.97 2.295 ;
 RECT 6.83 0.315 6.97 0.84 ;
 RECT 10.595 0.98 10.735 2.295 ;
 RECT 10.595 0.315 10.735 0.84 ;
 RECT 13.415 0.98 13.555 2.29 ;
 RECT 13.415 0.315 13.555 0.84 ;
 RECT 9.655 0.98 9.795 2.29 ;
 RECT 9.655 0.315 9.795 0.84 ;
 RECT 15.295 0.98 15.435 2.295 ;
 RECT 15.295 0.315 15.435 0.84 ;
 END
 ANTENNADIFFAREA 9.44 ;
 END SLEEPOUT

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 19.52 2.96 ;
 RECT 1.185 2.96 1.325 4.01 ;
 RECT 10.585 2.96 10.725 3.95 ;
 RECT 16.225 2.96 16.365 3.95 ;
 RECT 15.285 2.96 15.425 3.95 ;
 RECT 9.645 2.96 9.785 3.95 ;
 RECT 12.465 2.96 12.605 3.95 ;
 RECT 14.345 2.96 14.485 3.95 ;
 RECT 11.525 2.96 11.665 3.95 ;
 RECT 13.405 2.96 13.545 3.95 ;
 RECT 2.125 2.96 2.265 3.95 ;
 RECT 3.065 2.96 3.205 3.95 ;
 RECT 4.005 2.96 4.145 3.95 ;
 RECT 4.945 2.96 5.085 3.95 ;
 RECT 6.825 2.96 6.965 3.95 ;
 RECT 5.885 2.96 6.025 3.95 ;
 RECT 8.705 2.96 8.845 3.95 ;
 RECT 7.765 2.96 7.905 3.95 ;
 END
 END VDD

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0.615 4.275 17.385 4.475 ;
 RECT 1.62 3.33 1.985 3.725 ;
 RECT 2.595 3.335 2.735 4.275 ;
 RECT 3.535 3.335 3.675 4.275 ;
 RECT 4.475 3.335 4.615 4.275 ;
 RECT 5.415 3.335 5.555 4.275 ;
 RECT 7.295 3.335 7.435 4.275 ;
 RECT 8.235 3.335 8.375 4.275 ;
 RECT 6.355 3.335 6.495 4.275 ;
 RECT 13.875 3.335 14.015 4.275 ;
 RECT 10.115 3.335 10.255 4.275 ;
 RECT 11.055 3.335 11.195 4.275 ;
 RECT 11.995 3.335 12.135 4.275 ;
 RECT 12.935 3.335 13.075 4.275 ;
 RECT 14.815 3.335 14.955 4.275 ;
 RECT 15.755 3.335 15.895 4.275 ;
 RECT 9.175 3.335 9.315 4.275 ;
 RECT 0.615 3.485 0.815 4.275 ;
 RECT 17.185 3.73 17.385 4.275 ;
 RECT 17.01 3.415 17.38 3.42 ;
 RECT 17.01 3.42 17.385 3.73 ;
 RECT 1.695 3.965 1.895 4.275 ;
 RECT 1.62 3.725 1.895 3.965 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 19.52 0.08 ;
 RECT 13.885 0.08 14.025 0.595 ;
 RECT 12.005 0.08 12.145 0.595 ;
 RECT 16.71 0.08 16.85 0.595 ;
 RECT 4.48 0.08 4.62 0.595 ;
 RECT 6.36 0.08 6.5 0.595 ;
 RECT 5.42 0.08 5.56 0.595 ;
 RECT 1.66 0.08 1.8 0.595 ;
 RECT 9.185 0.08 9.325 0.595 ;
 RECT 2.6 0.08 2.74 0.595 ;
 RECT 3.54 0.08 3.68 0.595 ;
 RECT 7.3 0.08 7.44 0.595 ;
 RECT 8.24 0.08 8.38 0.595 ;
 RECT 10.125 0.08 10.265 0.595 ;
 RECT 12.945 0.08 13.085 0.595 ;
 RECT 11.065 0.08 11.205 0.595 ;
 RECT 14.825 0.08 14.965 0.595 ;
 RECT 15.765 0.08 15.905 0.595 ;
 RECT 18.465 0.08 18.665 1.01 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 19.52 5.84 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 7.55 3.1 7.65 4.48 ;
 RECT 5.2 3.1 5.3 4.48 ;
 RECT 8.49 3.1 8.59 4.48 ;
 RECT 5.67 3.1 5.77 4.48 ;
 RECT 6.14 2.99 6.24 3 ;
 RECT 6.14 3.1 6.24 4.48 ;
 RECT 8.02 3.1 8.12 4.48 ;
 RECT 6.61 3.1 6.71 4.48 ;
 RECT 7.08 3.1 7.18 4.48 ;
 RECT 4.73 3.1 4.83 4.48 ;
 RECT 4.26 3.1 4.36 4.48 ;
 RECT 3.32 3.1 3.42 4.48 ;
 RECT 3.79 3.1 3.89 4.48 ;
 RECT 2.38 3.1 2.48 4.48 ;
 RECT 2.85 3.1 2.95 4.48 ;
 RECT 1.44 3.1 1.54 4.48 ;
 RECT 1.91 3.1 2.01 4.48 ;
 RECT 0.595 3 16.11 3.1 ;
 RECT 16.01 3.1 16.11 4.48 ;
 RECT 14.6 3.1 14.7 4.48 ;
 RECT 11.31 3.1 11.41 4.48 ;
 RECT 13.19 3.1 13.29 4.48 ;
 RECT 1.025 0.87 1.255 0.925 ;
 RECT 1.025 1.025 1.255 1.08 ;
 RECT 0.595 0.925 1.255 1.025 ;
 RECT 1.915 1.105 2.015 1.36 ;
 RECT 1.915 1.46 2.015 2.81 ;
 RECT 8.965 0.095 9.065 1.36 ;
 RECT 8.965 1.46 9.065 2.81 ;
 RECT 6.615 0.095 6.715 1.36 ;
 RECT 6.615 1.46 6.715 2.81 ;
 RECT 8.495 0.095 8.595 1.36 ;
 RECT 8.495 1.46 8.595 2.81 ;
 RECT 8.025 0.095 8.125 1.36 ;
 RECT 8.025 1.46 8.125 2.81 ;
 RECT 7.555 0.095 7.655 1.36 ;
 RECT 7.555 1.46 7.655 2.81 ;
 RECT 7.085 0.095 7.185 1.36 ;
 RECT 7.085 1.46 7.185 2.81 ;
 RECT 6.145 0.095 6.245 1.36 ;
 RECT 6.145 1.46 6.245 2.81 ;
 RECT 5.675 0.095 5.775 1.36 ;
 RECT 5.675 1.46 5.775 2.81 ;
 RECT 5.205 0.095 5.305 1.36 ;
 RECT 5.205 1.46 5.305 2.81 ;
 RECT 4.735 0.095 4.835 1.36 ;
 RECT 4.735 1.46 4.835 2.81 ;
 RECT 4.265 0.095 4.365 1.36 ;
 RECT 4.265 1.46 4.365 2.81 ;
 RECT 3.795 0.095 3.895 1.36 ;
 RECT 3.795 1.46 3.895 2.81 ;
 RECT 2.385 0.095 2.485 1.36 ;
 RECT 2.385 1.46 2.485 2.81 ;
 RECT 3.325 0.095 3.425 1.36 ;
 RECT 3.325 1.46 3.425 2.81 ;
 RECT 2.855 0.095 2.955 1.36 ;
 RECT 2.855 1.46 2.955 2.81 ;
 RECT 16.49 0.095 16.59 1.36 ;
 RECT 1.91 1.36 16.59 1.46 ;
 RECT 16.49 1.46 16.59 2.81 ;
 RECT 14.61 0.095 14.71 1.36 ;
 RECT 14.61 1.46 14.71 2.81 ;
 RECT 12.73 0.095 12.83 1.36 ;
 RECT 12.73 1.46 12.83 2.81 ;
 RECT 14.14 0.095 14.24 1.36 ;
 RECT 14.14 1.46 14.24 2.81 ;
 RECT 10.38 0.095 10.48 1.36 ;
 RECT 10.38 1.46 10.48 2.81 ;
 RECT 13.67 0.095 13.77 1.36 ;
 RECT 13.67 1.46 13.77 2.81 ;
 RECT 12.26 0.095 12.36 1.36 ;
 RECT 12.26 1.46 12.36 2.81 ;
 RECT 16.02 0.095 16.12 1.36 ;
 RECT 16.02 1.46 16.12 2.81 ;
 RECT 13.2 0.095 13.3 1.36 ;
 RECT 13.2 1.46 13.3 2.81 ;
 RECT 11.79 0.095 11.89 1.36 ;
 RECT 11.79 1.46 11.89 2.81 ;
 RECT 15.55 0.095 15.65 1.36 ;
 RECT 15.55 1.46 15.65 2.81 ;
 RECT 11.32 0.095 11.42 1.36 ;
 RECT 11.32 1.46 11.42 2.81 ;
 RECT 10.85 0.095 10.95 1.36 ;
 RECT 10.85 1.46 10.95 2.81 ;
 RECT 15.08 0.095 15.18 1.36 ;
 RECT 15.08 1.46 15.18 2.81 ;
 RECT 9.91 0.095 10.01 1.36 ;
 RECT 9.91 1.46 10.01 2.81 ;
 RECT 9.44 0.095 9.54 1.36 ;
 RECT 9.44 1.46 9.54 2.81 ;
 RECT 1.915 0.095 2.015 0.895 ;
 RECT 1.75 0.895 2.015 1.105 ;
 RECT 1.445 0.095 1.545 0.59 ;
 RECT 0.515 0.59 1.545 0.69 ;
 RECT 1.445 0.69 1.545 2.81 ;
 RECT 0.52 0.485 0.75 0.59 ;
 RECT 0.52 0.69 0.75 0.695 ;
 RECT 17.2 2.655 17.3 3.445 ;
 RECT 17.2 3.655 17.3 3.71 ;
 RECT 17.14 2.445 17.37 2.655 ;
 RECT 17.135 3.445 17.365 3.655 ;
 RECT 0.595 1.025 0.695 3 ;
 RECT 8.96 3.1 9.06 4.48 ;
 RECT 12.25 3.1 12.35 4.48 ;
 RECT 13.66 3.1 13.76 4.48 ;
 RECT 9.43 3.1 9.53 4.48 ;
 RECT 9.9 3.1 10 4.48 ;
 RECT 15.07 3.1 15.17 4.48 ;
 RECT 15.54 2.99 15.64 3 ;
 RECT 15.54 3.1 15.64 4.48 ;
 RECT 11.78 3.1 11.88 4.48 ;
 RECT 10.37 3.1 10.47 4.48 ;
 RECT 12.72 3.1 12.82 4.48 ;
 RECT 14.13 3.1 14.23 4.48 ;
 RECT 10.84 3.1 10.94 4.48 ;
 LAYER CO ;
 RECT 16.715 2.315 16.845 2.445 ;
 RECT 14.83 2.315 14.96 2.445 ;
 RECT 12.95 2.315 13.08 2.445 ;
 RECT 16.715 0.395 16.845 0.525 ;
 RECT 15.3 2.115 15.43 2.245 ;
 RECT 12.95 0.395 13.08 0.525 ;
 RECT 13.42 2.11 13.55 2.24 ;
 RECT 9.66 2.11 9.79 2.24 ;
 RECT 15.3 0.395 15.43 0.525 ;
 RECT 11.07 0.395 11.2 0.525 ;
 RECT 12.01 0.395 12.14 0.525 ;
 RECT 14.83 0.395 14.96 0.525 ;
 RECT 13.89 0.395 14.02 0.525 ;
 RECT 12.48 2.115 12.61 2.245 ;
 RECT 9.66 0.395 9.79 0.525 ;
 RECT 15.77 0.395 15.9 0.525 ;
 RECT 13.89 2.315 14.02 2.445 ;
 RECT 12.48 0.395 12.61 0.525 ;
 RECT 10.6 2.115 10.73 2.245 ;
 RECT 18.5 0.685 18.63 0.815 ;
 RECT 18.5 0.425 18.63 0.555 ;
 RECT 0.65 3.91 0.78 4.04 ;
 RECT 0.65 3.65 0.78 3.78 ;
 RECT 9.18 3.385 9.31 3.515 ;
 RECT 15.29 3.645 15.42 3.775 ;
 RECT 16.23 3.645 16.36 3.775 ;
 RECT 11.53 3.385 11.66 3.515 ;
 RECT 13.41 3.385 13.54 3.515 ;
 RECT 13.41 3.645 13.54 3.775 ;
 RECT 11.06 3.645 11.19 3.775 ;
 RECT 12.94 3.385 13.07 3.515 ;
 RECT 14.82 3.385 14.95 3.515 ;
 RECT 11.53 3.645 11.66 3.775 ;
 RECT 15.76 3.385 15.89 3.515 ;
 RECT 9.65 3.385 9.78 3.515 ;
 RECT 10.12 3.385 10.25 3.515 ;
 RECT 14.35 3.385 14.48 3.515 ;
 RECT 12 3.385 12.13 3.515 ;
 RECT 10.59 3.385 10.72 3.515 ;
 RECT 13.88 3.385 14.01 3.515 ;
 RECT 16.23 3.385 16.36 3.515 ;
 RECT 12.47 3.385 12.6 3.515 ;
 RECT 10.12 3.645 10.25 3.775 ;
 RECT 13.88 3.645 14.01 3.775 ;
 RECT 12.94 3.645 13.07 3.775 ;
 RECT 12 3.645 12.13 3.775 ;
 RECT 10.59 3.645 10.72 3.775 ;
 RECT 15.29 3.385 15.42 3.515 ;
 RECT 15.76 3.645 15.89 3.775 ;
 RECT 12.47 3.645 12.6 3.775 ;
 RECT 9.65 3.645 9.78 3.775 ;
 RECT 14.82 3.645 14.95 3.775 ;
 RECT 14.35 3.645 14.48 3.775 ;
 RECT 11.06 3.385 11.19 3.515 ;
 RECT 6.835 2.04 6.965 2.17 ;
 RECT 5.895 0.42 6.025 0.55 ;
 RECT 9.19 2.315 9.32 2.445 ;
 RECT 9.19 0.395 9.32 0.525 ;
 RECT 5.895 2.11 6.025 2.24 ;
 RECT 7.305 0.395 7.435 0.525 ;
 RECT 8.245 0.395 8.375 0.525 ;
 RECT 8.715 2.115 8.845 2.245 ;
 RECT 8.715 0.395 8.845 0.525 ;
 RECT 6.835 0.435 6.965 0.565 ;
 RECT 8.245 2.315 8.375 2.445 ;
 RECT 7.305 2.315 7.435 2.445 ;
 RECT 7.775 2.115 7.905 2.245 ;
 RECT 7.775 0.395 7.905 0.525 ;
 RECT 6.365 0.395 6.495 0.525 ;
 RECT 6.365 2.315 6.495 2.445 ;
 RECT 6.36 3.385 6.49 3.515 ;
 RECT 6.36 3.645 6.49 3.775 ;
 RECT 7.77 3.385 7.9 3.515 ;
 RECT 7.3 3.645 7.43 3.775 ;
 RECT 7.77 3.645 7.9 3.775 ;
 RECT 5.89 3.385 6.02 3.515 ;
 RECT 5.42 3.385 5.55 3.515 ;
 RECT 8.24 3.385 8.37 3.515 ;
 RECT 6.83 3.385 6.96 3.515 ;
 RECT 8.71 3.385 8.84 3.515 ;
 RECT 5.42 3.645 5.55 3.775 ;
 RECT 8.24 3.645 8.37 3.775 ;
 RECT 6.83 3.645 6.96 3.775 ;
 RECT 8.71 3.645 8.84 3.775 ;
 RECT 5.89 3.645 6.02 3.775 ;
 RECT 7.3 3.385 7.43 3.515 ;
 RECT 4.48 3.385 4.61 3.515 ;
 RECT 4.95 3.385 5.08 3.515 ;
 RECT 4.48 3.645 4.61 3.775 ;
 RECT 4.95 3.645 5.08 3.775 ;
 RECT 3.54 3.385 3.67 3.515 ;
 RECT 4.01 3.385 4.14 3.515 ;
 RECT 3.54 3.645 3.67 3.775 ;
 RECT 4.01 3.645 4.14 3.775 ;
 RECT 16.24 2.115 16.37 2.245 ;
 RECT 14.36 2.04 14.49 2.17 ;
 RECT 12.01 2.315 12.14 2.445 ;
 RECT 16.24 0.395 16.37 0.525 ;
 RECT 11.07 2.315 11.2 2.445 ;
 RECT 13.42 0.42 13.55 0.55 ;
 RECT 11.54 2.115 11.67 2.245 ;
 RECT 14.36 0.435 14.49 0.565 ;
 RECT 11.54 0.395 11.67 0.525 ;
 RECT 15.77 2.315 15.9 2.445 ;
 RECT 10.6 0.395 10.73 0.525 ;
 RECT 10.13 0.395 10.26 0.525 ;
 RECT 10.13 2.315 10.26 2.445 ;
 RECT 9.18 3.645 9.31 3.775 ;
 RECT 17.19 2.485 17.32 2.615 ;
 RECT 1.075 0.91 1.205 1.04 ;
 RECT 1.8 0.935 1.93 1.065 ;
 RECT 0.57 0.525 0.7 0.655 ;
 RECT 17.185 3.485 17.315 3.615 ;
 RECT 2.6 3.385 2.73 3.515 ;
 RECT 3.07 3.385 3.2 3.515 ;
 RECT 2.6 3.645 2.73 3.775 ;
 RECT 3.07 3.645 3.2 3.775 ;
 RECT 5.425 2.315 5.555 2.445 ;
 RECT 5.425 0.395 5.555 0.525 ;
 RECT 4.485 0.395 4.615 0.525 ;
 RECT 4.955 2.115 5.085 2.245 ;
 RECT 4.955 0.395 5.085 0.525 ;
 RECT 4.485 2.315 4.615 2.445 ;
 RECT 4.015 2.115 4.145 2.245 ;
 RECT 4.015 0.395 4.145 0.525 ;
 RECT 3.075 0.395 3.205 0.525 ;
 RECT 2.605 0.395 2.735 0.525 ;
 RECT 2.135 2.11 2.265 2.24 ;
 RECT 1.19 2.32 1.32 2.45 ;
 RECT 2.135 0.395 2.265 0.525 ;
 RECT 1.66 3.385 1.79 3.515 ;
 RECT 1.66 3.645 1.79 3.775 ;
 RECT 2.13 3.645 2.26 3.775 ;
 RECT 1.19 0.325 1.32 0.455 ;
 RECT 1.19 3.385 1.32 3.515 ;
 RECT 3.075 2.115 3.205 2.245 ;
 RECT 3.545 2.315 3.675 2.445 ;
 RECT 1.665 0.395 1.795 0.525 ;
 RECT 1.665 2.315 1.795 2.445 ;
 RECT 2.605 2.315 2.735 2.445 ;
 RECT 3.545 0.395 3.675 0.525 ;
 RECT 2.13 3.385 2.26 3.515 ;
 RECT 1.19 3.645 1.32 3.775 ;
 LAYER M1 ;
 RECT 15.765 2.26 15.905 2.52 ;
 RECT 14.825 2.26 14.965 2.52 ;
 RECT 13.885 2.265 14.025 2.52 ;
 RECT 12.945 2.26 13.085 2.52 ;
 RECT 12.005 2.26 12.145 2.52 ;
 RECT 11.065 2.26 11.205 2.52 ;
 RECT 10.125 2.265 10.265 2.52 ;
 RECT 9.185 2.26 9.325 2.52 ;
 RECT 8.24 2.26 8.38 2.52 ;
 RECT 7.3 2.26 7.44 2.52 ;
 RECT 6.36 2.265 6.5 2.52 ;
 RECT 5.42 2.26 5.56 2.52 ;
 RECT 4.48 2.26 4.62 2.52 ;
 RECT 3.54 2.26 3.68 2.52 ;
 RECT 2.6 2.265 2.74 2.52 ;
 RECT 1.66 2.265 1.8 2.52 ;
 RECT 16.71 2.26 16.85 2.52 ;
 RECT 17.09 2.34 17.435 2.52 ;
 RECT 1.655 2.52 17.435 2.66 ;
 RECT 0.97 0.81 1.325 0.87 ;
 RECT 0.97 1.01 1.325 1.145 ;
 RECT 1.185 0.24 1.325 0.81 ;
 RECT 1.185 1.145 1.325 2.555 ;
 RECT 0.97 0.87 1.985 1.01 ;
 RECT 1.63 0.835 1.985 0.87 ;
 RECT 1.63 1.01 1.985 1.19 ;
 END
END HEAD2X32

MACRO HEAD2X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.76 BY 5.76 ;
 PIN SLEEP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.33 0.345 0.91 0.835 ;
 END
 ANTENNAGATEAREA 0.074 ;
 END SLEEP

 PIN SLEEPOUT
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.295 1.59 2.435 2.3 ;
 RECT 2.295 0.235 2.435 1 ;
 RECT 3.235 1.59 3.375 2.295 ;
 RECT 3.235 0.23 3.375 1.45 ;
 RECT 2.295 1 2.885 1.45 ;
 RECT 2.295 1.45 3.375 1.59 ;
 END
 ANTENNADIFFAREA 1.18 ;
 END SLEEPOUT

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.79 3.405 2.15 3.8 ;
 RECT 1.79 3.28 2.025 3.405 ;
 RECT 1.79 3.8 2.065 3.915 ;
 RECT 0.785 4.345 4.23 4.545 ;
 RECT 1.865 3.915 2.065 4.345 ;
 RECT 3.985 3.92 4.23 4.345 ;
 RECT 0.785 3.555 0.985 4.345 ;
 RECT 2.765 3.28 2.905 4.345 ;
 END
 END VDDG

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.76 2.96 ;
 RECT 2.295 2.96 2.435 4.16 ;
 RECT 1.355 2.96 1.495 4.09 ;
 RECT 3.235 2.96 3.375 4.065 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.76 0.08 ;
 RECT 4.08 0.08 4.345 0.835 ;
 RECT 2.765 0.08 2.905 0.555 ;
 RECT 1.825 0.08 1.965 0.555 ;
 RECT 3.705 0.08 3.845 0.56 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 5.76 5.84 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 4.055 2.56 4.155 3.95 ;
 RECT 4.055 2.34 4.155 2.35 ;
 RECT 3.995 3.95 4.225 4.16 ;
 RECT 3.99 2.35 4.22 2.56 ;
 RECT 1.61 0.1 1.71 0.59 ;
 RECT 1.61 0.69 1.71 2.81 ;
 RECT 0.52 0.485 0.75 0.59 ;
 RECT 0.52 0.69 0.75 0.695 ;
 RECT 0.52 0.59 1.71 0.69 ;
 RECT 0.765 1.025 0.865 3.01 ;
 RECT 3.02 3.11 3.12 4.605 ;
 RECT 2.55 3.11 2.65 4.605 ;
 RECT 1.61 3.11 1.71 4.605 ;
 RECT 2.08 3.11 2.18 4.605 ;
 RECT 0.765 3.11 0.865 3.125 ;
 RECT 1.15 0.87 1.38 0.925 ;
 RECT 1.15 1.025 1.38 1.08 ;
 RECT 0.765 0.925 1.38 1.025 ;
 RECT 0.765 3.01 3.12 3.11 ;
 RECT 2.08 1.105 2.18 1.21 ;
 RECT 2.08 1.31 2.18 2.81 ;
 RECT 2.08 1.21 3.59 1.31 ;
 RECT 3.49 0.1 3.59 1.21 ;
 RECT 3.49 1.31 3.59 2.81 ;
 RECT 2.55 0.1 2.65 1.21 ;
 RECT 2.55 1.31 2.65 2.81 ;
 RECT 3.02 0.1 3.12 1.21 ;
 RECT 3.02 1.31 3.12 2.825 ;
 RECT 2.08 0.1 2.18 0.895 ;
 RECT 1.92 0.895 2.18 1.105 ;
 LAYER CO ;
 RECT 3.71 0.325 3.84 0.455 ;
 RECT 3.24 0.6 3.37 0.73 ;
 RECT 3.24 0.34 3.37 0.47 ;
 RECT 2.77 0.325 2.9 0.455 ;
 RECT 2.3 0.34 2.43 0.47 ;
 RECT 2.77 2 2.9 2.13 ;
 RECT 3.24 1.59 3.37 1.72 ;
 RECT 3.24 1.85 3.37 1.98 ;
 RECT 2.3 1.59 2.43 1.72 ;
 RECT 2.3 1.85 2.43 1.98 ;
 RECT 3.24 3.36 3.37 3.49 ;
 RECT 3.24 3.88 3.37 4.01 ;
 RECT 3.24 3.62 3.37 3.75 ;
 RECT 2.77 3.365 2.9 3.495 ;
 RECT 2.77 3.905 2.9 4.035 ;
 RECT 2.77 3.635 2.9 3.765 ;
 RECT 2.3 3.895 2.43 4.025 ;
 RECT 1.36 3.9 1.49 4.03 ;
 RECT 1.83 0.325 1.96 0.455 ;
 RECT 2.77 2.26 2.9 2.39 ;
 RECT 2.3 3.375 2.43 3.505 ;
 RECT 1.36 3.38 1.49 3.51 ;
 RECT 2.3 2.11 2.43 2.24 ;
 RECT 1.36 2.32 1.49 2.45 ;
 RECT 1.83 3.46 1.96 3.59 ;
 RECT 1.83 2.315 1.96 2.445 ;
 RECT 3.24 2.115 3.37 2.245 ;
 RECT 3.71 2.31 3.84 2.44 ;
 RECT 2.3 0.6 2.43 0.73 ;
 RECT 1.36 0.325 1.49 0.455 ;
 RECT 4.135 0.335 4.265 0.465 ;
 RECT 4.135 0.595 4.265 0.725 ;
 RECT 0.82 3.72 0.95 3.85 ;
 RECT 0.82 3.98 0.95 4.11 ;
 RECT 4.045 3.99 4.175 4.12 ;
 RECT 4.04 2.39 4.17 2.52 ;
 RECT 0.57 0.525 0.7 0.655 ;
 RECT 1.2 0.91 1.33 1.04 ;
 RECT 1.97 0.935 2.1 1.065 ;
 LAYER M1 ;
 RECT 2.765 1.93 2.905 2.455 ;
 RECT 1.825 2.24 1.965 2.455 ;
 RECT 1.825 2.455 4.235 2.59 ;
 RECT 1.86 2.59 4.235 2.595 ;
 RECT 3.705 2.24 3.845 2.455 ;
 RECT 3.985 2.32 4.235 2.455 ;
 RECT 1.14 0.81 1.495 0.87 ;
 RECT 1.14 1.01 1.495 1.145 ;
 RECT 1.355 0.225 1.495 0.81 ;
 RECT 1.355 1.145 1.495 2.555 ;
 RECT 1.14 0.87 2.155 1.01 ;
 RECT 1.8 0.835 2.155 0.87 ;
 RECT 1.8 1.01 2.155 1.19 ;
 END
END HEAD2X4

MACRO HEAD2X8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.68 BY 5.76 ;
 PIN SLEEP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.63 0.345 1.175 0.78 ;
 END
 ANTENNAGATEAREA 0.072 ;
 END SLEEP

 PIN SLEEPOUT
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.86 0.98 3.35 1.18 ;
 RECT 2.86 0.81 3.35 0.84 ;
 RECT 3.5 0.98 3.64 2.295 ;
 RECT 3.5 0.315 3.64 0.84 ;
 RECT 2.56 0.98 2.7 2.29 ;
 RECT 2.56 0.315 2.7 0.84 ;
 RECT 4.44 0.98 4.58 2.295 ;
 RECT 4.44 0.315 4.58 0.84 ;
 RECT 2.56 0.84 5.52 0.98 ;
 RECT 5.38 0.98 5.52 2.295 ;
 RECT 5.38 0.315 5.52 0.84 ;
 END
 ANTENNADIFFAREA 2.36 ;
 END SLEEPOUT

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.68 2.96 ;
 RECT 2.56 2.96 2.7 3.95 ;
 RECT 1.62 2.96 1.76 4.01 ;
 RECT 3.5 2.96 3.64 3.95 ;
 RECT 4.44 2.96 4.58 3.95 ;
 RECT 5.38 2.96 5.52 3.95 ;
 END
 END VDD

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 2.055 3.33 2.42 3.725 ;
 RECT 1.05 4.47 6.37 4.475 ;
 RECT 1.05 4.275 6.375 4.47 ;
 RECT 1.05 3.485 1.25 4.275 ;
 RECT 3.03 3.335 3.17 4.275 ;
 RECT 3.97 3.335 4.11 4.275 ;
 RECT 4.91 3.335 5.05 4.275 ;
 RECT 6.175 3.73 6.375 4.275 ;
 RECT 6 3.415 6.37 3.42 ;
 RECT 6 3.42 6.375 3.73 ;
 RECT 2.055 3.725 2.33 3.965 ;
 RECT 2.13 3.965 2.33 4.275 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.68 0.08 ;
 RECT 6.835 0.08 7.035 1.01 ;
 RECT 3.97 0.08 4.11 0.61 ;
 RECT 2.09 0.08 2.23 0.65 ;
 RECT 3.03 0.08 3.17 0.61 ;
 RECT 4.91 0.08 5.05 0.61 ;
 RECT 5.85 0.08 5.99 0.61 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 7.68 5.84 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 1.03 1.025 1.13 3 ;
 RECT 5.165 3.1 5.265 4.48 ;
 RECT 4.695 3.1 4.795 4.48 ;
 RECT 3.755 3.1 3.855 4.48 ;
 RECT 4.225 3.1 4.325 4.48 ;
 RECT 2.815 3.1 2.915 4.48 ;
 RECT 3.285 3.1 3.385 4.48 ;
 RECT 1.875 3.1 1.975 4.48 ;
 RECT 2.345 3.1 2.445 4.48 ;
 RECT 1.03 3.1 1.13 3.105 ;
 RECT 1.46 0.87 1.69 0.925 ;
 RECT 1.46 1.025 1.69 1.08 ;
 RECT 1.03 0.925 1.69 1.025 ;
 RECT 1.03 3 5.265 3.1 ;
 RECT 2.345 1.105 2.445 1.36 ;
 RECT 2.345 1.46 2.445 2.81 ;
 RECT 5.635 0.09 5.735 1.36 ;
 RECT 2.345 1.36 5.735 1.46 ;
 RECT 5.635 1.46 5.735 2.81 ;
 RECT 5.165 0.09 5.265 1.36 ;
 RECT 5.165 1.46 5.265 2.81 ;
 RECT 4.695 0.09 4.795 1.36 ;
 RECT 4.695 1.46 4.795 2.81 ;
 RECT 4.225 0.09 4.325 1.36 ;
 RECT 4.225 1.46 4.325 2.81 ;
 RECT 2.815 0.09 2.915 1.36 ;
 RECT 2.815 1.46 2.915 2.81 ;
 RECT 3.755 0.09 3.855 1.36 ;
 RECT 3.755 1.46 3.855 2.81 ;
 RECT 3.285 0.09 3.385 1.36 ;
 RECT 3.285 1.46 3.385 2.81 ;
 RECT 2.345 0.09 2.445 0.895 ;
 RECT 2.185 0.895 2.445 1.105 ;
 RECT 1.875 0.09 1.975 0.59 ;
 RECT 1.875 0.69 1.975 2.81 ;
 RECT 0.785 0.485 1.015 0.59 ;
 RECT 0.785 0.69 1.015 0.695 ;
 RECT 0.785 0.59 1.975 0.69 ;
 RECT 6.255 2.655 6.355 3.445 ;
 RECT 6.255 3.655 6.355 3.71 ;
 RECT 6.19 2.445 6.42 2.655 ;
 RECT 6.125 3.445 6.355 3.655 ;
 LAYER CO ;
 RECT 4.915 3.385 5.045 3.515 ;
 RECT 5.385 3.385 5.515 3.515 ;
 RECT 4.915 3.645 5.045 3.775 ;
 RECT 5.385 3.645 5.515 3.775 ;
 RECT 3.975 3.385 4.105 3.515 ;
 RECT 4.445 3.385 4.575 3.515 ;
 RECT 3.975 3.645 4.105 3.775 ;
 RECT 4.445 3.645 4.575 3.775 ;
 RECT 3.035 3.385 3.165 3.515 ;
 RECT 3.505 3.385 3.635 3.515 ;
 RECT 3.035 3.645 3.165 3.775 ;
 RECT 3.505 3.645 3.635 3.775 ;
 RECT 5.855 2.315 5.985 2.445 ;
 RECT 5.855 0.395 5.985 0.525 ;
 RECT 4.915 0.395 5.045 0.525 ;
 RECT 5.385 2.115 5.515 2.245 ;
 RECT 5.385 0.395 5.515 0.525 ;
 RECT 4.915 2.315 5.045 2.445 ;
 RECT 4.445 2.115 4.575 2.245 ;
 RECT 4.445 0.395 4.575 0.525 ;
 RECT 3.505 0.395 3.635 0.525 ;
 RECT 3.035 0.395 3.165 0.525 ;
 RECT 2.565 2.11 2.695 2.24 ;
 RECT 1.625 2.32 1.755 2.45 ;
 RECT 2.565 0.395 2.695 0.525 ;
 RECT 2.095 3.385 2.225 3.515 ;
 RECT 2.095 3.645 2.225 3.775 ;
 RECT 2.565 3.645 2.695 3.775 ;
 RECT 1.625 0.325 1.755 0.455 ;
 RECT 1.625 3.385 1.755 3.515 ;
 RECT 3.505 2.115 3.635 2.245 ;
 RECT 3.975 2.315 4.105 2.445 ;
 RECT 2.095 0.395 2.225 0.525 ;
 RECT 2.095 2.315 2.225 2.445 ;
 RECT 3.035 2.315 3.165 2.445 ;
 RECT 3.975 0.395 4.105 0.525 ;
 RECT 2.565 3.385 2.695 3.515 ;
 RECT 1.625 3.645 1.755 3.775 ;
 RECT 6.87 0.685 7 0.815 ;
 RECT 6.87 0.425 7 0.555 ;
 RECT 1.085 3.91 1.215 4.04 ;
 RECT 1.085 3.65 1.215 3.78 ;
 RECT 6.24 2.485 6.37 2.615 ;
 RECT 1.51 0.91 1.64 1.04 ;
 RECT 2.235 0.935 2.365 1.065 ;
 RECT 0.835 0.525 0.965 0.655 ;
 RECT 6.175 3.485 6.305 3.615 ;
 LAYER M1 ;
 RECT 4.91 2.26 5.05 2.52 ;
 RECT 3.97 2.26 4.11 2.52 ;
 RECT 3.03 2.265 3.17 2.52 ;
 RECT 2.09 2.265 2.23 2.52 ;
 RECT 5.85 2.26 5.99 2.52 ;
 RECT 6.19 2.34 6.535 2.52 ;
 RECT 2.09 2.52 6.535 2.66 ;
 RECT 1.405 0.81 1.76 0.87 ;
 RECT 1.405 1.01 1.76 1.145 ;
 RECT 1.62 0.24 1.76 0.81 ;
 RECT 1.62 1.145 1.76 2.555 ;
 RECT 1.405 0.87 2.42 1.01 ;
 RECT 2.065 0.835 2.42 0.87 ;
 RECT 2.065 1.01 2.42 1.19 ;
 END
END HEAD2X8

MACRO HEADX16
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.52 BY 5.76 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.52 2.96 ;
 RECT 2.04 1.885 2.18 2.8 ;
 RECT 3.015 1.855 3.155 2.8 ;
 RECT 5.94 1.9 6.08 2.8 ;
 RECT 4.965 1.855 5.105 2.8 ;
 RECT 3.99 1.855 4.13 2.8 ;
 RECT 6.935 1.855 7.075 2.8 ;
 RECT 7.91 1.855 8.05 2.8 ;
 RECT 9.86 1.9 10 2.8 ;
 RECT 8.885 1.855 9.025 2.8 ;
 END
 END VDD

 PIN SLEEP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.225 0.74 2.555 1.1 ;
 END
 ANTENNAGATEAREA 1.792 ;
 END SLEEP

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 6.44 2.09 6.58 2.485 ;
 RECT 6.22 1.715 6.795 2.09 ;
 RECT 6.22 1.695 7.555 1.715 ;
 RECT 4.47 1.7 4.61 2.485 ;
 RECT 1.63 1.7 3.635 1.715 ;
 RECT 5.485 1.495 9.505 1.5 ;
 RECT 5.445 1.7 5.585 2.485 ;
 RECT 7.415 1.715 7.555 2.485 ;
 RECT 8.39 1.695 8.53 2.485 ;
 RECT 9.365 1.695 9.505 2.485 ;
 RECT 1.63 1.695 5.615 1.7 ;
 RECT 1.63 1.715 1.77 2.475 ;
 RECT 2.52 1.715 2.66 2.485 ;
 RECT 3.495 1.715 3.635 2.485 ;
 RECT 1.63 1.5 9.505 1.695 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.52 0.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 11.52 5.84 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 9.62 1.33 9.72 2.79 ;
 RECT 9.15 1.31 9.25 2.79 ;
 RECT 8.645 1.33 8.745 2.79 ;
 RECT 8.175 1.295 8.275 2.79 ;
 RECT 7.69 1.28 9.72 1.38 ;
 RECT 7.2 1.29 7.3 2.79 ;
 RECT 6.695 1.33 6.795 2.79 ;
 RECT 7.67 1.33 7.77 2.79 ;
 RECT 6.225 1.28 7.77 1.38 ;
 RECT 6.225 1.29 6.325 2.79 ;
 RECT 5.23 1.31 5.33 2.79 ;
 RECT 4.725 1.33 4.825 2.79 ;
 RECT 4.255 1.295 4.355 2.79 ;
 RECT 5.7 1.33 5.8 2.79 ;
 RECT 3.77 1.28 6.335 1.38 ;
 RECT 3.75 1.33 3.85 2.79 ;
 RECT 3.28 1.29 3.38 2.79 ;
 RECT 2.775 1.33 2.875 2.79 ;
 RECT 2.365 1.28 3.85 1.38 ;
 RECT 2.305 0.845 2.405 2.79 ;
 RECT 2.285 0.845 2.515 1.075 ;
 LAYER CO ;
 RECT 9.865 2.27 9.995 2.4 ;
 RECT 7.915 1.97 8.045 2.1 ;
 RECT 9.37 1.97 9.5 2.1 ;
 RECT 6.94 1.935 7.07 2.065 ;
 RECT 9.865 1.97 9.995 2.1 ;
 RECT 6.94 2.27 7.07 2.4 ;
 RECT 8.395 2.27 8.525 2.4 ;
 RECT 8.89 1.935 9.02 2.065 ;
 RECT 8.89 2.27 9.02 2.4 ;
 RECT 8.89 2.27 9.02 2.4 ;
 RECT 6.445 2.27 6.575 2.4 ;
 RECT 6.94 2.27 7.07 2.4 ;
 RECT 8.395 1.97 8.525 2.1 ;
 RECT 6.445 1.97 6.575 2.1 ;
 RECT 7.42 2.27 7.55 2.4 ;
 RECT 9.37 2.27 9.5 2.4 ;
 RECT 7.915 2.27 8.045 2.4 ;
 RECT 7.915 2.27 8.045 2.4 ;
 RECT 7.42 1.97 7.55 2.1 ;
 RECT 4.475 2.27 4.605 2.4 ;
 RECT 4.97 2.27 5.1 2.4 ;
 RECT 4.475 1.97 4.605 2.1 ;
 RECT 5.45 2.27 5.58 2.4 ;
 RECT 3.995 2.27 4.125 2.4 ;
 RECT 5.945 2.27 6.075 2.4 ;
 RECT 5.45 1.97 5.58 2.1 ;
 RECT 5.945 1.97 6.075 2.1 ;
 RECT 4.97 1.935 5.1 2.065 ;
 RECT 4.97 2.27 5.1 2.4 ;
 RECT 3.5 2.27 3.63 2.4 ;
 RECT 3.995 2.27 4.125 2.4 ;
 RECT 3.5 1.97 3.63 2.1 ;
 RECT 3.995 1.97 4.125 2.1 ;
 RECT 3.02 1.935 3.15 2.065 ;
 RECT 3.02 2.27 3.15 2.4 ;
 RECT 2.525 2.27 2.655 2.4 ;
 RECT 2.525 1.97 2.655 2.1 ;
 RECT 1.635 2.015 1.765 2.145 ;
 RECT 1.635 2.275 1.765 2.405 ;
 RECT 2.335 0.895 2.465 1.025 ;
 RECT 3.02 2.27 3.15 2.4 ;
 RECT 2.045 1.935 2.175 2.065 ;
 RECT 2.045 2.27 2.175 2.4 ;
 END
END HEADX16

MACRO HEADX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 5.76 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 3.015 1.9 3.155 2.8 ;
 RECT 2.04 1.935 2.18 2.8 ;
 END
 END VDD

 PIN SLEEP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.225 0.76 2.555 1.17 ;
 END
 ANTENNAGATEAREA 0.224 ;
 END SLEEP

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.6 1.525 2.875 1.725 ;
 RECT 1.6 1.725 1.8 2.505 ;
 RECT 2.52 1.725 2.875 2.09 ;
 RECT 2.52 2.09 2.66 2.485 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 4.8 5.84 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 2.775 1.33 2.875 2.79 ;
 RECT 2.365 1.295 2.875 1.395 ;
 RECT 2.305 1.075 2.405 2.79 ;
 RECT 2.285 0.865 2.515 1.095 ;
 LAYER CO ;
 RECT 2.525 2.27 2.655 2.4 ;
 RECT 2.525 1.97 2.655 2.1 ;
 RECT 1.635 2.015 1.765 2.145 ;
 RECT 1.635 2.275 1.765 2.405 ;
 RECT 2.335 0.915 2.465 1.045 ;
 RECT 3.02 2.27 3.15 2.4 ;
 RECT 3.02 1.97 3.15 2.1 ;
 RECT 2.045 2.01 2.175 2.14 ;
 RECT 2.045 2.27 2.175 2.4 ;
 END
END HEADX2

MACRO HEADX32
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 19.52 BY 5.76 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 19.52 2.96 ;
 RECT 2.04 1.855 2.18 2.8 ;
 RECT 3.015 1.855 3.155 2.8 ;
 RECT 5.94 1.9 6.08 2.8 ;
 RECT 4.965 1.855 5.105 2.8 ;
 RECT 3.99 1.855 4.13 2.8 ;
 RECT 6.935 1.855 7.075 2.8 ;
 RECT 7.91 1.855 8.05 2.8 ;
 RECT 9.86 1.9 10 2.8 ;
 RECT 8.885 1.855 9.025 2.8 ;
 RECT 17.68 1.9 17.82 2.8 ;
 RECT 10.835 1.855 10.975 2.8 ;
 RECT 16.705 1.855 16.845 2.8 ;
 RECT 15.73 1.855 15.87 2.8 ;
 RECT 11.81 1.855 11.95 2.8 ;
 RECT 13.76 1.9 13.9 2.8 ;
 RECT 12.785 1.855 12.925 2.8 ;
 RECT 14.755 1.855 14.895 2.8 ;
 END
 END VDD

 PIN SLEEP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.29 0.815 9.585 1.105 ;
 END
 ANTENNAGATEAREA 3.584 ;
 END SLEEP

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.63 1.41 17.325 1.61 ;
 RECT 11.115 1.61 11.67 2.09 ;
 RECT 2.52 1.61 2.66 2.485 ;
 RECT 4.47 1.61 4.61 2.485 ;
 RECT 8.39 1.61 8.53 2.485 ;
 RECT 6.44 1.61 6.58 2.485 ;
 RECT 14.26 1.61 14.4 2.485 ;
 RECT 12.29 1.61 12.43 2.485 ;
 RECT 16.21 1.61 16.35 2.485 ;
 RECT 10.34 1.61 10.48 2.485 ;
 RECT 1.63 1.61 1.77 2.47 ;
 RECT 3.495 1.61 3.635 2.485 ;
 RECT 5.445 1.61 5.585 2.485 ;
 RECT 9.365 1.61 9.505 2.485 ;
 RECT 15.235 1.61 15.375 2.485 ;
 RECT 17.185 1.61 17.325 2.485 ;
 RECT 13.265 1.61 13.405 2.485 ;
 RECT 7.415 1.61 7.555 2.485 ;
 RECT 11.315 2.09 11.455 2.485 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 19.52 0.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 19.52 5.84 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 17.44 1.33 17.54 2.79 ;
 RECT 16.97 1.31 17.07 2.79 ;
 RECT 15.995 1.295 16.095 2.79 ;
 RECT 16.465 1.33 16.565 2.79 ;
 RECT 15.51 1.28 17.54 1.38 ;
 RECT 14.515 1.33 14.615 2.79 ;
 RECT 15.49 1.33 15.59 2.79 ;
 RECT 15.02 1.29 15.12 2.79 ;
 RECT 2.775 1.33 2.875 2.79 ;
 RECT 2.305 1.29 2.405 2.79 ;
 RECT 3.28 1.29 3.38 2.79 ;
 RECT 14.045 1.28 15.59 1.38 ;
 RECT 13.52 1.33 13.62 2.79 ;
 RECT 13.05 1.31 13.15 2.79 ;
 RECT 14.045 1.29 14.145 2.79 ;
 RECT 12.545 1.33 12.645 2.79 ;
 RECT 12.075 1.295 12.175 2.79 ;
 RECT 2.305 1.28 3.85 1.38 ;
 RECT 5.23 1.31 5.33 2.79 ;
 RECT 4.725 1.33 4.825 2.79 ;
 RECT 4.255 1.295 4.355 2.79 ;
 RECT 5.7 1.33 5.8 2.79 ;
 RECT 3.75 1.33 3.85 2.79 ;
 RECT 11.59 1.28 14.155 1.38 ;
 RECT 10.125 1.29 10.225 2.79 ;
 RECT 11.1 1.29 11.2 2.79 ;
 RECT 10.595 1.33 10.695 2.79 ;
 RECT 11.57 1.33 11.67 2.79 ;
 RECT 3.77 1.28 6.335 1.38 ;
 RECT 7.2 1.29 7.3 2.79 ;
 RECT 6.695 1.33 6.795 2.79 ;
 RECT 6.225 1.29 6.325 2.79 ;
 RECT 9.685 1.28 11.67 1.38 ;
 RECT 6.225 1.28 7.77 1.38 ;
 RECT 9.62 1.33 9.72 2.79 ;
 RECT 9.15 1.31 9.25 2.79 ;
 RECT 8.645 1.33 8.745 2.79 ;
 RECT 8.175 1.295 8.275 2.79 ;
 RECT 7.67 1.33 7.77 2.79 ;
 RECT 7.69 1.28 9.72 1.38 ;
 RECT 9.325 1.09 9.555 1.33 ;
 RECT 9.325 0.86 9.555 1.09 ;
 LAYER CO ;
 RECT 13.765 2.27 13.895 2.4 ;
 RECT 11.815 1.97 11.945 2.1 ;
 RECT 13.27 1.97 13.4 2.1 ;
 RECT 10.84 1.935 10.97 2.065 ;
 RECT 16.71 2.27 16.84 2.4 ;
 RECT 15.735 2.27 15.865 2.4 ;
 RECT 17.19 1.97 17.32 2.1 ;
 RECT 14.265 2.27 14.395 2.4 ;
 RECT 15.24 1.97 15.37 2.1 ;
 RECT 13.765 1.97 13.895 2.1 ;
 RECT 10.84 2.27 10.97 2.4 ;
 RECT 14.76 1.935 14.89 2.065 ;
 RECT 14.76 2.27 14.89 2.4 ;
 RECT 12.295 2.27 12.425 2.4 ;
 RECT 12.79 1.935 12.92 2.065 ;
 RECT 17.685 1.97 17.815 2.1 ;
 RECT 16.215 1.97 16.345 2.1 ;
 RECT 12.79 2.27 12.92 2.4 ;
 RECT 12.79 2.27 12.92 2.4 ;
 RECT 10.345 2.27 10.475 2.4 ;
 RECT 10.84 2.27 10.97 2.4 ;
 RECT 14.76 2.27 14.89 2.4 ;
 RECT 14.265 1.97 14.395 2.1 ;
 RECT 12.295 1.97 12.425 2.1 ;
 RECT 10.345 1.97 10.475 2.1 ;
 RECT 16.215 2.27 16.345 2.4 ;
 RECT 11.32 2.27 11.45 2.4 ;
 RECT 9.865 2.27 9.995 2.4 ;
 RECT 16.71 1.935 16.84 2.065 ;
 RECT 15.24 2.27 15.37 2.4 ;
 RECT 13.27 2.27 13.4 2.4 ;
 RECT 11.815 2.27 11.945 2.4 ;
 RECT 17.685 2.27 17.815 2.4 ;
 RECT 17.19 2.27 17.32 2.4 ;
 RECT 11.815 2.27 11.945 2.4 ;
 RECT 11.32 1.97 11.45 2.1 ;
 RECT 15.735 1.97 15.865 2.1 ;
 RECT 16.71 2.27 16.84 2.4 ;
 RECT 15.735 2.27 15.865 2.4 ;
 RECT 9.865 2.27 9.995 2.4 ;
 RECT 7.915 1.97 8.045 2.1 ;
 RECT 9.37 1.97 9.5 2.1 ;
 RECT 6.94 1.935 7.07 2.065 ;
 RECT 9.865 1.97 9.995 2.1 ;
 RECT 6.94 2.27 7.07 2.4 ;
 RECT 8.395 2.27 8.525 2.4 ;
 RECT 8.89 1.935 9.02 2.065 ;
 RECT 8.89 2.27 9.02 2.4 ;
 RECT 8.89 2.27 9.02 2.4 ;
 RECT 6.445 2.27 6.575 2.4 ;
 RECT 6.94 2.27 7.07 2.4 ;
 RECT 8.395 1.97 8.525 2.1 ;
 RECT 6.445 1.97 6.575 2.1 ;
 RECT 7.42 2.27 7.55 2.4 ;
 RECT 9.37 2.27 9.5 2.4 ;
 RECT 7.915 2.27 8.045 2.4 ;
 RECT 7.915 2.27 8.045 2.4 ;
 RECT 7.42 1.97 7.55 2.1 ;
 RECT 4.475 2.27 4.605 2.4 ;
 RECT 4.97 2.27 5.1 2.4 ;
 RECT 4.475 1.97 4.605 2.1 ;
 RECT 5.45 2.27 5.58 2.4 ;
 RECT 3.995 2.27 4.125 2.4 ;
 RECT 5.945 2.27 6.075 2.4 ;
 RECT 5.45 1.97 5.58 2.1 ;
 RECT 5.945 1.97 6.075 2.1 ;
 RECT 4.97 1.935 5.1 2.065 ;
 RECT 4.97 2.27 5.1 2.4 ;
 RECT 3.5 2.27 3.63 2.4 ;
 RECT 3.995 2.27 4.125 2.4 ;
 RECT 3.5 1.97 3.63 2.1 ;
 RECT 3.995 1.97 4.125 2.1 ;
 RECT 3.02 1.935 3.15 2.065 ;
 RECT 3.02 2.27 3.15 2.4 ;
 RECT 2.525 2.27 2.655 2.4 ;
 RECT 2.525 1.97 2.655 2.1 ;
 RECT 1.635 2.015 1.765 2.145 ;
 RECT 1.635 2.275 1.765 2.405 ;
 RECT 9.375 0.91 9.505 1.04 ;
 RECT 3.02 2.27 3.15 2.4 ;
 RECT 2.045 1.935 2.175 2.065 ;
 RECT 2.045 2.27 2.175 2.4 ;
 END
END HEADX32

MACRO HEADX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.76 BY 5.76 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.76 2.96 ;
 RECT 2.04 2.005 2.18 2.8 ;
 RECT 3.99 1.9 4.13 2.8 ;
 RECT 3.015 2.175 3.155 2.8 ;
 END
 END VDD

 PIN SLEEP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.225 0.765 2.555 1.125 ;
 END
 ANTENNAGATEAREA 0.448 ;
 END SLEEP

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.6 1.745 1.8 2.505 ;
 RECT 2.49 1.745 2.875 2.09 ;
 RECT 2.49 2.09 2.69 2.515 ;
 RECT 3.465 1.745 3.665 2.515 ;
 RECT 1.6 1.545 3.665 1.745 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.76 0.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 5.76 5.84 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 3.75 1.33 3.85 2.79 ;
 RECT 3.28 1.305 3.38 2.79 ;
 RECT 2.775 1.33 2.875 2.79 ;
 RECT 2.365 1.295 3.85 1.395 ;
 RECT 2.305 1.06 2.405 2.79 ;
 RECT 2.285 0.87 2.515 1.1 ;
 LAYER CO ;
 RECT 3.5 2.27 3.63 2.4 ;
 RECT 3.995 2.27 4.125 2.4 ;
 RECT 3.5 1.97 3.63 2.1 ;
 RECT 3.995 1.97 4.125 2.1 ;
 RECT 3.02 2.27 3.15 2.4 ;
 RECT 2.525 2.27 2.655 2.4 ;
 RECT 2.525 1.97 2.655 2.1 ;
 RECT 1.635 2.015 1.765 2.145 ;
 RECT 1.635 2.275 1.765 2.405 ;
 RECT 2.335 0.92 2.465 1.05 ;
 RECT 3.02 2.27 3.15 2.4 ;
 RECT 2.045 2.27 2.175 2.4 ;
 END
END HEADX4

MACRO HEADX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.68 BY 5.76 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.68 2.96 ;
 RECT 2.04 1.93 2.18 2.8 ;
 RECT 3.99 1.945 4.13 2.8 ;
 RECT 3.015 2.105 3.155 2.8 ;
 RECT 5.94 1.9 6.08 2.8 ;
 RECT 4.965 1.885 5.105 2.8 ;
 END
 END VDD

 PIN SLEEP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.225 0.75 2.555 1.11 ;
 END
 ANTENNAGATEAREA 0.896 ;
 END SLEEP

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.6 1.745 1.8 2.505 ;
 RECT 2.49 1.745 2.875 2.09 ;
 RECT 2.49 2.09 2.69 2.515 ;
 RECT 4.44 1.745 4.64 2.515 ;
 RECT 1.6 1.545 5.615 1.745 ;
 RECT 3.465 1.745 3.665 2.515 ;
 RECT 5.415 1.745 5.615 2.515 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.68 0.08 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 7.68 5.84 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 5.23 1.31 5.33 2.79 ;
 RECT 4.725 1.33 4.825 2.79 ;
 RECT 4.255 1.295 4.355 2.79 ;
 RECT 5.7 1.33 5.8 2.79 ;
 RECT 3.77 1.295 5.8 1.395 ;
 RECT 3.75 1.33 3.85 2.79 ;
 RECT 3.28 1.29 3.38 2.79 ;
 RECT 2.775 1.33 2.875 2.79 ;
 RECT 2.365 1.295 3.85 1.395 ;
 RECT 2.305 1.03 2.405 2.79 ;
 RECT 2.285 0.855 2.515 1.085 ;
 LAYER CO ;
 RECT 4.475 2.27 4.605 2.4 ;
 RECT 4.97 2.27 5.1 2.4 ;
 RECT 4.475 1.97 4.605 2.1 ;
 RECT 5.45 2.27 5.58 2.4 ;
 RECT 3.995 2.27 4.125 2.4 ;
 RECT 5.945 2.27 6.075 2.4 ;
 RECT 5.45 1.97 5.58 2.1 ;
 RECT 5.945 1.97 6.075 2.1 ;
 RECT 4.97 1.95 5.1 2.08 ;
 RECT 4.97 2.27 5.1 2.4 ;
 RECT 3.5 2.27 3.63 2.4 ;
 RECT 3.995 2.27 4.125 2.4 ;
 RECT 3.5 1.97 3.63 2.1 ;
 RECT 3.995 2.01 4.125 2.14 ;
 RECT 3.02 2.27 3.15 2.4 ;
 RECT 2.525 2.27 2.655 2.4 ;
 RECT 2.525 1.97 2.655 2.1 ;
 RECT 1.635 2.015 1.765 2.145 ;
 RECT 1.635 2.275 1.765 2.405 ;
 RECT 2.335 0.905 2.465 1.035 ;
 RECT 3.02 2.27 3.15 2.4 ;
 RECT 2.045 2.27 2.175 2.4 ;
 END
END HEADX8

MACRO NMT1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN G
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.985 0.82 1.385 1.11 ;
 END
 ANTENNAGATEAREA 0.048 ;
 END G

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.095 0.83 0.47 1.11 ;
 RECT 0.095 0.305 0.635 0.445 ;
 RECT 0.095 0.445 0.235 0.83 ;
 END
 ANTENNADIFFAREA 0.144 ;
 END D

 PIN S
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.875 0.305 1.655 0.445 ;
 RECT 1.295 0.445 1.655 0.625 ;
 RECT 1.295 0.235 1.655 0.305 ;
 END
 ANTENNADIFFAREA 0.144 ;
 END S

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 RECT 2 0.08 2.16 0.755 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.705 0.09 0.805 0.92 ;
 RECT 0.705 0.92 1.15 1.02 ;
 RECT 0.985 0.84 1.215 1.07 ;
 LAYER CO ;
 RECT 1.035 0.89 1.165 1.02 ;
 RECT 2.015 0.31 2.145 0.44 ;
 RECT 2.015 0.575 2.145 0.705 ;
 RECT 0.925 0.31 1.055 0.44 ;
 RECT 0.455 0.31 0.585 0.44 ;
 END
END NMT1

MACRO NMT2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN G
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.945 1.77 1.36 2.11 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END G

 PIN S
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.17 0.83 0.47 1.08 ;
 RECT 0.265 1.22 1.53 1.36 ;
 RECT 0.265 0.315 0.625 0.455 ;
 RECT 0.265 1.08 0.405 1.22 ;
 RECT 0.265 0.455 0.405 0.83 ;
 RECT 1.39 0.26 1.53 1.22 ;
 END
 ANTENNADIFFAREA 0.288 ;
 END S

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.92 0.53 1.06 0.82 ;
 RECT 0.655 0.82 1.06 1.08 ;
 END
 ANTENNADIFFAREA 0.178 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 RECT 2 0.08 2.16 0.755 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.705 0.09 0.805 0.92 ;
 RECT 0.705 0.92 1.275 1.02 ;
 RECT 1.175 0.09 1.275 1.005 ;
 RECT 1.1 0.97 1.2 1.86 ;
 RECT 1.025 1.79 1.255 2.02 ;
 LAYER CO ;
 RECT 1.075 1.84 1.205 1.97 ;
 RECT 2.015 0.31 2.145 0.44 ;
 RECT 2.015 0.575 2.145 0.705 ;
 RECT 1.395 0.31 1.525 0.44 ;
 RECT 0.925 0.58 1.055 0.71 ;
 RECT 0.445 0.32 0.575 0.45 ;
 END
END NMT2

MACRO NMT3
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 2.88 ;
 PIN G
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.12 1.775 1.43 2.1 ;
 END
 ANTENNAGATEAREA 0.192 ;
 END G

 PIN S
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.33 1.22 2.59 1.36 ;
 RECT 0.33 1.13 0.635 1.22 ;
 RECT 0.55 0.225 1.64 0.365 ;
 RECT 0.33 1.36 0.635 1.43 ;
 RECT 2.45 0.26 2.59 1.22 ;
 RECT 0.375 0.585 0.69 0.725 ;
 RECT 1.5 0.365 1.64 0.49 ;
 RECT 0.55 0.365 0.69 0.585 ;
 RECT 0.375 0.725 0.515 1.13 ;
 END
 ANTENNADIFFAREA 0.471 ;
 END S

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.955 0.51 1.34 0.77 ;
 RECT 1.97 0.53 2.11 0.94 ;
 RECT 1.03 0.94 2.11 1.08 ;
 RECT 1.03 0.77 1.17 0.94 ;
 END
 ANTENNADIFFAREA 0.358 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 3.28 0.08 3.44 0.755 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 2.23 0.09 2.33 1.02 ;
 RECT 1.755 0.09 1.855 1.005 ;
 RECT 0.815 0.09 0.915 0.92 ;
 RECT 0.815 0.92 2.33 1.02 ;
 RECT 1.285 0.09 1.385 1.005 ;
 RECT 1.21 0.97 1.31 1.86 ;
 RECT 1.135 1.79 1.365 2.02 ;
 LAYER CO ;
 RECT 1.185 1.84 1.315 1.97 ;
 RECT 3.295 0.31 3.425 0.44 ;
 RECT 3.295 0.575 3.425 0.705 ;
 RECT 2.455 0.31 2.585 0.44 ;
 RECT 1.975 0.58 2.105 0.71 ;
 RECT 1.505 0.31 1.635 0.44 ;
 RECT 1.035 0.58 1.165 0.71 ;
 RECT 0.555 0.32 0.685 0.45 ;
 END
END NMT3

MACRO PMT1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.24 BY 2.88 ;
 PIN G
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.345 0.73 0.635 1.105 ;
 END
 ANTENNAGATEAREA 0.112 ;
 END G

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.985 0.815 1.27 1.1 ;
 RECT 0.985 1.1 1.125 2.615 ;
 END
 ANTENNADIFFAREA 0.347 ;
 END D

 PIN S
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.505 1.745 0.645 2.615 ;
 RECT 0.075 1.535 0.645 1.745 ;
 RECT 0.075 1.455 0.64 1.535 ;
 END
 ANTENNADIFFAREA 0.336 ;
 END S

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.24 2.96 ;
 RECT 1.69 1.865 1.83 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.24 0.08 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.76 1.305 0.86 2.785 ;
 RECT 0.345 1.235 0.86 1.335 ;
 RECT 0.345 0.905 0.445 1.3 ;
 RECT 0.345 0.825 0.575 1.055 ;
 LAYER CO ;
 RECT 0.395 0.875 0.525 1.005 ;
 RECT 1.695 1.915 1.825 2.045 ;
 RECT 1.695 2.175 1.825 2.305 ;
 RECT 0.51 1.89 0.64 2.02 ;
 RECT 0.51 1.62 0.64 1.75 ;
 RECT 0.99 1.635 1.12 1.765 ;
 RECT 0.99 1.895 1.12 2.025 ;
 RECT 0.99 2.165 1.12 2.295 ;
 RECT 0.99 2.435 1.12 2.565 ;
 RECT 0.51 2.16 0.64 2.29 ;
 RECT 0.51 2.435 0.64 2.565 ;
 END
END PMT1

MACRO DFFNASX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.84 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.84 2.96 ;
 RECT 1.98 2.62 2.23 2.8 ;
 RECT 4.495 2.635 4.755 2.8 ;
 RECT 1.5 2.05 1.64 2.8 ;
 RECT 0.54 1.76 0.68 2.8 ;
 RECT 8.26 2.055 8.4 2.8 ;
 RECT 9.38 1.48 9.52 2.8 ;
 RECT 5.485 2.38 5.625 2.8 ;
 RECT 10.415 1.48 10.555 2.8 ;
 RECT 11.36 1.48 11.5 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.84 0.08 ;
 RECT 1.5 0.08 1.64 1.075 ;
 RECT 10.285 0.08 10.565 0.245 ;
 RECT 2.075 0.08 2.305 0.385 ;
 RECT 4.465 0.08 4.605 0.38 ;
 RECT 9.315 0.08 9.455 0.655 ;
 RECT 0.54 0.08 0.68 0.795 ;
 RECT 7.775 0.08 7.915 1.07 ;
 RECT 11.355 0.08 11.495 0.85 ;
 END
 END VSS

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.03 0.44 7.365 0.785 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END SETB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.135 1.78 1.77 1.88 ;
 RECT 1.75 1.505 2.025 1.555 ;
 RECT 1.75 1.555 2.03 1.615 ;
 RECT 1.135 1.615 2.03 1.78 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 0.29 1.325 0.6 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.88 2.11 10.215 2.36 ;
 RECT 9.88 2.36 10.02 2.51 ;
 RECT 9.88 0.675 10.02 2.11 ;
 END
 ANTENNADIFFAREA 0.714 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.885 2.11 11.175 2.36 ;
 RECT 10.885 2.36 11.025 2.51 ;
 RECT 10.885 0.58 11.025 2.11 ;
 END
 ANTENNADIFFAREA 0.622 ;
 END Q

 OBS
 LAYER PO ;
 RECT 2.285 1.675 2.635 1.69 ;
 RECT 4.25 0.285 4.35 1.24 ;
 RECT 2.6 0.185 4.35 0.285 ;
 RECT 2.535 1.355 2.635 1.44 ;
 RECT 2.6 0.285 2.7 1.255 ;
 RECT 3.42 1.675 3.52 2.5 ;
 RECT 2.535 1.69 2.635 2.275 ;
 RECT 2.535 1.255 2.7 1.355 ;
 RECT 5.155 0.575 5.905 0.675 ;
 RECT 5.805 0.675 5.905 1.35 ;
 RECT 7.56 0.265 7.66 1.32 ;
 RECT 5.805 0.265 5.905 0.575 ;
 RECT 5.155 0.455 5.385 0.575 ;
 RECT 5.155 0.675 5.385 0.685 ;
 RECT 6.25 1.545 6.35 2.435 ;
 RECT 5.805 0.165 7.66 0.265 ;
 RECT 5.805 1.35 6.095 1.445 ;
 RECT 5.805 1.445 6.35 1.45 ;
 RECT 5.995 1.45 6.35 1.545 ;
 RECT 11.14 0.14 11.24 1.135 ;
 RECT 11.14 1.235 11.24 2.79 ;
 RECT 10.56 1.07 10.77 1.135 ;
 RECT 10.56 1.235 10.77 1.305 ;
 RECT 10.56 1.135 11.24 1.235 ;
 RECT 10.67 0.14 10.77 1.07 ;
 RECT 10.67 1.305 10.77 2.79 ;
 RECT 8.03 1.53 8.615 1.63 ;
 RECT 8.39 1.63 8.615 1.94 ;
 RECT 8.03 0.65 8.13 1.53 ;
 RECT 8.515 1.94 8.615 2.56 ;
 RECT 4.575 0.625 4.675 1.58 ;
 RECT 4.705 1.82 4.805 2.455 ;
 RECT 4.575 1.58 4.815 1.82 ;
 RECT 3.915 1.43 4.015 1.475 ;
 RECT 3.915 1.71 4.015 2.505 ;
 RECT 3.935 0.65 4.035 1.33 ;
 RECT 3.915 1.33 4.035 1.43 ;
 RECT 3.785 1.475 4.015 1.71 ;
 RECT 4.22 1.795 4.32 2.685 ;
 RECT 2.84 2.08 3.05 2.685 ;
 RECT 2.84 2.685 4.32 2.785 ;
 RECT 3.465 0.47 3.75 0.705 ;
 RECT 3.465 0.705 3.565 1.145 ;
 RECT 2.88 1.145 3.565 1.395 ;
 RECT 1.76 0.675 1.86 1.5 ;
 RECT 1.76 1.5 2.03 1.74 ;
 RECT 1.76 1.74 1.86 2.39 ;
 RECT 5.525 1.095 5.625 1.64 ;
 RECT 5.525 1.64 5.84 1.87 ;
 RECT 5.355 0.865 5.625 1.095 ;
 RECT 6.745 0.645 6.845 1.24 ;
 RECT 6.745 1.24 6.99 1.45 ;
 RECT 6.745 1.45 6.845 2.37 ;
 RECT 6.275 0.685 6.375 1.23 ;
 RECT 6.2 0.455 6.43 0.685 ;
 RECT 9.065 1.18 10.295 1.28 ;
 RECT 9.065 1.28 9.275 1.415 ;
 RECT 9.645 0.145 9.745 1.18 ;
 RECT 9.645 1.28 9.745 2.79 ;
 RECT 10.195 1.28 10.295 2.79 ;
 RECT 10.135 0.14 10.235 1.18 ;
 RECT 1.08 0.33 1.385 0.57 ;
 RECT 1.285 0.57 1.385 2.485 ;
 RECT 5.195 1.375 5.295 2.69 ;
 RECT 4.875 1.275 5.295 1.375 ;
 RECT 5.195 2.69 7.32 2.79 ;
 RECT 7.22 0.72 7.32 2.69 ;
 RECT 7.085 0.5 7.32 0.72 ;
 RECT 7.085 0.49 7.315 0.5 ;
 RECT 4.875 0.635 4.975 1.275 ;
 RECT 7.83 2.47 8.145 2.71 ;
 RECT 8.045 1.84 8.145 2.47 ;
 RECT 2.285 1.575 3.52 1.675 ;
 RECT 2.285 1.44 2.635 1.575 ;
 LAYER CO ;
 RECT 3.835 1.525 3.965 1.655 ;
 RECT 4.545 2.64 4.675 2.77 ;
 RECT 10.6 1.12 10.73 1.25 ;
 RECT 11.36 0.65 11.49 0.78 ;
 RECT 11.365 1.79 11.495 1.92 ;
 RECT 11.365 2.05 11.495 2.18 ;
 RECT 7.895 2.525 8.025 2.655 ;
 RECT 11.365 2.31 11.495 2.44 ;
 RECT 11.365 1.53 11.495 1.66 ;
 RECT 10.89 2.05 11.02 2.18 ;
 RECT 10.89 1.79 11.02 1.92 ;
 RECT 5.66 1.69 5.79 1.82 ;
 RECT 5.42 0.915 5.55 1.045 ;
 RECT 5.205 0.505 5.335 0.635 ;
 RECT 6.495 1.9 6.625 2.03 ;
 RECT 6.025 0.87 6.155 1 ;
 RECT 6.25 0.505 6.38 0.635 ;
 RECT 6.805 1.28 6.935 1.41 ;
 RECT 9.105 1.23 9.235 1.36 ;
 RECT 10.42 1.53 10.55 1.66 ;
 RECT 10.42 1.79 10.55 1.92 ;
 RECT 10.42 2.05 10.55 2.18 ;
 RECT 10.42 2.31 10.55 2.44 ;
 RECT 9.385 1.53 9.515 1.66 ;
 RECT 9.385 1.79 9.515 1.92 ;
 RECT 9.385 2.05 9.515 2.18 ;
 RECT 9.385 2.31 9.515 2.44 ;
 RECT 2.82 0.905 2.95 1.035 ;
 RECT 5.095 0.88 5.225 1.01 ;
 RECT 4.47 0.2 4.6 0.33 ;
 RECT 2.755 1.81 2.885 1.94 ;
 RECT 3.57 0.525 3.7 0.655 ;
 RECT 7.125 0.54 7.255 0.67 ;
 RECT 0.545 2.105 0.675 2.235 ;
 RECT 2.11 0.895 2.24 1.025 ;
 RECT 9.885 0.725 10.015 0.855 ;
 RECT 1.13 0.385 1.26 0.515 ;
 RECT 7.78 0.87 7.91 1 ;
 RECT 0.545 1.845 0.675 1.975 ;
 RECT 1.505 2.12 1.635 2.25 ;
 RECT 2.355 1.495 2.485 1.625 ;
 RECT 2.05 2.63 2.18 2.76 ;
 RECT 3.665 2.07 3.795 2.2 ;
 RECT 3.685 0.88 3.815 1.01 ;
 RECT 3.17 2.105 3.3 2.235 ;
 RECT 3.215 0.88 3.345 1.01 ;
 RECT 6 1.815 6.13 1.945 ;
 RECT 5.49 2.44 5.62 2.57 ;
 RECT 6.495 0.87 6.625 1 ;
 RECT 7.445 1.965 7.575 2.095 ;
 RECT 6.965 1.965 7.095 2.095 ;
 RECT 8.25 0.87 8.38 1 ;
 RECT 8.265 2.115 8.395 2.245 ;
 RECT 7.795 2.11 7.925 2.24 ;
 RECT 8.825 2.13 8.955 2.26 ;
 RECT 8.44 1.76 8.57 1.89 ;
 RECT 4.645 1.63 4.775 1.76 ;
 RECT 4.93 2.015 5.06 2.145 ;
 RECT 2.125 0.25 2.255 0.38 ;
 RECT 2.88 2.135 3.01 2.265 ;
 RECT 2.95 1.2 3.08 1.33 ;
 RECT 0.545 0.61 0.675 0.74 ;
 RECT 0.545 0.35 0.675 0.48 ;
 RECT 1.505 0.895 1.635 1.025 ;
 RECT 1.86 1.555 1.99 1.685 ;
 RECT 1.035 0.895 1.165 1.025 ;
 RECT 1.035 2.11 1.165 2.24 ;
 RECT 0.545 2.365 0.675 2.495 ;
 RECT 1.98 2.015 2.11 2.145 ;
 RECT 10.89 1.53 11.02 1.66 ;
 RECT 10.89 2.31 11.02 2.44 ;
 RECT 10.89 0.65 11.02 0.78 ;
 RECT 10.355 0.11 10.485 0.24 ;
 RECT 9.32 0.475 9.45 0.605 ;
 RECT 9.885 1.79 10.015 1.92 ;
 RECT 9.885 1.53 10.015 1.66 ;
 RECT 9.885 2.05 10.015 2.18 ;
 RECT 9.885 2.31 10.015 2.44 ;
 LAYER M1 ;
 RECT 4.925 1.04 5.6 1.05 ;
 RECT 4.36 0.91 5.6 1.04 ;
 RECT 4.36 0.9 5.23 0.91 ;
 RECT 4.925 1.08 5.065 2.2 ;
 RECT 4.925 1.05 5.23 1.08 ;
 RECT 3.785 1.52 4.5 1.66 ;
 RECT 5.09 0.81 5.23 0.9 ;
 RECT 4.36 1.04 4.5 1.52 ;
 RECT 3.5 0.52 5.41 0.66 ;
 RECT 5.125 0.47 5.41 0.52 ;
 RECT 5.205 1.36 5.345 2.1 ;
 RECT 5.205 2.24 5.345 2.355 ;
 RECT 4.13 2.355 5.345 2.495 ;
 RECT 2.465 2.515 4.27 2.655 ;
 RECT 2.105 0.845 2.245 1.125 ;
 RECT 2.35 2.15 2.49 2.34 ;
 RECT 4.13 2.495 4.27 2.515 ;
 RECT 2.465 2.48 2.605 2.515 ;
 RECT 2.35 2.34 2.605 2.48 ;
 RECT 2.105 1.125 2.49 1.265 ;
 RECT 2.35 1.265 2.49 2.01 ;
 RECT 1.91 2.01 2.49 2.15 ;
 RECT 6.61 2.32 6.75 2.52 ;
 RECT 5.74 0.5 6.455 0.64 ;
 RECT 5.74 0.64 5.88 1.22 ;
 RECT 5.205 2.1 6.105 2.18 ;
 RECT 5.205 2.18 6.75 2.24 ;
 RECT 5.965 2.24 6.75 2.32 ;
 RECT 5.205 1.22 5.88 1.36 ;
 RECT 6.61 2.52 8.105 2.66 ;
 RECT 2.815 1.41 3.015 1.725 ;
 RECT 2.815 0.83 2.955 1.15 ;
 RECT 2.815 1.15 3.085 1.41 ;
 RECT 2.75 1.725 3.015 2.335 ;
 RECT 3.505 1.805 4.78 1.945 ;
 RECT 3.505 1.945 3.87 1.96 ;
 RECT 3.505 1.22 3.82 1.36 ;
 RECT 3.68 0.805 3.82 1.22 ;
 RECT 3.59 1.96 3.87 2.215 ;
 RECT 3.505 1.36 3.645 1.805 ;
 RECT 4.64 1.56 4.78 1.805 ;
 RECT 6.96 2.1 7.145 2.24 ;
 RECT 7.79 2.03 7.93 2.24 ;
 RECT 6.915 1.96 7.145 2.1 ;
 RECT 6.96 2.24 7.93 2.38 ;
 RECT 6.49 1.815 6.7 1.895 ;
 RECT 6.49 0.805 6.63 1.675 ;
 RECT 7.395 1.815 7.625 2.1 ;
 RECT 6.42 1.895 6.7 2.035 ;
 RECT 6.49 1.675 8.68 1.815 ;
 RECT 9.1 1.18 9.24 2.505 ;
 RECT 8.38 1.815 8.68 1.915 ;
 RECT 8.54 1.915 8.68 2.505 ;
 RECT 8.54 2.505 9.24 2.645 ;
 RECT 5.65 1.685 6.16 1.81 ;
 RECT 5.65 1.81 6.2 1.825 ;
 RECT 6.02 0.78 6.16 1.685 ;
 RECT 5.65 1.615 5.79 1.685 ;
 RECT 5.65 1.825 5.79 1.895 ;
 RECT 5.93 1.825 6.2 1.95 ;
 RECT 8.82 1.005 8.96 1.395 ;
 RECT 6.8 1.395 8.96 1.535 ;
 RECT 8.82 1.535 8.96 2.32 ;
 RECT 6.8 1.21 6.94 1.395 ;
 RECT 9.595 0.535 9.735 0.865 ;
 RECT 9.595 0.38 9.735 0.395 ;
 RECT 8.2 0.865 9.735 1.005 ;
 RECT 9.595 0.395 10.735 0.535 ;
 RECT 10.595 0.535 10.735 1.315 ;
 RECT 0.82 1.355 0.96 2.105 ;
 RECT 0.82 1.03 0.96 1.215 ;
 RECT 0.82 2.105 1.235 2.245 ;
 RECT 0.82 0.89 1.24 1.03 ;
 RECT 1.78 0.665 1.92 1.215 ;
 RECT 3.21 0.665 3.35 0.875 ;
 RECT 0.82 1.215 1.92 1.355 ;
 RECT 3.225 1.015 3.365 2.035 ;
 RECT 1.78 0.525 3.35 0.665 ;
 RECT 3.165 2.035 3.365 2.305 ;
 RECT 3.165 0.875 3.42 1.015 ;
 END
END DFFNASX2

MACRO DFFNX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.92 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.92 2.96 ;
 RECT 4.29 2.635 4.55 2.8 ;
 RECT 1.93 2.635 2.18 2.8 ;
 RECT 8.84 1.7 8.98 2.8 ;
 RECT 1.275 1.98 1.415 2.8 ;
 RECT 7.2 1.955 7.34 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.92 0.08 ;
 RECT 7.205 0.08 7.46 0.285 ;
 RECT 1.275 0.08 1.415 1.055 ;
 RECT 1.905 0.08 2.205 0.26 ;
 RECT 4.225 0.08 4.365 0.58 ;
 RECT 8.89 0.08 9.03 0.815 ;
 RECT 0.3 0.08 0.44 0.775 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.3 1.475 1.585 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.305 1.15 0.75 1.41 ;
 RECT 0.61 1.41 0.75 1.42 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.325 2.085 8.665 2.39 ;
 RECT 8.325 0.56 8.465 2.085 ;
 END
 ANTENNADIFFAREA 0.492 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.315 2.12 9.605 2.385 ;
 RECT 9.37 2.385 9.51 2.52 ;
 RECT 9.37 0.61 9.51 2.12 ;
 END
 ANTENNADIFFAREA 0.441 ;
 END Q

 OBS
 LAYER PO ;
 RECT 1.06 0.63 1.16 1.24 ;
 RECT 1.06 1.34 1.16 2.72 ;
 RECT 0.565 1.17 0.785 1.24 ;
 RECT 0.565 1.34 0.785 1.4 ;
 RECT 0.565 1.24 1.16 1.34 ;
 RECT 6.985 1.64 7.085 2.585 ;
 RECT 5.765 2.47 5.985 2.585 ;
 RECT 5.765 2.685 5.985 2.71 ;
 RECT 5.765 2.585 7.085 2.685 ;
 RECT 9.155 0.33 9.255 1.08 ;
 RECT 8.955 1.08 9.255 1.315 ;
 RECT 9.155 1.315 9.255 2.79 ;
 RECT 8.58 0.095 8.68 1.225 ;
 RECT 8.58 1.455 8.68 2.775 ;
 RECT 8 1.225 8.68 1.455 ;
 RECT 5.145 0.875 5.475 1.105 ;
 RECT 5.375 1.105 5.475 1.64 ;
 RECT 5.375 1.64 5.61 1.87 ;
 RECT 5.725 0.265 5.825 0.575 ;
 RECT 5.725 0.675 5.825 1.35 ;
 RECT 4.92 0.575 5.825 0.675 ;
 RECT 6.17 1.545 6.27 2.405 ;
 RECT 7.06 0.265 7.16 1.32 ;
 RECT 4.92 0.46 5.15 0.575 ;
 RECT 4.92 0.675 5.15 0.69 ;
 RECT 5.915 1.45 6.27 1.545 ;
 RECT 5.725 0.165 7.16 0.265 ;
 RECT 5.725 1.35 6.015 1.445 ;
 RECT 5.725 1.445 6.27 1.45 ;
 RECT 6.665 0.645 6.765 1.24 ;
 RECT 6.665 1.45 6.765 2.37 ;
 RECT 6.645 1.24 6.88 1.45 ;
 RECT 6.195 0.685 6.295 1.255 ;
 RECT 6.12 0.455 6.35 0.685 ;
 RECT 7.475 0.65 7.575 1.48 ;
 RECT 7.475 1.72 7.575 2.56 ;
 RECT 7.38 1.48 7.61 1.72 ;
 RECT 4.45 0.635 4.55 1.54 ;
 RECT 4.45 1.54 4.77 1.77 ;
 RECT 4.45 1.77 4.55 2.52 ;
 RECT 1.535 0.655 1.635 1.48 ;
 RECT 1.34 1.48 1.635 1.72 ;
 RECT 1.535 1.72 1.635 2.37 ;
 RECT 2.715 2.33 2.815 2.685 ;
 RECT 2.715 2.685 4.11 2.785 ;
 RECT 4.01 1.7 4.11 2.685 ;
 RECT 2.595 2.09 2.815 2.33 ;
 RECT 3.69 1.37 3.83 1.475 ;
 RECT 3.69 1.71 3.79 2.475 ;
 RECT 3.69 1.33 3.81 1.37 ;
 RECT 3.575 1.475 3.83 1.5 ;
 RECT 3.575 1.5 3.805 1.71 ;
 RECT 3.71 0.65 3.81 1.33 ;
 RECT 3.24 0.705 3.34 1.21 ;
 RECT 2.67 1.16 2.915 1.21 ;
 RECT 2.67 1.21 3.34 1.31 ;
 RECT 2.67 1.31 2.915 1.405 ;
 RECT 3.24 0.47 3.525 0.705 ;
 RECT 1.875 1.52 2.475 1.585 ;
 RECT 1.875 1.585 3.295 1.62 ;
 RECT 1.875 1.62 2.12 1.69 ;
 RECT 2.31 1.62 3.295 1.685 ;
 RECT 2.31 1.685 2.41 2.27 ;
 RECT 2.695 0.185 4.11 0.285 ;
 RECT 2.375 0.685 2.475 1.52 ;
 RECT 2.695 0.285 2.795 0.585 ;
 RECT 1.875 1.44 2.12 1.52 ;
 RECT 3.195 1.685 3.295 2.495 ;
 RECT 4.01 0.285 4.11 1.26 ;
 RECT 2.375 0.585 2.795 0.685 ;
 LAYER CO ;
 RECT 3.625 1.525 3.755 1.655 ;
 RECT 4.875 0.88 5.005 1.01 ;
 RECT 4.87 2.015 5 2.145 ;
 RECT 2.025 0.125 2.155 0.255 ;
 RECT 4.34 2.64 4.47 2.77 ;
 RECT 1.935 1.495 2.065 1.625 ;
 RECT 2 2.64 2.13 2.77 ;
 RECT 3.44 2.07 3.57 2.2 ;
 RECT 3.46 0.88 3.59 1.01 ;
 RECT 2.945 2.105 3.075 2.235 ;
 RECT 2.99 0.88 3.12 1.01 ;
 RECT 2.725 1.205 2.855 1.335 ;
 RECT 2.595 0.905 2.725 1.035 ;
 RECT 1.39 1.535 1.52 1.665 ;
 RECT 1.805 1.995 1.935 2.125 ;
 RECT 1.885 0.875 2.015 1.005 ;
 RECT 1.28 2.05 1.41 2.18 ;
 RECT 1.28 0.875 1.41 1.005 ;
 RECT 0.81 2.04 0.94 2.17 ;
 RECT 0.81 0.875 0.94 1.005 ;
 RECT 4.96 0.51 5.09 0.64 ;
 RECT 7.435 1.535 7.565 1.665 ;
 RECT 2.645 2.145 2.775 2.275 ;
 RECT 2.53 1.825 2.66 1.955 ;
 RECT 3.345 0.525 3.475 0.655 ;
 RECT 0.615 1.22 0.745 1.35 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 5.815 2.525 5.945 2.655 ;
 RECT 5.92 1.815 6.05 1.945 ;
 RECT 8.995 1.13 9.125 1.26 ;
 RECT 9.375 0.68 9.505 0.81 ;
 RECT 8.845 1.77 8.975 1.9 ;
 RECT 8.845 2.03 8.975 2.16 ;
 RECT 8.845 2.29 8.975 2.42 ;
 RECT 9.375 2.32 9.505 2.45 ;
 RECT 8.05 1.275 8.18 1.405 ;
 RECT 9.375 1.8 9.505 1.93 ;
 RECT 9.375 2.06 9.505 2.19 ;
 RECT 8.895 0.615 9.025 0.745 ;
 RECT 8.33 1.87 8.46 2 ;
 RECT 8.33 2.13 8.46 2.26 ;
 RECT 8.33 0.63 8.46 0.76 ;
 RECT 5.43 1.69 5.56 1.82 ;
 RECT 5.215 0.915 5.345 1.045 ;
 RECT 7.28 0.15 7.41 0.28 ;
 RECT 4.23 0.38 4.36 0.51 ;
 RECT 6.415 1.9 6.545 2.03 ;
 RECT 6.415 0.87 6.545 1 ;
 RECT 5.945 0.87 6.075 1 ;
 RECT 6.17 0.505 6.3 0.635 ;
 RECT 6.695 1.28 6.825 1.41 ;
 RECT 7.695 0.87 7.825 1 ;
 RECT 7.205 2.01 7.335 2.14 ;
 RECT 7.765 2.13 7.895 2.26 ;
 RECT 4.585 1.58 4.715 1.71 ;
 LAYER M1 ;
 RECT 6.69 1.245 7.905 1.385 ;
 RECT 7.76 1.105 7.9 1.245 ;
 RECT 7.76 1.385 7.9 2.33 ;
 RECT 7.69 0.36 7.83 0.965 ;
 RECT 7.69 0.965 7.9 1.105 ;
 RECT 6.69 1.21 6.83 1.245 ;
 RECT 6.69 1.385 6.83 1.465 ;
 RECT 8.61 0.36 8.75 1.125 ;
 RECT 7.69 0.22 8.75 0.36 ;
 RECT 8.99 1.055 9.13 1.125 ;
 RECT 8.99 1.265 9.13 1.335 ;
 RECT 8.61 1.125 9.13 1.265 ;
 RECT 3.275 0.52 3.875 0.66 ;
 RECT 3.735 0.66 3.875 0.79 ;
 RECT 4.505 0.505 5.14 0.645 ;
 RECT 3.735 0.79 4.645 0.93 ;
 RECT 4.505 0.645 4.645 0.79 ;
 RECT 4.865 1.05 5.005 1.185 ;
 RECT 4.08 1.185 5.005 1.325 ;
 RECT 4.865 1.325 5.005 2.215 ;
 RECT 4.865 1.015 5.415 1.05 ;
 RECT 3.56 1.52 4.22 1.66 ;
 RECT 4.805 0.91 5.415 1.015 ;
 RECT 4.805 0.875 5.075 0.91 ;
 RECT 4.08 1.325 4.22 1.52 ;
 RECT 0.89 1.01 1.03 1.195 ;
 RECT 0.89 1.335 1.03 2.035 ;
 RECT 0.74 0.87 1.03 1.01 ;
 RECT 0.74 2.035 1.03 2.175 ;
 RECT 1.555 0.67 1.695 1.195 ;
 RECT 0.89 1.195 1.695 1.335 ;
 RECT 1.555 0.53 2.505 0.67 ;
 RECT 2.365 0.22 3.125 0.36 ;
 RECT 2.985 0.36 3.125 0.875 ;
 RECT 2.94 2.035 3.14 2.17 ;
 RECT 2.94 2.17 3.08 2.305 ;
 RECT 3 1.015 3.14 2.035 ;
 RECT 2.365 0.36 2.505 0.53 ;
 RECT 2.92 0.875 3.195 1.015 ;
 RECT 2.59 1.385 2.73 1.82 ;
 RECT 2.46 1.825 2.78 1.96 ;
 RECT 2.46 1.82 2.73 1.825 ;
 RECT 2.64 1.96 2.78 2.345 ;
 RECT 2.59 0.84 2.73 1.155 ;
 RECT 2.59 1.155 2.86 1.385 ;
 RECT 2.32 2.515 3.855 2.65 ;
 RECT 2.32 2.65 3.61 2.655 ;
 RECT 3.175 2.51 3.855 2.515 ;
 RECT 2.32 2.49 2.46 2.515 ;
 RECT 1.8 1.63 1.94 2.35 ;
 RECT 1.8 1.475 2.14 1.63 ;
 RECT 1.88 0.825 2.02 1.475 ;
 RECT 3.715 2.495 3.855 2.51 ;
 RECT 1.8 2.35 2.46 2.49 ;
 RECT 5.585 0.58 6.375 0.64 ;
 RECT 5.585 0.64 6.045 0.72 ;
 RECT 5.865 0.5 6.375 0.58 ;
 RECT 5.145 1.21 5.725 1.35 ;
 RECT 5.745 2.24 5.885 2.52 ;
 RECT 5.145 1.35 5.285 2.1 ;
 RECT 5.145 2.24 5.285 2.355 ;
 RECT 5.145 2.1 5.885 2.24 ;
 RECT 3.715 2.355 5.285 2.495 ;
 RECT 5.585 0.72 5.725 1.21 ;
 RECT 5.745 2.52 6.015 2.66 ;
 RECT 3.28 1.82 4.72 1.96 ;
 RECT 3.28 1.22 3.595 1.36 ;
 RECT 3.455 0.805 3.595 1.22 ;
 RECT 4.58 1.51 4.72 1.82 ;
 RECT 3.365 1.96 3.645 2.215 ;
 RECT 3.28 1.36 3.42 1.82 ;
 RECT 6.41 1.815 6.62 1.895 ;
 RECT 6.41 0.805 6.55 1.675 ;
 RECT 6.34 1.895 6.62 2.035 ;
 RECT 6.41 1.675 7.27 1.815 ;
 RECT 7.13 1.67 7.27 1.675 ;
 RECT 8.045 1.205 8.185 2.505 ;
 RECT 7.13 1.53 7.62 1.67 ;
 RECT 7.48 2.505 8.185 2.645 ;
 RECT 7.48 1.67 7.62 2.505 ;
 RECT 5.425 1.685 6.08 1.81 ;
 RECT 5.94 1.005 6.08 1.685 ;
 RECT 5.425 1.81 6.12 1.825 ;
 RECT 5.425 1.825 5.565 1.89 ;
 RECT 5.425 1.62 5.565 1.685 ;
 RECT 5.85 1.825 6.12 1.95 ;
 RECT 5.87 0.865 6.15 1.005 ;
 END
END DFFNX1

MACRO PMT2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.115 1.63 1.17 1.77 ;
 RECT 0.115 1.77 0.49 1.92 ;
 RECT 0.115 1.61 0.49 1.63 ;
 END
 ANTENNADIFFAREA 0.426 ;
 END D

 PIN S
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.46 2.43 1.64 2.57 ;
 RECT 0.995 2.11 1.265 2.43 ;
 END
 ANTENNADIFFAREA 0.672 ;
 END S

 PIN G
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.645 0.73 0.995 1.105 ;
 END
 ANTENNAGATEAREA 0.224 ;
 END G

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 RECT 2 1.565 2.16 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 1.24 1.305 1.34 2.785 ;
 RECT 0.76 1.245 1.34 1.345 ;
 RECT 0.76 1.025 0.86 2.785 ;
 RECT 0.705 0.795 0.935 1.025 ;
 LAYER CO ;
 RECT 0.755 0.845 0.885 0.975 ;
 RECT 2.015 1.62 2.145 1.75 ;
 RECT 2.015 1.88 2.145 2.01 ;
 RECT 1.46 2.435 1.59 2.565 ;
 RECT 0.99 1.635 1.12 1.765 ;
 RECT 0.51 2.435 0.64 2.565 ;
 END
END PMT2

MACRO PMT3
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN S
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.115 1.63 2.11 1.77 ;
 RECT 0.115 1.77 0.475 1.91 ;
 END
 ANTENNADIFFAREA 0.84 ;
 END S

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.46 2.43 2.58 2.57 ;
 RECT 0.965 2.11 1.275 2.43 ;
 END
 ANTENNADIFFAREA 1.086 ;
 END D

 PIN G
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.655 0.745 1 1.11 ;
 END
 ANTENNAGATEAREA 0.448 ;
 END G

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 2.96 1.835 3.12 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 2.18 1.305 2.28 2.785 ;
 RECT 1.71 1.305 1.81 2.785 ;
 RECT 1.24 1.305 1.34 2.785 ;
 RECT 0.76 1.25 2.28 1.35 ;
 RECT 0.76 1.04 0.86 2.785 ;
 RECT 0.695 0.81 0.925 1.04 ;
 LAYER CO ;
 RECT 0.745 0.86 0.875 0.99 ;
 RECT 2.975 1.885 3.105 2.015 ;
 RECT 2.975 2.175 3.105 2.305 ;
 RECT 1.93 1.635 2.06 1.765 ;
 RECT 2.4 2.435 2.53 2.565 ;
 RECT 1.46 2.435 1.59 2.565 ;
 RECT 0.99 1.635 1.12 1.765 ;
 RECT 0.51 2.435 0.64 2.565 ;
 END
END PMT3

MACRO RSDFFNSRARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 28.48 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.185 1.16 19.55 1.4 ;
 RECT 19.41 0.51 19.55 1.16 ;
 RECT 20.47 1.905 20.61 1.91 ;
 RECT 19.41 1.765 20.61 1.905 ;
 RECT 20.47 0.56 20.61 1.765 ;
 RECT 19.41 1.905 19.55 1.915 ;
 RECT 19.41 1.4 19.55 1.765 ;
 END
 ANTENNADIFFAREA 0.689 ;
 END Q

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.495 0.455 7.825 0.485 ;
 RECT 11.335 0.245 13.46 0.385 ;
 RECT 7.525 0.755 8.6 0.875 ;
 RECT 7.48 0.485 7.825 0.735 ;
 RECT 7.48 0.735 8.6 0.755 ;
 RECT 8.46 0.22 10.095 0.36 ;
 RECT 8.46 0.36 8.6 0.735 ;
 RECT 9.955 0.525 10.5 0.665 ;
 RECT 10.36 1.005 11.455 1.01 ;
 RECT 10.36 0.87 11.475 1.005 ;
 RECT 13.315 0.385 13.455 1.09 ;
 RECT 13.315 1.09 15.715 1.23 ;
 RECT 15.575 0.81 15.715 1.09 ;
 RECT 15.575 0.6 15.865 0.81 ;
 RECT 9.955 0.36 10.095 0.525 ;
 RECT 11.335 0.385 11.475 0.87 ;
 RECT 10.36 0.665 10.5 0.87 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.79 1.475 5.12 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.35 1.15 10.68 1.49 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.685 1.84 18.04 1.99 ;
 RECT 17.685 1.75 19.045 1.84 ;
 RECT 18.905 0.915 19.045 1.7 ;
 RECT 17.9 1.7 19.045 1.75 ;
 RECT 17.9 0.905 18.04 1.7 ;
 RECT 18.905 1.84 19.045 1.885 ;
 END
 ANTENNADIFFAREA 0.352 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 28.48 2.96 ;
 RECT 1.36 2.005 1.5 2.8 ;
 RECT 3.27 2.03 3.41 2.8 ;
 RECT 4.74 1.98 4.88 2.8 ;
 RECT 0.385 1.74 0.525 2.8 ;
 RECT 5.415 2.34 5.665 2.8 ;
 RECT 8.67 2.07 8.81 2.8 ;
 RECT 10.77 2.375 10.91 2.8 ;
 RECT 16.32 2.57 16.46 2.8 ;
 RECT 18.305 2.57 18.445 2.8 ;
 RECT 15.42 2.57 15.56 2.8 ;
 RECT 19.885 2.57 20.025 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 28.48 0.08 ;
 RECT 10.895 0.59 11.17 0.73 ;
 RECT 18.335 0.28 18.6 0.44 ;
 RECT 4.74 0.08 4.88 1.055 ;
 RECT 3.27 0.08 3.41 0.78 ;
 RECT 1.36 0.08 1.5 0.97 ;
 RECT 0.35 0.08 0.49 0.775 ;
 RECT 8.085 0.08 8.32 0.595 ;
 RECT 5.485 0.08 5.625 0.39 ;
 RECT 14.82 0.08 14.96 0.945 ;
 RECT 16.325 0.08 16.465 0.525 ;
 RECT 22.995 0.08 23.135 0.31 ;
 RECT 19.97 0.08 20.11 0.82 ;
 RECT 25.345 0.08 25.585 0.31 ;
 RECT 24.21 0.08 24.35 0.325 ;
 RECT 10.96 0.08 11.1 0.59 ;
 RECT 18.39 0.08 18.53 0.28 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.33 1.155 2.75 1.415 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.18 1.475 1.705 1.75 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.965 1.13 2.105 1.48 ;
 RECT 1.87 1.63 2.815 1.79 ;
 RECT 1.87 1.48 2.115 1.63 ;
 RECT 2.665 1.79 2.805 1.845 ;
 RECT 2.665 1.57 2.805 1.63 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.905 1.41 27.245 1.775 ;
 RECT 25.225 1.965 27.09 2.105 ;
 RECT 22.995 2.195 25.365 2.335 ;
 RECT 25.225 1.41 25.365 1.965 ;
 RECT 26.95 1.775 27.09 1.965 ;
 RECT 22.995 1.365 23.135 2.195 ;
 RECT 24.38 1.345 24.52 2.195 ;
 RECT 25.225 2.105 25.365 2.195 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 21.565 0.57 22.045 0.78 ;
 RECT 21.565 0.78 21.935 0.865 ;
 RECT 21.565 0.565 21.935 0.57 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 OBS
 LAYER PO ;
 RECT 25.645 0.09 26.755 0.19 ;
 RECT 25.645 0.19 25.745 0.94 ;
 RECT 22.02 2.64 26.755 2.74 ;
 RECT 22.02 1.075 22.35 1.175 ;
 RECT 22.78 0.87 22.88 2.175 ;
 RECT 21.815 0.77 23.35 0.78 ;
 RECT 22.78 0.73 23.35 0.77 ;
 RECT 25.48 1.125 25.58 2.175 ;
 RECT 21.82 0.78 23.35 0.83 ;
 RECT 21.82 0.83 22.88 0.87 ;
 RECT 23.25 0.19 23.35 0.73 ;
 RECT 22.78 0.185 22.88 0.73 ;
 RECT 21.815 0.57 22.045 0.77 ;
 RECT 22.78 2.175 25.58 2.275 ;
 RECT 25.955 0.37 26.055 1.01 ;
 RECT 25.955 1.01 26.205 1.22 ;
 RECT 25.955 1.22 26.055 2.245 ;
 RECT 25.955 2.245 26.24 2.455 ;
 RECT 24.47 0.355 24.57 0.985 ;
 RECT 24.64 1.215 24.74 1.815 ;
 RECT 24.08 1.115 24.74 1.215 ;
 RECT 24.08 0.985 24.57 1.115 ;
 RECT 24.975 0.355 25.205 0.465 ;
 RECT 24.47 0.255 25.205 0.355 ;
 RECT 23.12 1.01 23.355 1.22 ;
 RECT 23.255 1.22 23.355 1.995 ;
 RECT 11.615 2.69 13.265 2.695 ;
 RECT 13.09 2.54 13.265 2.69 ;
 RECT 12.405 2.695 13.265 2.79 ;
 RECT 11.615 0.655 11.715 2.595 ;
 RECT 11.615 2.595 12.505 2.69 ;
 RECT 13.09 2.33 13.32 2.54 ;
 RECT 15.675 0.81 15.775 2.21 ;
 RECT 15.635 0.6 15.865 0.81 ;
 RECT 9.4 1.575 9.5 2.485 ;
 RECT 9.91 1.41 10.14 1.475 ;
 RECT 9.91 1.575 10.14 1.62 ;
 RECT 9.4 1.475 10.14 1.575 ;
 RECT 10.325 1.45 10.425 1.655 ;
 RECT 10.325 1.755 10.425 2.57 ;
 RECT 10.325 0.655 10.425 1.13 ;
 RECT 10.325 1.23 10.425 1.24 ;
 RECT 9.41 0.66 9.51 1.13 ;
 RECT 10.325 1.655 11.285 1.755 ;
 RECT 11.185 1.755 11.285 2.355 ;
 RECT 10.325 1.24 10.58 1.45 ;
 RECT 9.41 1.13 10.425 1.23 ;
 RECT 17.155 0.29 18.265 0.39 ;
 RECT 18.165 0.39 18.265 1.4 ;
 RECT 18.165 1.5 18.265 2.11 ;
 RECT 18.655 0.505 18.755 1.4 ;
 RECT 18.655 1.5 18.755 2.11 ;
 RECT 17.155 0.225 17.385 0.29 ;
 RECT 17.155 0.39 17.385 0.435 ;
 RECT 18.165 1.4 18.755 1.5 ;
 RECT 15.205 0.835 15.305 2.21 ;
 RECT 15.205 0.47 15.37 0.625 ;
 RECT 14.32 0.455 15.37 0.47 ;
 RECT 14.32 0.47 14.55 0.665 ;
 RECT 14.43 0.37 15.37 0.455 ;
 RECT 15.205 0.625 15.435 0.835 ;
 RECT 16.575 1.635 16.675 1.66 ;
 RECT 16.575 1.66 16.83 1.87 ;
 RECT 16.575 1.87 16.675 2.565 ;
 RECT 12.945 0.885 13.175 0.925 ;
 RECT 12.945 0.925 13.79 1.025 ;
 RECT 12.945 1.025 13.175 1.095 ;
 RECT 13.625 0.795 13.79 0.925 ;
 RECT 13.625 0.585 13.855 0.795 ;
 RECT 5.775 1.62 5.875 2.375 ;
 RECT 5.84 0.185 12.75 0.19 ;
 RECT 5.84 0.19 7.995 0.285 ;
 RECT 5.84 0.285 5.94 1.52 ;
 RECT 12.65 1.29 13.67 1.39 ;
 RECT 12.65 0.19 12.75 1.29 ;
 RECT 6.66 1.565 6.76 2.375 ;
 RECT 5.34 1.44 5.585 1.52 ;
 RECT 5.34 1.62 5.585 1.69 ;
 RECT 5.34 1.52 5.94 1.62 ;
 RECT 7.895 0.285 7.995 1.24 ;
 RECT 7.895 0.09 12.75 0.185 ;
 RECT 13.44 1.285 13.67 1.29 ;
 RECT 13.44 1.39 13.67 1.615 ;
 RECT 5.775 2.375 6.76 2.475 ;
 RECT 8.945 0.47 9.13 0.5 ;
 RECT 16.58 0.19 16.68 1.18 ;
 RECT 14.04 0.09 16.68 0.19 ;
 RECT 14.04 0.19 14.14 1.795 ;
 RECT 13.155 1.71 13.255 1.795 ;
 RECT 12.685 1.71 12.785 2.445 ;
 RECT 12.135 0.47 12.235 1.61 ;
 RECT 13.155 1.795 14.14 1.895 ;
 RECT 12.135 1.61 13.255 1.71 ;
 RECT 8.945 0.37 12.235 0.47 ;
 RECT 8.9 0.5 9.13 0.71 ;
 RECT 16.85 1.25 17.11 1.3 ;
 RECT 17.01 0.61 17.11 1.25 ;
 RECT 16.85 1.4 17.11 1.46 ;
 RECT 17.01 1.46 17.11 2.56 ;
 RECT 17.54 0.84 17.64 1.3 ;
 RECT 16.85 1.3 17.64 1.4 ;
 RECT 17.525 0.63 17.755 0.84 ;
 RECT 2.755 1.82 2.855 2.735 ;
 RECT 2.615 1.59 2.855 1.82 ;
 RECT 1.95 0.555 2.05 1.145 ;
 RECT 1.91 1.145 2.155 1.385 ;
 RECT 3.525 0.335 3.625 1.155 ;
 RECT 3.525 1.365 3.625 2.745 ;
 RECT 3.335 1.155 3.625 1.365 ;
 RECT 1.145 1.475 1.715 1.75 ;
 RECT 1.145 0.555 1.245 1.475 ;
 RECT 1.145 1.75 1.245 2.685 ;
 RECT 1.615 0.555 1.715 1.475 ;
 RECT 1.615 1.75 1.715 2.735 ;
 RECT 2.335 1.41 2.435 1.645 ;
 RECT 2.565 0.555 2.665 1.18 ;
 RECT 2.285 1.745 2.385 2.735 ;
 RECT 2.285 1.645 2.435 1.745 ;
 RECT 2.335 1.18 2.665 1.41 ;
 RECT 5 0.57 5.1 1.495 ;
 RECT 4.805 1.495 5.1 1.745 ;
 RECT 5 1.745 5.1 2.37 ;
 RECT 7.155 1.33 7.295 1.475 ;
 RECT 7.155 1.71 7.255 2.475 ;
 RECT 7.195 0.65 7.295 1.33 ;
 RECT 7.155 1.475 7.385 1.71 ;
 RECT 2.85 0.175 3.155 0.405 ;
 RECT 3.055 0.405 3.155 2.735 ;
 RECT 7.595 0.715 7.695 1.61 ;
 RECT 7.63 1.71 7.73 2.48 ;
 RECT 7.595 1.61 7.73 1.71 ;
 RECT 7.475 0.485 7.715 0.715 ;
 RECT 4.285 0.27 4.625 0.52 ;
 RECT 4.525 0.52 4.625 2.465 ;
 RECT 11.22 0.655 11.32 1.24 ;
 RECT 11.09 1.24 11.32 1.475 ;
 RECT 8.76 1.61 9.025 1.82 ;
 RECT 8.925 1.82 9.025 2.49 ;
 RECT 8.555 0.66 8.655 1.51 ;
 RECT 8.555 1.51 9.025 1.61 ;
 RECT 8.24 2.465 8.555 2.71 ;
 RECT 8.455 1.79 8.555 2.465 ;
 RECT 6.705 0.705 6.805 1.17 ;
 RECT 6.705 0.47 6.99 0.705 ;
 RECT 6.12 1.27 6.365 1.46 ;
 RECT 6.12 1.17 6.805 1.27 ;
 RECT 19.655 1.285 20.35 1.385 ;
 RECT 20.25 0.19 20.35 1.285 ;
 RECT 19.655 1.385 19.865 1.435 ;
 RECT 19.655 1.2 19.865 1.285 ;
 RECT 19.67 0.385 19.77 1.2 ;
 RECT 19.67 1.435 19.77 2.645 ;
 RECT 20.25 1.385 20.35 2.645 ;
 RECT 20.25 0.09 21.395 0.19 ;
 RECT 21.165 0.19 21.395 0.435 ;
 RECT 23.56 0.19 23.66 0.97 ;
 RECT 23.56 0.97 23.8 1.18 ;
 RECT 23.56 1.18 23.66 1.975 ;
 RECT 22.02 1.175 22.305 1.305 ;
 RECT 22.02 1.305 22.12 2.64 ;
 RECT 26.655 0.19 26.755 2.64 ;
 LAYER CO ;
 RECT 11.875 0.875 12.005 1.005 ;
 RECT 7.205 1.525 7.335 1.655 ;
 RECT 4.345 0.325 4.475 0.455 ;
 RECT 25.395 0.115 25.525 0.245 ;
 RECT 24.215 0.11 24.345 0.24 ;
 RECT 22.53 1.4 22.66 1.53 ;
 RECT 24.695 0.59 24.825 0.72 ;
 RECT 3.745 2.05 3.875 2.18 ;
 RECT 1.37 1.55 1.5 1.68 ;
 RECT 3.275 2.09 3.405 2.22 ;
 RECT 2.49 1.23 2.62 1.36 ;
 RECT 1.365 2.315 1.495 2.445 ;
 RECT 2.67 1.64 2.8 1.77 ;
 RECT 25.23 1.465 25.36 1.595 ;
 RECT 24.385 1.42 24.515 1.55 ;
 RECT 26.175 1.44 26.305 1.57 ;
 RECT 23 1.45 23.13 1.58 ;
 RECT 12.905 1.87 13.035 2 ;
 RECT 4.865 1.55 4.995 1.68 ;
 RECT 6.925 0.88 7.055 1.01 ;
 RECT 12.4 0.595 12.53 0.725 ;
 RECT 10.075 1.885 10.205 2.015 ;
 RECT 5.995 1.825 6.125 1.955 ;
 RECT 12.4 1.9 12.53 2.03 ;
 RECT 7.855 1.825 7.985 1.955 ;
 RECT 8.205 2.125 8.335 2.255 ;
 RECT 4.275 2.115 4.405 2.245 ;
 RECT 0.355 0.59 0.485 0.72 ;
 RECT 11.875 1.945 12.005 2.075 ;
 RECT 10.075 0.88 10.205 1.01 ;
 RECT 5.4 1.495 5.53 1.625 ;
 RECT 19.89 2.64 20.02 2.77 ;
 RECT 7.53 0.53 7.66 0.66 ;
 RECT 11.14 1.28 11.27 1.41 ;
 RECT 17.905 1.705 18.035 1.835 ;
 RECT 5.22 1.995 5.35 2.125 ;
 RECT 20.475 1.71 20.605 1.84 ;
 RECT 16.33 0.33 16.46 0.46 ;
 RECT 18.91 1.705 19.04 1.835 ;
 RECT 12.905 0.595 13.035 0.725 ;
 RECT 17.23 1.78 17.36 1.91 ;
 RECT 18.395 0.305 18.525 0.435 ;
 RECT 19.975 0.62 20.105 0.75 ;
 RECT 6.905 2.07 7.035 2.2 ;
 RECT 6.175 1.265 6.305 1.395 ;
 RECT 21.215 0.265 21.345 0.395 ;
 RECT 23.62 1.01 23.75 1.14 ;
 RECT 26.025 1.05 26.155 1.18 ;
 RECT 22.125 1.135 22.255 1.265 ;
 RECT 21.865 0.61 21.995 0.74 ;
 RECT 24.13 1.025 24.26 1.155 ;
 RECT 26.06 2.285 26.19 2.415 ;
 RECT 25.025 0.295 25.155 0.425 ;
 RECT 23.17 1.05 23.3 1.18 ;
 RECT 15.255 0.665 15.385 0.795 ;
 RECT 13.14 2.37 13.27 2.5 ;
 RECT 15.685 0.64 15.815 0.77 ;
 RECT 9.96 1.45 10.09 1.58 ;
 RECT 10.4 1.28 10.53 1.41 ;
 RECT 12.995 0.925 13.125 1.055 ;
 RECT 17.205 0.265 17.335 0.395 ;
 RECT 17.575 0.67 17.705 0.8 ;
 RECT 14.37 0.495 14.5 0.625 ;
 RECT 16.65 1.7 16.78 1.83 ;
 RECT 13.675 0.625 13.805 0.755 ;
 RECT 13.49 1.445 13.62 1.575 ;
 RECT 8.95 0.54 9.08 0.67 ;
 RECT 16.9 1.29 17.03 1.42 ;
 RECT 1.365 0.775 1.495 0.905 ;
 RECT 3.275 2.35 3.405 2.48 ;
 RECT 2.505 2.115 2.635 2.245 ;
 RECT 1.365 2.055 1.495 2.185 ;
 RECT 0.895 2.055 1.025 2.185 ;
 RECT 3.745 1.79 3.875 1.92 ;
 RECT 1.97 1.195 2.1 1.325 ;
 RECT 3.385 1.195 3.515 1.325 ;
 RECT 2.9 0.225 3.03 0.355 ;
 RECT 0.895 0.775 1.025 0.905 ;
 RECT 3.745 0.775 3.875 0.905 ;
 RECT 3.275 0.585 3.405 0.715 ;
 RECT 2.31 0.775 2.44 0.905 ;
 RECT 17.905 0.975 18.035 1.105 ;
 RECT 5.49 0.21 5.62 0.34 ;
 RECT 18.31 2.64 18.44 2.77 ;
 RECT 9.145 2.015 9.275 2.145 ;
 RECT 7.375 2.125 7.505 2.255 ;
 RECT 14.955 1.7 15.085 1.83 ;
 RECT 5.485 2.345 5.615 2.475 ;
 RECT 19.695 1.25 19.825 1.38 ;
 RECT 0.355 0.33 0.485 0.46 ;
 RECT 26.175 0.59 26.305 0.72 ;
 RECT 23.78 1.46 23.91 1.59 ;
 RECT 23.78 0.41 23.91 0.54 ;
 RECT 24.86 1.38 24.99 1.51 ;
 RECT 22.28 0.505 22.41 0.635 ;
 RECT 26.955 1.45 27.085 1.58 ;
 RECT 23 0.11 23.13 0.24 ;
 RECT 16.325 2.64 16.455 2.77 ;
 RECT 0.39 2.085 0.52 2.215 ;
 RECT 10.775 2.445 10.905 2.575 ;
 RECT 4.275 0.79 4.405 0.92 ;
 RECT 15.425 2.64 15.555 2.77 ;
 RECT 18.91 0.975 19.04 1.105 ;
 RECT 0.39 1.825 0.52 1.955 ;
 RECT 15.895 1.705 16.025 1.835 ;
 RECT 6.81 0.525 6.94 0.655 ;
 RECT 6.455 0.88 6.585 1.01 ;
 RECT 19.415 0.62 19.545 0.75 ;
 RECT 8.28 2.515 8.41 2.645 ;
 RECT 8.135 0.455 8.265 0.585 ;
 RECT 6.06 0.905 6.19 1.035 ;
 RECT 17.23 0.83 17.36 0.96 ;
 RECT 20.475 0.63 20.605 0.76 ;
 RECT 14.825 0.745 14.955 0.875 ;
 RECT 4.745 2.05 4.875 2.18 ;
 RECT 10.965 0.595 11.095 0.725 ;
 RECT 6.41 2.105 6.54 2.235 ;
 RECT 9.63 2.07 9.76 2.2 ;
 RECT 8.675 2.135 8.805 2.265 ;
 RECT 8.815 1.63 8.945 1.76 ;
 RECT 19.415 1.725 19.545 1.855 ;
 RECT 5.35 0.88 5.48 1.01 ;
 RECT 9.63 0.88 9.76 1.01 ;
 RECT 15.93 0.96 16.06 1.09 ;
 RECT 0.39 2.345 0.52 2.475 ;
 RECT 4.745 0.79 4.875 0.92 ;
 RECT 9.145 0.93 9.275 1.06 ;
 LAYER M1 ;
 RECT 9.14 1.44 9.28 2.215 ;
 RECT 7.865 1.3 9.28 1.44 ;
 RECT 5.26 1.63 5.4 1.99 ;
 RECT 5.26 1.475 5.605 1.63 ;
 RECT 5.345 0.81 5.485 1.475 ;
 RECT 5.15 1.99 5.4 2.13 ;
 RECT 6.83 1.96 7.11 2.215 ;
 RECT 6.92 0.805 7.06 1.22 ;
 RECT 6.85 1.22 7.06 1.36 ;
 RECT 6.85 1.36 6.99 1.82 ;
 RECT 6.83 1.89 8.325 1.96 ;
 RECT 6.85 1.82 8.325 1.89 ;
 RECT 8.185 1.79 8.325 1.82 ;
 RECT 8.76 1.58 9 1.65 ;
 RECT 8.76 1.79 9 1.835 ;
 RECT 8.185 1.65 9 1.79 ;
 RECT 2.96 0.91 3.1 1.19 ;
 RECT 2.96 1.33 3.1 2.11 ;
 RECT 2.255 0.77 3.1 0.91 ;
 RECT 2.45 2.11 3.1 2.25 ;
 RECT 2.96 1.19 3.52 1.33 ;
 RECT 3.38 1.145 3.52 1.19 ;
 RECT 3.38 1.33 3.52 1.375 ;
 RECT 24.08 1.195 24.22 1.32 ;
 RECT 23.775 1.46 23.915 1.735 ;
 RECT 24.095 0.705 24.235 0.985 ;
 RECT 23.775 0.33 23.915 0.565 ;
 RECT 23.775 1.32 24.22 1.46 ;
 RECT 24.08 0.985 24.31 1.195 ;
 RECT 23.775 0.565 24.235 0.705 ;
 RECT 24.855 1.22 24.995 1.58 ;
 RECT 24.69 0.48 24.83 1.08 ;
 RECT 25.975 1.01 26.205 1.08 ;
 RECT 24.69 1.08 26.205 1.22 ;
 RECT 25.065 0.465 25.205 0.685 ;
 RECT 24.975 0.255 25.205 0.465 ;
 RECT 25.065 0.685 26.625 0.825 ;
 RECT 26.485 0.825 26.625 1.36 ;
 RECT 26.17 1.5 26.31 1.705 ;
 RECT 26.17 0.485 26.31 0.685 ;
 RECT 26.17 1.36 26.625 1.5 ;
 RECT 22.525 1.2 22.665 1.725 ;
 RECT 22.075 1.17 22.665 1.2 ;
 RECT 22.075 1.2 22.305 1.305 ;
 RECT 22.35 0.64 22.49 0.99 ;
 RECT 22.215 0.99 22.525 1.03 ;
 RECT 22.23 0.5 22.49 0.64 ;
 RECT 23.12 1.01 23.35 1.03 ;
 RECT 22.07 1.03 23.35 1.17 ;
 RECT 23.12 1.17 23.35 1.22 ;
 RECT 21.165 0.36 21.395 0.435 ;
 RECT 22.63 0.36 22.77 0.54 ;
 RECT 21.165 0.225 22.77 0.36 ;
 RECT 21.17 0.22 22.77 0.225 ;
 RECT 23.495 0.535 23.635 0.54 ;
 RECT 23.495 0.68 23.635 0.97 ;
 RECT 23.495 0.97 23.8 1.18 ;
 RECT 22.63 0.54 23.635 0.68 ;
 RECT 17.525 0.72 17.755 0.84 ;
 RECT 17.52 0.58 18.94 0.72 ;
 RECT 18.8 0.37 18.94 0.58 ;
 RECT 19.69 0.37 19.83 1.46 ;
 RECT 18.8 0.23 19.83 0.37 ;
 RECT 15.205 0.36 15.435 0.835 ;
 RECT 16.005 0.36 16.145 0.665 ;
 RECT 15.205 0.22 16.15 0.36 ;
 RECT 17.225 0.435 17.365 0.665 ;
 RECT 16.005 0.665 17.365 0.805 ;
 RECT 17.225 0.805 17.365 1.98 ;
 RECT 17.225 0.22 17.365 0.225 ;
 RECT 17.155 0.225 17.385 0.435 ;
 RECT 12.9 0.525 13.04 0.885 ;
 RECT 12.9 1.095 13.04 2.065 ;
 RECT 12.9 0.885 13.175 1.095 ;
 RECT 9.625 0.82 9.765 2.225 ;
 RECT 10.475 2.165 10.615 2.225 ;
 RECT 9.625 2.225 10.615 2.365 ;
 RECT 11.87 0.765 12.01 2.025 ;
 RECT 12.395 0.525 12.535 2.025 ;
 RECT 10.475 2.025 12.535 2.165 ;
 RECT 13.625 0.585 14.55 0.63 ;
 RECT 13.625 0.63 13.855 0.795 ;
 RECT 13.65 0.49 14.55 0.585 ;
 RECT 14.32 0.455 14.55 0.49 ;
 RECT 14.32 0.63 14.55 0.665 ;
 RECT 6.055 1.435 6.195 1.82 ;
 RECT 6.055 1.96 6.195 2.51 ;
 RECT 6.055 0.5 6.195 1.225 ;
 RECT 6.055 1.225 6.355 1.435 ;
 RECT 5.925 1.82 6.195 1.96 ;
 RECT 6.055 2.51 8.53 2.65 ;
 RECT 4.05 1.335 4.19 2.11 ;
 RECT 4.05 2.25 4.19 2.255 ;
 RECT 4.05 0.925 4.19 1.195 ;
 RECT 4.05 2.11 4.475 2.25 ;
 RECT 4.05 0.785 4.475 0.925 ;
 RECT 4.05 1.195 5.16 1.335 ;
 RECT 5.02 0.67 5.16 1.195 ;
 RECT 6.45 0.36 6.59 0.9 ;
 RECT 6.525 1.08 6.665 1.945 ;
 RECT 5.765 0.22 6.59 0.36 ;
 RECT 6.405 2.17 6.545 2.305 ;
 RECT 6.405 1.945 6.665 2.17 ;
 RECT 6.45 0.9 6.665 1.08 ;
 RECT 5.765 0.36 5.905 0.53 ;
 RECT 5.02 0.53 5.905 0.67 ;
 RECT 6.74 0.52 7.34 0.66 ;
 RECT 7.2 0.66 7.34 1.015 ;
 RECT 8.745 0.505 9.13 0.71 ;
 RECT 7.2 1.015 8.885 1.155 ;
 RECT 8.745 0.71 8.885 1.015 ;
 RECT 8.9 0.5 9.13 0.505 ;
 RECT 0.89 0.72 1.03 1.195 ;
 RECT 0.89 1.335 1.03 2.27 ;
 RECT 0.89 1.195 1.815 1.335 ;
 RECT 1.675 0.36 1.815 1.195 ;
 RECT 1.675 0.22 3.1 0.36 ;
 RECT 3.74 0.57 3.88 2.25 ;
 RECT 4.235 0.22 4.6 0.43 ;
 RECT 4.235 0.57 4.6 0.615 ;
 RECT 3.74 0.43 4.6 0.57 ;
 RECT 13.09 2.42 13.32 2.54 ;
 RECT 21.555 2.42 21.695 2.505 ;
 RECT 13.09 2.28 21.695 2.42 ;
 RECT 26.01 2.455 26.15 2.505 ;
 RECT 26.01 2.245 26.24 2.455 ;
 RECT 21.555 2.505 26.15 2.645 ;
 RECT 14.95 1.51 15.09 1.695 ;
 RECT 14.88 1.695 15.16 1.835 ;
 RECT 15.89 1.51 16.03 1.7 ;
 RECT 15.925 1.095 16.065 1.37 ;
 RECT 14.95 1.37 17.08 1.51 ;
 RECT 16.85 1.25 17.08 1.37 ;
 RECT 15.825 1.7 16.1 1.84 ;
 RECT 15.855 0.955 16.135 1.095 ;
 RECT 10.07 1.62 10.21 1.735 ;
 RECT 10.07 1.875 10.21 2.085 ;
 RECT 10.07 0.81 10.21 1.41 ;
 RECT 9.91 1.41 10.21 1.62 ;
 RECT 11.135 1.415 11.275 1.735 ;
 RECT 10.07 1.735 11.275 1.875 ;
 RECT 11.07 1.275 11.34 1.415 ;
 RECT 16.6 1.87 16.785 1.985 ;
 RECT 13.435 1.43 13.67 1.615 ;
 RECT 13.44 1.405 13.67 1.43 ;
 RECT 13.435 1.615 13.575 1.985 ;
 RECT 16.6 1.66 16.83 1.87 ;
 RECT 13.435 1.985 16.785 2.125 ;
 RECT 7.305 2.12 8.405 2.26 ;
 RECT 7.135 1.52 8.005 1.66 ;
 RECT 7.865 1.44 8.005 1.52 ;
 RECT 9.14 0.865 9.28 1.3 ;
 END
END RSDFFNSRARX1

MACRO RSDFFNSRARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 29.44 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.41 1.765 21.55 1.905 ;
 RECT 19.185 1.16 19.55 1.4 ;
 RECT 19.41 0.51 19.55 1.16 ;
 RECT 21.41 1.905 21.55 1.91 ;
 RECT 21.41 0.56 21.55 1.765 ;
 RECT 20.47 1.905 20.61 1.91 ;
 RECT 20.47 0.56 20.61 1.765 ;
 RECT 19.41 1.905 19.55 1.915 ;
 RECT 19.41 1.4 19.55 1.765 ;
 END
 ANTENNADIFFAREA 1.434 ;
 END Q

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.495 0.455 7.825 0.485 ;
 RECT 11.335 0.245 13.46 0.385 ;
 RECT 7.525 0.755 8.6 0.875 ;
 RECT 7.48 0.485 7.825 0.735 ;
 RECT 7.48 0.735 8.6 0.755 ;
 RECT 8.46 0.36 8.6 0.735 ;
 RECT 11.335 1.02 11.475 1.025 ;
 RECT 10.36 0.88 11.475 1.02 ;
 RECT 13.315 0.385 13.455 1.09 ;
 RECT 13.315 1.09 15.715 1.23 ;
 RECT 15.575 0.81 15.715 1.09 ;
 RECT 15.575 0.6 15.865 0.81 ;
 RECT 10.36 0.36 10.5 0.88 ;
 RECT 8.46 0.22 10.5 0.36 ;
 RECT 11.335 0.385 11.475 0.88 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.79 1.475 5.12 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.35 1.16 10.68 1.49 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.695 1.295 18.05 1.535 ;
 RECT 17.9 0.905 18.04 1.295 ;
 RECT 18.905 1.84 19.045 1.885 ;
 RECT 18.905 0.915 19.045 1.7 ;
 RECT 17.9 1.7 19.045 1.84 ;
 RECT 17.9 1.535 18.04 1.7 ;
 RECT 17.9 1.84 18.04 1.885 ;
 END
 ANTENNADIFFAREA 0.657 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 29.44 2.96 ;
 RECT 1.36 2.005 1.5 2.8 ;
 RECT 0.385 1.74 0.525 2.8 ;
 RECT 5.415 2.34 5.665 2.8 ;
 RECT 3.27 2.03 3.41 2.8 ;
 RECT 4.74 1.98 4.88 2.8 ;
 RECT 8.67 2.07 8.81 2.8 ;
 RECT 10.77 2.375 10.91 2.8 ;
 RECT 15.42 2.57 15.56 2.8 ;
 RECT 16.32 2.57 16.46 2.8 ;
 RECT 18.305 2.57 18.445 2.8 ;
 RECT 19.885 2.57 20.025 2.8 ;
 RECT 20.94 2.57 21.08 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 29.44 0.08 ;
 RECT 10.895 0.585 11.17 0.725 ;
 RECT 18.335 0.28 18.6 0.44 ;
 RECT 1.36 0.08 1.5 0.97 ;
 RECT 0.35 0.08 0.49 0.775 ;
 RECT 4.74 0.08 4.88 1.055 ;
 RECT 3.27 0.08 3.41 0.78 ;
 RECT 5.485 0.08 5.625 0.39 ;
 RECT 8.085 0.08 8.32 0.595 ;
 RECT 14.82 0.08 14.96 0.945 ;
 RECT 16.325 0.08 16.465 0.525 ;
 RECT 19.97 0.08 20.11 0.82 ;
 RECT 23.94 0.08 24.08 0.355 ;
 RECT 20.94 0.08 21.08 0.82 ;
 RECT 26.29 0.08 26.53 0.255 ;
 RECT 25.155 0.08 25.295 0.345 ;
 RECT 10.96 0.08 11.1 0.585 ;
 RECT 18.39 0.08 18.53 0.28 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.33 1.155 2.75 1.415 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.18 1.475 1.705 1.75 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.965 1.13 2.105 1.48 ;
 RECT 1.87 1.63 2.815 1.79 ;
 RECT 1.87 1.48 2.115 1.63 ;
 RECT 2.665 1.79 2.805 1.845 ;
 RECT 2.665 1.57 2.805 1.63 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.62 0.585 22.99 0.885 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 27.85 1.43 28.19 1.795 ;
 RECT 26.17 1.985 28.035 2.125 ;
 RECT 23.94 2.215 26.31 2.355 ;
 RECT 26.17 1.43 26.31 1.985 ;
 RECT 27.895 1.795 28.035 1.985 ;
 RECT 23.94 1.385 24.08 2.215 ;
 RECT 25.325 1.365 25.465 2.215 ;
 RECT 26.17 2.125 26.31 2.215 ;
 END
 END VDDG

 OBS
 LAYER PO ;
 RECT 25.78 0.375 26.01 0.43 ;
 RECT 24.995 0.93 25.225 0.955 ;
 RECT 24.995 1.055 25.225 1.14 ;
 RECT 24.995 0.955 25.515 1.055 ;
 RECT 23.725 0.205 23.825 0.755 ;
 RECT 23.725 0.855 23.825 2.195 ;
 RECT 26.59 1.12 26.69 2.195 ;
 RECT 22.76 0.755 24.295 0.835 ;
 RECT 22.76 0.835 24.29 0.855 ;
 RECT 24.195 0.21 24.295 0.755 ;
 RECT 22.76 0.59 22.99 0.755 ;
 RECT 23.725 2.195 26.69 2.295 ;
 RECT 11.615 2.69 13.265 2.695 ;
 RECT 13.09 2.54 13.265 2.69 ;
 RECT 12.405 2.695 13.265 2.79 ;
 RECT 11.615 0.655 11.715 2.595 ;
 RECT 11.615 2.595 12.505 2.69 ;
 RECT 13.09 2.33 13.32 2.54 ;
 RECT 15.675 0.81 15.775 2.21 ;
 RECT 15.635 0.6 15.865 0.81 ;
 RECT 9.4 1.575 9.5 2.485 ;
 RECT 9.91 1.41 10.14 1.475 ;
 RECT 9.91 1.575 10.14 1.62 ;
 RECT 9.4 1.475 10.14 1.575 ;
 RECT 10.325 1.45 10.425 1.655 ;
 RECT 10.325 1.755 10.425 2.57 ;
 RECT 10.325 0.655 10.425 1.13 ;
 RECT 10.325 1.23 10.425 1.24 ;
 RECT 9.41 0.66 9.51 1.13 ;
 RECT 10.325 1.655 11.285 1.755 ;
 RECT 11.185 1.755 11.285 2.355 ;
 RECT 10.325 1.24 10.58 1.45 ;
 RECT 9.41 1.13 10.425 1.23 ;
 RECT 17.155 0.29 18.265 0.39 ;
 RECT 18.165 0.39 18.265 1.4 ;
 RECT 18.165 1.5 18.265 2.385 ;
 RECT 18.655 0.505 18.755 1.4 ;
 RECT 18.655 1.5 18.755 2.385 ;
 RECT 17.155 0.225 17.385 0.29 ;
 RECT 17.155 0.39 17.385 0.435 ;
 RECT 18.165 1.4 18.755 1.5 ;
 RECT 15.205 0.835 15.305 2.21 ;
 RECT 15.205 0.47 15.37 0.625 ;
 RECT 14.32 0.455 15.37 0.47 ;
 RECT 14.32 0.47 14.55 0.665 ;
 RECT 14.43 0.37 15.37 0.455 ;
 RECT 15.205 0.625 15.435 0.835 ;
 RECT 16.575 1.635 16.675 1.66 ;
 RECT 16.575 1.66 16.83 1.87 ;
 RECT 16.575 1.87 16.675 2.565 ;
 RECT 12.945 0.885 13.175 0.925 ;
 RECT 12.945 0.925 13.79 1.025 ;
 RECT 12.945 1.025 13.175 1.095 ;
 RECT 13.625 0.795 13.79 0.925 ;
 RECT 13.625 0.585 13.855 0.795 ;
 RECT 5.775 1.62 5.875 2.69 ;
 RECT 5.84 0.185 12.75 0.19 ;
 RECT 5.84 0.19 7.995 0.285 ;
 RECT 5.84 0.285 5.94 1.52 ;
 RECT 12.65 1.29 13.67 1.39 ;
 RECT 12.65 0.19 12.75 1.29 ;
 RECT 6.66 1.565 6.76 2.69 ;
 RECT 5.34 1.44 5.585 1.52 ;
 RECT 5.34 1.62 5.585 1.69 ;
 RECT 5.34 1.52 5.94 1.62 ;
 RECT 7.895 0.285 7.995 1.24 ;
 RECT 7.895 0.09 12.75 0.185 ;
 RECT 13.44 1.285 13.67 1.29 ;
 RECT 13.44 1.39 13.67 1.615 ;
 RECT 5.775 2.69 6.76 2.79 ;
 RECT 8.945 0.47 9.13 0.5 ;
 RECT 16.58 0.19 16.68 1.18 ;
 RECT 14.04 0.09 16.68 0.19 ;
 RECT 14.04 0.19 14.14 1.795 ;
 RECT 13.155 1.71 13.255 1.795 ;
 RECT 13.155 1.895 13.255 1.905 ;
 RECT 14.04 1.895 14.14 1.91 ;
 RECT 12.135 1.61 13.255 1.71 ;
 RECT 12.135 0.47 12.235 1.61 ;
 RECT 12.685 1.71 12.785 2.445 ;
 RECT 13.155 1.795 14.14 1.895 ;
 RECT 8.945 0.37 12.235 0.47 ;
 RECT 8.9 0.5 9.13 0.71 ;
 RECT 16.85 1.25 17.11 1.3 ;
 RECT 17.01 0.61 17.11 1.25 ;
 RECT 16.85 1.4 17.11 1.46 ;
 RECT 17.01 1.46 17.11 2.56 ;
 RECT 17.54 0.84 17.64 1.3 ;
 RECT 16.85 1.3 17.64 1.4 ;
 RECT 17.525 0.63 17.755 0.84 ;
 RECT 2.755 1.82 2.855 2.735 ;
 RECT 2.615 1.59 2.855 1.82 ;
 RECT 1.95 0.555 2.05 1.145 ;
 RECT 1.91 1.145 2.155 1.385 ;
 RECT 3.525 0.335 3.625 1.155 ;
 RECT 3.525 1.365 3.625 2.745 ;
 RECT 3.335 1.155 3.625 1.365 ;
 RECT 2.335 1.41 2.435 1.645 ;
 RECT 2.565 0.555 2.665 1.18 ;
 RECT 2.285 1.745 2.385 2.735 ;
 RECT 2.285 1.645 2.435 1.745 ;
 RECT 2.335 1.18 2.665 1.41 ;
 RECT 5 0.57 5.1 1.495 ;
 RECT 4.805 1.495 5.1 1.745 ;
 RECT 5 1.745 5.1 2.37 ;
 RECT 7.155 1.33 7.295 1.475 ;
 RECT 7.155 1.71 7.255 2.475 ;
 RECT 7.195 0.65 7.295 1.33 ;
 RECT 7.155 1.475 7.385 1.71 ;
 RECT 2.85 0.175 3.155 0.405 ;
 RECT 3.055 0.405 3.155 2.735 ;
 RECT 1.145 1.475 1.715 1.75 ;
 RECT 1.615 0.555 1.715 1.475 ;
 RECT 1.615 1.75 1.715 2.735 ;
 RECT 1.145 0.555 1.245 1.475 ;
 RECT 1.145 1.75 1.245 2.685 ;
 RECT 7.595 0.715 7.695 1.61 ;
 RECT 7.63 1.71 7.73 2.48 ;
 RECT 7.595 1.61 7.73 1.71 ;
 RECT 7.475 0.485 7.715 0.715 ;
 RECT 4.285 0.27 4.625 0.52 ;
 RECT 4.525 0.52 4.625 2.465 ;
 RECT 11.22 0.655 11.32 1.24 ;
 RECT 11.09 1.24 11.32 1.475 ;
 RECT 8.76 1.61 9.025 1.82 ;
 RECT 8.925 1.82 9.025 2.49 ;
 RECT 8.555 0.66 8.655 1.51 ;
 RECT 8.555 1.51 9.025 1.61 ;
 RECT 8.24 2.465 8.555 2.71 ;
 RECT 8.455 1.79 8.555 2.465 ;
 RECT 6.705 0.705 6.805 1.165 ;
 RECT 6.265 1.27 6.365 1.445 ;
 RECT 6.705 0.47 6.99 0.705 ;
 RECT 6.265 1.17 6.805 1.265 ;
 RECT 6.495 1.165 6.805 1.17 ;
 RECT 6.265 1.265 6.64 1.27 ;
 RECT 6.12 1.445 6.365 1.69 ;
 RECT 27.6 0.19 27.7 2.66 ;
 RECT 26.59 0.09 27.7 0.19 ;
 RECT 22.965 1.25 23.065 2.66 ;
 RECT 22.965 1.195 23.25 1.25 ;
 RECT 26.59 0.19 26.69 0.94 ;
 RECT 23.02 1.04 23.25 1.095 ;
 RECT 22.965 2.66 27.7 2.76 ;
 RECT 22.965 1.095 23.295 1.195 ;
 RECT 24.2 1.245 24.3 2.015 ;
 RECT 24.07 1.035 24.3 1.245 ;
 RECT 24.505 0.21 24.605 0.99 ;
 RECT 24.505 0.99 24.745 1.2 ;
 RECT 24.505 1.2 24.605 1.995 ;
 RECT 20.25 0.385 20.35 1.285 ;
 RECT 20.25 1.385 20.35 2.585 ;
 RECT 19.67 0.385 19.77 1.2 ;
 RECT 19.655 1.285 21.295 1.385 ;
 RECT 21.195 0.19 21.295 1.285 ;
 RECT 22.18 0.19 22.28 0.22 ;
 RECT 19.67 1.435 19.77 2.585 ;
 RECT 19.655 1.2 19.865 1.285 ;
 RECT 19.655 1.385 19.865 1.435 ;
 RECT 20.725 0.385 20.825 1.285 ;
 RECT 20.725 1.385 20.825 2.585 ;
 RECT 21.195 1.385 21.295 2.585 ;
 RECT 21.195 0.09 22.28 0.19 ;
 RECT 22.18 0.22 22.41 0.43 ;
 RECT 26.9 2.265 27.185 2.475 ;
 RECT 26.9 1.195 27 2.265 ;
 RECT 26.9 0.37 27 0.985 ;
 RECT 26.9 0.985 27.15 1.195 ;
 RECT 25.415 1.055 25.515 1.135 ;
 RECT 25.415 0.375 25.515 0.955 ;
 RECT 25.415 1.135 25.685 1.235 ;
 RECT 25.585 1.235 25.685 1.835 ;
 RECT 25.78 0.22 26.01 0.275 ;
 RECT 25.415 0.275 26.01 0.375 ;
 LAYER CO ;
 RECT 7.855 1.825 7.985 1.955 ;
 RECT 8.205 2.125 8.335 2.255 ;
 RECT 4.275 2.115 4.405 2.245 ;
 RECT 0.355 0.59 0.485 0.72 ;
 RECT 11.875 1.945 12.005 2.075 ;
 RECT 10.075 0.88 10.205 1.01 ;
 RECT 5.4 1.495 5.53 1.625 ;
 RECT 19.89 2.64 20.02 2.77 ;
 RECT 7.53 0.53 7.66 0.66 ;
 RECT 11.14 1.28 11.27 1.41 ;
 RECT 17.905 1.705 18.035 1.835 ;
 RECT 5.22 1.995 5.35 2.125 ;
 RECT 20.475 1.71 20.605 1.84 ;
 RECT 16.33 0.33 16.46 0.46 ;
 RECT 18.91 1.705 19.04 1.835 ;
 RECT 12.905 0.595 13.035 0.725 ;
 RECT 17.23 1.78 17.36 1.91 ;
 RECT 18.395 0.305 18.525 0.435 ;
 RECT 19.975 0.62 20.105 0.75 ;
 RECT 6.905 2.07 7.035 2.2 ;
 RECT 23.07 1.08 23.2 1.21 ;
 RECT 24.12 1.075 24.25 1.205 ;
 RECT 24.565 1.03 24.695 1.16 ;
 RECT 27.005 2.305 27.135 2.435 ;
 RECT 22.23 0.26 22.36 0.39 ;
 RECT 25.83 0.26 25.96 0.39 ;
 RECT 26.97 1.025 27.1 1.155 ;
 RECT 25.045 0.97 25.175 1.1 ;
 RECT 22.81 0.63 22.94 0.76 ;
 RECT 15.255 0.665 15.385 0.795 ;
 RECT 13.14 2.37 13.27 2.5 ;
 RECT 15.685 0.64 15.815 0.77 ;
 RECT 9.96 1.45 10.09 1.58 ;
 RECT 10.4 1.28 10.53 1.41 ;
 RECT 12.995 0.925 13.125 1.055 ;
 RECT 17.205 0.265 17.335 0.395 ;
 RECT 17.575 0.67 17.705 0.8 ;
 RECT 14.37 0.495 14.5 0.625 ;
 RECT 16.65 1.7 16.78 1.83 ;
 RECT 13.675 0.625 13.805 0.755 ;
 RECT 13.49 1.445 13.62 1.575 ;
 RECT 8.95 0.54 9.08 0.67 ;
 RECT 16.9 1.29 17.03 1.42 ;
 RECT 2.505 2.115 2.635 2.245 ;
 RECT 1.365 2.055 1.495 2.185 ;
 RECT 0.895 2.055 1.025 2.185 ;
 RECT 3.745 1.79 3.875 1.92 ;
 RECT 1.97 1.195 2.1 1.325 ;
 RECT 3.385 1.195 3.515 1.325 ;
 RECT 2.9 0.225 3.03 0.355 ;
 RECT 0.895 0.775 1.025 0.905 ;
 RECT 3.745 0.775 3.875 0.905 ;
 RECT 3.275 0.585 3.405 0.715 ;
 RECT 2.31 0.775 2.44 0.905 ;
 RECT 17.905 0.975 18.035 1.105 ;
 RECT 5.49 0.21 5.62 0.34 ;
 RECT 18.31 2.64 18.44 2.77 ;
 RECT 9.145 2.015 9.275 2.145 ;
 RECT 7.375 2.125 7.505 2.255 ;
 RECT 14.955 1.7 15.085 1.83 ;
 RECT 5.485 2.345 5.615 2.475 ;
 RECT 19.695 1.25 19.825 1.38 ;
 RECT 0.355 0.33 0.485 0.46 ;
 RECT 25.33 1.44 25.46 1.57 ;
 RECT 26.175 1.485 26.305 1.615 ;
 RECT 27.12 1.46 27.25 1.59 ;
 RECT 23.945 1.47 24.075 1.6 ;
 RECT 23.475 1.42 23.605 1.55 ;
 RECT 25.805 1.4 25.935 1.53 ;
 RECT 25.16 0.115 25.29 0.245 ;
 RECT 23.945 0.13 24.075 0.26 ;
 RECT 27.9 1.47 28.03 1.6 ;
 RECT 26.34 0.115 26.47 0.245 ;
 RECT 25.665 0.59 25.795 0.72 ;
 RECT 23.225 0.505 23.355 0.635 ;
 RECT 24.725 1.48 24.855 1.61 ;
 RECT 24.725 0.43 24.855 0.56 ;
 RECT 27.12 0.59 27.25 0.72 ;
 RECT 16.325 2.64 16.455 2.77 ;
 RECT 0.39 2.085 0.52 2.215 ;
 RECT 10.775 2.445 10.905 2.575 ;
 RECT 4.275 0.79 4.405 0.92 ;
 RECT 15.425 2.64 15.555 2.77 ;
 RECT 18.91 0.975 19.04 1.105 ;
 RECT 0.39 1.825 0.52 1.955 ;
 RECT 15.895 1.705 16.025 1.835 ;
 RECT 6.81 0.525 6.94 0.655 ;
 RECT 6.455 0.88 6.585 1.01 ;
 RECT 19.415 0.62 19.545 0.75 ;
 RECT 8.28 2.515 8.41 2.645 ;
 RECT 8.135 0.455 8.265 0.585 ;
 RECT 6.06 0.905 6.19 1.035 ;
 RECT 17.23 0.83 17.36 0.96 ;
 RECT 20.475 0.63 20.605 0.76 ;
 RECT 14.825 0.745 14.955 0.875 ;
 RECT 4.745 2.05 4.875 2.18 ;
 RECT 10.965 0.59 11.095 0.72 ;
 RECT 6.41 2.105 6.54 2.235 ;
 RECT 9.63 2.07 9.76 2.2 ;
 RECT 8.675 2.135 8.805 2.265 ;
 RECT 8.815 1.63 8.945 1.76 ;
 RECT 19.415 1.725 19.545 1.855 ;
 RECT 5.35 0.88 5.48 1.01 ;
 RECT 9.63 0.88 9.76 1.01 ;
 RECT 15.93 0.96 16.06 1.09 ;
 RECT 0.39 2.345 0.52 2.475 ;
 RECT 4.745 0.79 4.875 0.92 ;
 RECT 9.145 0.93 9.275 1.06 ;
 RECT 11.875 0.875 12.005 1.005 ;
 RECT 7.205 1.525 7.335 1.655 ;
 RECT 4.345 0.325 4.475 0.455 ;
 RECT 21.415 1.71 21.545 1.84 ;
 RECT 20.945 0.62 21.075 0.75 ;
 RECT 20.945 2.64 21.075 2.77 ;
 RECT 3.745 2.05 3.875 2.18 ;
 RECT 1.37 1.55 1.5 1.68 ;
 RECT 3.275 2.09 3.405 2.22 ;
 RECT 2.49 1.23 2.62 1.36 ;
 RECT 1.365 2.315 1.495 2.445 ;
 RECT 2.67 1.64 2.8 1.77 ;
 RECT 1.365 0.775 1.495 0.905 ;
 RECT 3.275 2.35 3.405 2.48 ;
 RECT 21.415 0.63 21.545 0.76 ;
 RECT 12.905 1.87 13.035 2 ;
 RECT 4.865 1.55 4.995 1.68 ;
 RECT 6.925 0.88 7.055 1.01 ;
 RECT 12.4 0.595 12.53 0.725 ;
 RECT 10.075 1.995 10.205 2.125 ;
 RECT 5.995 1.825 6.125 1.955 ;
 RECT 6.175 1.49 6.305 1.62 ;
 RECT 12.4 1.9 12.53 2.03 ;
 LAYER M1 ;
 RECT 8.76 1.79 9 1.835 ;
 RECT 8.185 1.65 9 1.79 ;
 RECT 10.07 1.62 10.21 1.735 ;
 RECT 10.07 1.875 10.21 2.18 ;
 RECT 10.07 0.81 10.21 1.41 ;
 RECT 9.91 1.41 10.21 1.62 ;
 RECT 11.135 1.415 11.275 1.735 ;
 RECT 10.07 1.735 11.275 1.875 ;
 RECT 11.075 1.275 11.34 1.415 ;
 RECT 2.96 0.91 3.1 1.19 ;
 RECT 2.96 1.33 3.1 2.11 ;
 RECT 2.255 0.77 3.1 0.91 ;
 RECT 2.45 2.11 3.1 2.25 ;
 RECT 2.96 1.19 3.52 1.33 ;
 RECT 3.38 1.145 3.52 1.19 ;
 RECT 3.38 1.33 3.52 1.375 ;
 RECT 5.26 1.63 5.4 1.99 ;
 RECT 5.26 1.475 5.605 1.63 ;
 RECT 5.345 0.81 5.485 1.475 ;
 RECT 5.15 1.99 5.4 2.13 ;
 RECT 25.78 0.285 26.15 0.43 ;
 RECT 26.01 0.43 26.15 0.705 ;
 RECT 25.78 0.22 26.01 0.285 ;
 RECT 27.43 0.845 27.57 1.38 ;
 RECT 27.115 1.52 27.255 1.725 ;
 RECT 26.01 0.705 27.57 0.845 ;
 RECT 27.115 0.505 27.255 0.705 ;
 RECT 27.115 1.38 27.57 1.52 ;
 RECT 25.04 1.14 25.18 1.34 ;
 RECT 24.72 1.48 24.86 1.755 ;
 RECT 25.04 0.725 25.18 0.93 ;
 RECT 24.72 0.35 24.86 0.585 ;
 RECT 24.72 1.34 25.18 1.48 ;
 RECT 24.995 0.93 25.225 1.14 ;
 RECT 24.72 0.585 25.18 0.725 ;
 RECT 23.02 1.22 23.25 1.25 ;
 RECT 23.02 1.19 23.61 1.22 ;
 RECT 23.16 1.01 23.47 1.04 ;
 RECT 23.02 1.04 23.47 1.05 ;
 RECT 23.295 0.64 23.435 1.01 ;
 RECT 23.47 1.22 23.61 1.745 ;
 RECT 23.175 0.5 23.435 0.64 ;
 RECT 24.07 1.035 24.3 1.05 ;
 RECT 24.07 1.19 24.3 1.245 ;
 RECT 23.02 1.05 24.3 1.19 ;
 RECT 22.18 0.36 22.41 0.43 ;
 RECT 23.575 0.36 23.715 0.56 ;
 RECT 22.18 0.22 23.715 0.36 ;
 RECT 24.315 0.7 24.455 0.745 ;
 RECT 24.44 0.99 24.745 1.2 ;
 RECT 24.44 0.885 24.58 0.99 ;
 RECT 24.315 0.745 24.58 0.885 ;
 RECT 23.575 0.56 24.455 0.7 ;
 RECT 17.525 0.72 17.755 0.84 ;
 RECT 17.52 0.58 18.94 0.72 ;
 RECT 18.8 0.37 18.94 0.58 ;
 RECT 19.69 0.37 19.83 1.46 ;
 RECT 18.8 0.23 19.83 0.37 ;
 RECT 12.9 0.525 13.04 0.885 ;
 RECT 12.9 1.095 13.04 2.065 ;
 RECT 12.9 0.885 13.175 1.095 ;
 RECT 9.625 0.82 9.765 2.33 ;
 RECT 9.625 2.47 9.765 2.475 ;
 RECT 10.475 2.165 10.615 2.33 ;
 RECT 10.475 2.47 10.615 2.475 ;
 RECT 9.625 2.33 10.615 2.47 ;
 RECT 11.555 2.165 11.695 2.295 ;
 RECT 11.87 0.765 12.01 2.295 ;
 RECT 11.87 2.435 12.01 2.44 ;
 RECT 12.395 0.525 12.535 2.295 ;
 RECT 12.395 2.435 12.535 2.44 ;
 RECT 10.475 2.025 11.695 2.165 ;
 RECT 11.555 2.295 12.535 2.435 ;
 RECT 15.205 0.36 15.435 0.835 ;
 RECT 16.005 0.36 16.145 0.665 ;
 RECT 15.205 0.22 16.15 0.36 ;
 RECT 17.225 0.22 17.365 0.225 ;
 RECT 17.225 0.435 17.365 0.665 ;
 RECT 16.005 0.665 17.365 0.805 ;
 RECT 17.225 0.805 17.365 1.98 ;
 RECT 17.155 0.225 17.385 0.435 ;
 RECT 13.625 0.585 14.55 0.63 ;
 RECT 13.625 0.63 13.855 0.795 ;
 RECT 13.65 0.49 14.55 0.585 ;
 RECT 14.32 0.455 14.55 0.49 ;
 RECT 14.32 0.63 14.55 0.665 ;
 RECT 6.74 0.52 7.34 0.66 ;
 RECT 7.2 0.66 7.34 1.015 ;
 RECT 8.745 0.505 9.13 0.71 ;
 RECT 7.2 1.015 8.885 1.155 ;
 RECT 8.745 0.71 8.885 1.015 ;
 RECT 8.9 0.5 9.13 0.505 ;
 RECT 6.055 1.67 6.195 1.82 ;
 RECT 6.055 1.96 6.195 2.51 ;
 RECT 6.055 0.5 6.195 1.44 ;
 RECT 6.055 1.44 6.31 1.67 ;
 RECT 5.925 1.82 6.195 1.96 ;
 RECT 6.055 2.51 8.53 2.65 ;
 RECT 4.05 1.335 4.19 2.11 ;
 RECT 4.05 2.25 4.19 2.255 ;
 RECT 4.05 0.925 4.19 1.195 ;
 RECT 4.05 2.11 4.475 2.25 ;
 RECT 4.05 0.785 4.475 0.925 ;
 RECT 4.05 1.195 5.16 1.335 ;
 RECT 5.02 0.67 5.16 1.195 ;
 RECT 6.45 0.36 6.59 2.035 ;
 RECT 5.765 0.22 6.59 0.36 ;
 RECT 6.405 2.17 6.545 2.305 ;
 RECT 6.405 2.035 6.59 2.17 ;
 RECT 5.02 0.53 5.905 0.67 ;
 RECT 5.765 0.36 5.905 0.53 ;
 RECT 3.74 0.57 3.88 2.25 ;
 RECT 4.235 0.22 4.6 0.43 ;
 RECT 4.235 0.57 4.6 0.615 ;
 RECT 3.74 0.43 4.6 0.57 ;
 RECT 0.89 0.72 1.03 1.195 ;
 RECT 0.89 1.335 1.03 2.27 ;
 RECT 0.89 1.195 1.815 1.335 ;
 RECT 1.675 0.36 1.815 1.195 ;
 RECT 1.675 0.22 3.1 0.36 ;
 RECT 13.09 2.42 13.32 2.54 ;
 RECT 22.615 2.42 22.755 2.515 ;
 RECT 22.615 2.275 22.755 2.28 ;
 RECT 13.09 2.28 22.755 2.42 ;
 RECT 26.955 2.475 27.095 2.515 ;
 RECT 22.615 2.515 27.095 2.655 ;
 RECT 26.955 2.265 27.185 2.475 ;
 RECT 25.8 1.175 25.94 1.6 ;
 RECT 25.66 0.725 25.8 1.035 ;
 RECT 25.595 0.585 25.87 0.725 ;
 RECT 26.92 0.985 27.15 1.035 ;
 RECT 26.92 1.175 27.15 1.195 ;
 RECT 25.66 1.035 27.15 1.175 ;
 RECT 14.95 1.51 15.09 1.695 ;
 RECT 14.88 1.695 15.16 1.835 ;
 RECT 15.89 1.51 16.03 1.7 ;
 RECT 15.925 1.095 16.065 1.37 ;
 RECT 16.85 1.25 17.08 1.37 ;
 RECT 14.95 1.37 17.08 1.51 ;
 RECT 15.825 1.7 16.1 1.84 ;
 RECT 15.855 0.955 16.135 1.095 ;
 RECT 13.435 2.05 13.575 2.055 ;
 RECT 13.43 1.915 14.735 1.985 ;
 RECT 13.43 1.91 14.73 1.915 ;
 RECT 13.435 1.615 13.575 1.91 ;
 RECT 16.6 1.87 16.785 1.985 ;
 RECT 13.43 1.985 16.785 2.05 ;
 RECT 14.59 2.05 16.785 2.125 ;
 RECT 13.435 1.43 13.67 1.615 ;
 RECT 13.44 1.405 13.67 1.43 ;
 RECT 16.6 1.66 16.83 1.87 ;
 RECT 7.305 2.12 8.405 2.26 ;
 RECT 7.135 1.52 8.005 1.66 ;
 RECT 7.865 1.44 8.005 1.52 ;
 RECT 9.14 0.865 9.28 1.3 ;
 RECT 9.14 1.44 9.28 2.215 ;
 RECT 7.865 1.3 9.28 1.44 ;
 RECT 6.745 1.22 7.06 1.36 ;
 RECT 6.92 0.805 7.06 1.22 ;
 RECT 6.83 1.96 7.11 2.215 ;
 RECT 6.745 1.36 6.885 1.82 ;
 RECT 6.745 1.82 8.325 1.96 ;
 RECT 8.185 1.79 8.325 1.82 ;
 RECT 8.76 1.58 9 1.65 ;
 END
END RSDFFNSRARX2

MACRO RSDFFNSRASRNX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 29.44 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.695 0.59 23.065 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 27.925 1.435 28.265 1.8 ;
 RECT 26.245 1.99 28.11 2.13 ;
 RECT 24.015 2.22 26.385 2.36 ;
 RECT 26.245 1.435 26.385 1.99 ;
 RECT 27.97 1.8 28.11 1.99 ;
 RECT 24.015 1.39 24.155 2.22 ;
 RECT 25.4 1.37 25.54 2.22 ;
 RECT 26.245 2.13 26.385 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 5.155 0.08 5.435 0.295 ;
 RECT 9.085 0.31 9.375 0.45 ;
 RECT 12.77 0.59 13.04 0.73 ;
 RECT 16.695 0.275 17.72 0.415 ;
 RECT 21.055 0.475 21.32 0.635 ;
 RECT 26.365 0.08 26.605 0.26 ;
 RECT 17.58 0.75 18.525 0.89 ;
 RECT 0.31 0.08 0.45 0.775 ;
 RECT 1.28 0.08 1.42 0.93 ;
 RECT 4.635 0.08 4.775 0.97 ;
 RECT 3.19 0.08 3.33 0.74 ;
 RECT 7.98 0.08 8.215 0.46 ;
 RECT 24.015 0.08 24.155 0.36 ;
 RECT 25.23 0.08 25.37 0.35 ;
 RECT 0 -0.08 29.44 0.08 ;
 RECT 9.165 0.08 9.305 0.31 ;
 RECT 12.835 0.08 12.975 0.59 ;
 RECT 16.695 0.415 16.835 0.945 ;
 RECT 16.695 0.08 16.835 0.275 ;
 RECT 21.11 0.635 21.25 0.715 ;
 RECT 21.11 0.08 21.25 0.475 ;
 RECT 18.385 0.89 18.525 1.11 ;
 RECT 17.58 0.415 17.72 0.75 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.62 1.2 20.91 1.44 ;
 RECT 20.62 0.915 20.76 1.2 ;
 RECT 21.625 1.84 21.765 1.885 ;
 RECT 21.625 0.915 21.765 1.7 ;
 RECT 20.62 1.84 20.76 1.885 ;
 RECT 20.62 1.7 21.765 1.84 ;
 RECT 20.62 1.44 20.76 1.7 ;
 END
 ANTENNADIFFAREA 0.479 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 29.44 2.96 ;
 RECT 20.965 2.6 21.23 2.8 ;
 RECT 12.58 2.215 12.855 2.355 ;
 RECT 1.28 1.965 1.42 2.8 ;
 RECT 0.31 1.74 0.45 2.8 ;
 RECT 5.31 2.34 5.56 2.8 ;
 RECT 4.635 1.98 4.775 2.8 ;
 RECT 3.19 1.99 3.33 2.8 ;
 RECT 8.685 2.07 8.825 2.8 ;
 RECT 10.195 2.225 10.335 2.8 ;
 RECT 9.165 2.19 9.305 2.8 ;
 RECT 15.605 2.335 15.875 2.8 ;
 RECT 12.645 2.355 12.785 2.8 ;
 RECT 12.645 2.195 12.785 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.685 1.475 5.015 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.225 1.16 12.6 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.375 0.485 7.69 0.605 ;
 RECT 12.295 0.87 13.35 1.01 ;
 RECT 12.295 0.745 12.435 0.87 ;
 RECT 13.205 0.245 15.355 0.255 ;
 RECT 13.205 0.255 15.36 0.385 ;
 RECT 15.22 1.09 17.21 1.23 ;
 RECT 17.415 1.56 17.645 1.6 ;
 RECT 17.07 1.42 17.645 1.56 ;
 RECT 17.415 1.39 17.645 1.42 ;
 RECT 7.375 0.605 12.435 0.745 ;
 RECT 13.21 0.385 13.35 0.87 ;
 RECT 15.22 0.385 15.36 1.09 ;
 RECT 17.07 1.23 17.21 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.985 1.79 10.425 2.075 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.1 1.435 1.625 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.78 1.59 2.735 1.75 ;
 RECT 1.885 1.09 2.025 1.44 ;
 RECT 1.78 1.44 2.025 1.59 ;
 RECT 2.585 1.75 2.725 1.805 ;
 RECT 2.585 1.53 2.725 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.25 1.115 2.67 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 OBS
 LAYER PO ;
 RECT 24.145 1.035 24.375 1.245 ;
 RECT 15.915 0.105 18.74 0.205 ;
 RECT 15.915 0.205 16.015 1.91 ;
 RECT 18.64 0.205 18.74 1.265 ;
 RECT 15.095 1.71 15.195 1.91 ;
 RECT 14.01 1.61 15.195 1.71 ;
 RECT 14.01 0.475 14.11 1.61 ;
 RECT 14.56 1.71 14.66 2.425 ;
 RECT 10.675 0.475 10.775 0.895 ;
 RECT 15.095 1.91 16.015 2.01 ;
 RECT 10.675 0.375 14.11 0.475 ;
 RECT 10.55 0.895 10.78 1.105 ;
 RECT 16.225 0.455 18.155 0.535 ;
 RECT 17.925 0.535 18.155 0.6 ;
 RECT 17.925 0.39 18.155 0.435 ;
 RECT 16.305 0.435 18.155 0.455 ;
 RECT 16.225 0.535 16.455 0.665 ;
 RECT 17.08 0.535 17.31 0.835 ;
 RECT 17.08 0.835 17.18 2.39 ;
 RECT 24.58 0.215 24.68 0.995 ;
 RECT 24.58 0.995 24.82 1.205 ;
 RECT 24.58 1.205 24.68 2 ;
 RECT 26.975 0.375 27.075 0.99 ;
 RECT 26.975 0.99 27.225 1.2 ;
 RECT 26.975 1.2 27.075 2.27 ;
 RECT 26.975 2.27 27.26 2.48 ;
 RECT 13.49 0.655 13.59 2.305 ;
 RECT 13.795 2.3 14.025 2.305 ;
 RECT 13.795 2.405 14.025 2.51 ;
 RECT 13.49 2.305 14.025 2.405 ;
 RECT 23.8 0.21 23.9 0.755 ;
 RECT 23.8 0.855 23.9 2.2 ;
 RECT 26.665 1.125 26.765 2.2 ;
 RECT 22.835 0.755 24.37 0.84 ;
 RECT 22.835 0.84 24.365 0.855 ;
 RECT 24.27 0.215 24.37 0.755 ;
 RECT 22.835 0.595 23.065 0.755 ;
 RECT 23.8 2.2 26.765 2.3 ;
 RECT 12.2 1.28 12.455 1.45 ;
 RECT 12.2 1.45 12.3 1.655 ;
 RECT 12.2 0.655 12.3 1.18 ;
 RECT 12.2 1.655 13.16 1.755 ;
 RECT 13.06 1.755 13.16 2.355 ;
 RECT 11.285 0.66 11.385 1.18 ;
 RECT 12.2 1.755 12.3 2.51 ;
 RECT 11.285 1.24 12.455 1.28 ;
 RECT 11.285 1.18 12.3 1.24 ;
 RECT 25.49 0.38 25.59 0.96 ;
 RECT 25.49 1.06 25.59 1.14 ;
 RECT 25.07 0.935 25.3 0.96 ;
 RECT 25.07 0.96 25.59 1.06 ;
 RECT 25.07 1.06 25.3 1.145 ;
 RECT 25.49 1.14 25.76 1.24 ;
 RECT 25.66 1.24 25.76 1.84 ;
 RECT 25.855 0.22 26.085 0.28 ;
 RECT 25.855 0.38 26.085 0.43 ;
 RECT 25.49 0.28 26.085 0.38 ;
 RECT 11.275 1.575 11.375 2.485 ;
 RECT 11.785 1.575 12.015 1.685 ;
 RECT 11.275 1.475 12.015 1.575 ;
 RECT 27.675 0.195 27.775 2.665 ;
 RECT 26.665 0.095 27.775 0.195 ;
 RECT 23.04 1.245 23.14 2.665 ;
 RECT 26.665 0.195 26.765 0.945 ;
 RECT 23.04 1.2 23.325 1.245 ;
 RECT 23.095 1.035 23.325 1.1 ;
 RECT 23.04 2.665 27.775 2.765 ;
 RECT 23.04 1.1 23.37 1.2 ;
 RECT 15.5 0.795 15.665 0.925 ;
 RECT 14.82 0.885 15.05 0.925 ;
 RECT 14.82 1.025 15.05 1.095 ;
 RECT 14.82 0.925 15.665 1.025 ;
 RECT 15.5 0.585 15.73 0.795 ;
 RECT 13.095 0.655 13.195 1.24 ;
 RECT 12.965 1.24 13.195 1.475 ;
 RECT 4.895 0.49 4.995 1.495 ;
 RECT 4.7 1.495 4.995 1.745 ;
 RECT 4.895 1.745 4.995 2.37 ;
 RECT 7.49 0.715 7.59 1.61 ;
 RECT 7.525 1.71 7.625 2.48 ;
 RECT 7.49 1.61 7.625 1.71 ;
 RECT 7.37 0.485 7.61 0.715 ;
 RECT 7.05 1.33 7.19 1.475 ;
 RECT 7.05 1.71 7.15 2.475 ;
 RECT 7.09 0.65 7.19 1.33 ;
 RECT 7.05 1.475 7.28 1.71 ;
 RECT 4.18 0.27 4.52 0.52 ;
 RECT 4.42 0.52 4.52 2.465 ;
 RECT 1.87 0.515 1.97 1.105 ;
 RECT 1.83 1.105 2.075 1.345 ;
 RECT 6.6 0.705 6.7 1.165 ;
 RECT 6.16 1.27 6.26 1.445 ;
 RECT 6.6 0.47 6.885 0.705 ;
 RECT 6.16 1.17 6.7 1.265 ;
 RECT 6.39 1.165 6.7 1.17 ;
 RECT 6.16 1.265 6.535 1.27 ;
 RECT 6.015 1.445 6.26 1.69 ;
 RECT 1.065 1.435 1.635 1.71 ;
 RECT 1.535 0.515 1.635 1.435 ;
 RECT 1.535 1.71 1.635 2.695 ;
 RECT 1.065 0.515 1.165 1.435 ;
 RECT 1.065 1.71 1.165 2.645 ;
 RECT 2.535 1.55 2.775 1.78 ;
 RECT 2.675 1.78 2.775 2.695 ;
 RECT 2.255 1.37 2.355 1.605 ;
 RECT 2.485 0.515 2.585 1.14 ;
 RECT 2.205 1.705 2.305 2.695 ;
 RECT 2.205 1.605 2.355 1.705 ;
 RECT 2.255 1.14 2.585 1.37 ;
 RECT 2.975 0.135 3.075 0.22 ;
 RECT 2.815 0.22 3.075 0.43 ;
 RECT 2.975 0.43 3.075 2.695 ;
 RECT 3.445 0.295 3.545 1.115 ;
 RECT 3.28 1.115 3.545 1.325 ;
 RECT 3.445 1.325 3.545 2.74 ;
 RECT 20.885 1.52 20.985 2.255 ;
 RECT 20.105 1.42 21.475 1.455 ;
 RECT 20.885 1.4 21.475 1.42 ;
 RECT 20.885 0.67 20.985 1.4 ;
 RECT 20.115 1.455 21.475 1.5 ;
 RECT 20.115 1.5 20.985 1.52 ;
 RECT 21.375 0.675 21.475 1.4 ;
 RECT 21.375 1.5 21.475 2.26 ;
 RECT 20.105 1.245 20.335 1.42 ;
 RECT 8.31 2.445 8.57 2.655 ;
 RECT 8.47 1.79 8.57 2.445 ;
 RECT 18.58 1.445 18.68 2.035 ;
 RECT 18.565 2.035 18.795 2.245 ;
 RECT 19.05 0.55 19.15 2.69 ;
 RECT 9.98 2.015 10.08 2.69 ;
 RECT 9.98 1.58 10.08 1.805 ;
 RECT 9.72 1.01 9.82 1.48 ;
 RECT 9.98 1.805 10.215 2.015 ;
 RECT 9.98 2.69 19.15 2.79 ;
 RECT 9.72 1.48 10.08 1.58 ;
 RECT 9.42 1.005 9.52 1.615 ;
 RECT 9.28 1.615 9.52 1.825 ;
 RECT 9.42 1.825 9.52 2.69 ;
 RECT 19.52 0.55 19.71 0.56 ;
 RECT 19.61 0.325 19.71 0.55 ;
 RECT 19.52 0.77 19.62 2.155 ;
 RECT 19.52 0.56 19.775 0.77 ;
 RECT 22.055 0.22 22.285 0.225 ;
 RECT 22.055 0.325 22.285 0.43 ;
 RECT 19.61 0.225 22.285 0.325 ;
 RECT 17.55 0.73 17.65 1.39 ;
 RECT 17.415 1.39 17.65 1.6 ;
 RECT 17.55 1.6 17.65 2.39 ;
 RECT 5.735 0.285 5.835 1.52 ;
 RECT 5.235 1.52 5.835 1.62 ;
 RECT 5.735 0.185 14.625 0.195 ;
 RECT 7.79 0.095 14.625 0.185 ;
 RECT 5.735 0.195 7.89 0.285 ;
 RECT 14.525 0.195 14.625 1.29 ;
 RECT 15.42 1.39 15.615 1.405 ;
 RECT 6.555 1.565 6.655 2.675 ;
 RECT 5.67 1.62 5.77 2.675 ;
 RECT 5.235 1.44 5.48 1.52 ;
 RECT 5.235 1.62 5.48 1.69 ;
 RECT 7.79 0.285 7.89 1.24 ;
 RECT 14.525 1.29 15.615 1.39 ;
 RECT 5.67 2.675 6.655 2.775 ;
 RECT 15.42 1.405 15.65 1.615 ;
 RECT 24.275 1.245 24.375 2.02 ;
 LAYER CO ;
 RECT 25.74 0.595 25.87 0.725 ;
 RECT 3.195 0.545 3.325 0.675 ;
 RECT 27.195 0.595 27.325 0.725 ;
 RECT 14.275 0.595 14.405 0.725 ;
 RECT 5.115 1.995 5.245 2.125 ;
 RECT 13.75 1.945 13.88 2.075 ;
 RECT 6.35 0.88 6.48 1.01 ;
 RECT 0.815 2.015 0.945 2.145 ;
 RECT 2.865 0.26 2.995 0.39 ;
 RECT 3.33 1.155 3.46 1.285 ;
 RECT 20.155 1.285 20.285 1.415 ;
 RECT 17.975 0.43 18.105 0.56 ;
 RECT 19.595 0.6 19.725 0.73 ;
 RECT 8.36 2.485 8.49 2.615 ;
 RECT 18.615 2.075 18.745 2.205 ;
 RECT 10.035 1.845 10.165 1.975 ;
 RECT 9.33 1.655 9.46 1.785 ;
 RECT 22.105 0.26 22.235 0.39 ;
 RECT 27.045 1.03 27.175 1.16 ;
 RECT 16.275 0.495 16.405 0.625 ;
 RECT 17.465 1.43 17.595 1.56 ;
 RECT 15.55 0.625 15.68 0.755 ;
 RECT 15.47 1.445 15.6 1.575 ;
 RECT 24.195 1.075 24.325 1.205 ;
 RECT 10.6 0.935 10.73 1.065 ;
 RECT 25.12 0.975 25.25 1.105 ;
 RECT 17.13 0.665 17.26 0.795 ;
 RECT 24.64 1.035 24.77 1.165 ;
 RECT 27.08 2.31 27.21 2.44 ;
 RECT 13.845 2.34 13.975 2.47 ;
 RECT 22.885 0.635 23.015 0.765 ;
 RECT 12.275 1.28 12.405 1.41 ;
 RECT 25.905 0.26 26.035 0.39 ;
 RECT 11.835 1.515 11.965 1.645 ;
 RECT 23.145 1.075 23.275 1.205 ;
 RECT 14.87 0.925 15 1.055 ;
 RECT 7.27 2.11 7.4 2.24 ;
 RECT 12.84 0.595 12.97 0.725 ;
 RECT 0.315 2.345 0.445 2.475 ;
 RECT 0.315 1.825 0.445 1.955 ;
 RECT 20.625 1.705 20.755 1.835 ;
 RECT 16.83 1.835 16.96 1.965 ;
 RECT 5.38 2.345 5.51 2.475 ;
 RECT 9.98 1.23 10.11 1.36 ;
 RECT 0.315 0.33 0.445 0.46 ;
 RECT 4.64 0.74 4.77 0.87 ;
 RECT 9.17 2.265 9.3 2.395 ;
 RECT 5.955 0.79 6.085 0.92 ;
 RECT 27.975 1.475 28.105 1.605 ;
 RECT 19.865 0.92 19.995 1.05 ;
 RECT 8.69 2.135 8.82 2.265 ;
 RECT 26.415 0.12 26.545 0.25 ;
 RECT 5.225 0.145 5.355 0.275 ;
 RECT 21.63 1.705 21.76 1.835 ;
 RECT 21.03 2.64 21.16 2.77 ;
 RECT 17.805 1.035 17.935 1.165 ;
 RECT 11.03 0.905 11.16 1.035 ;
 RECT 14.78 0.595 14.91 0.725 ;
 RECT 25.405 1.445 25.535 1.575 ;
 RECT 4.24 0.325 4.37 0.455 ;
 RECT 10.2 2.3 10.33 2.43 ;
 RECT 9.17 0.315 9.3 0.445 ;
 RECT 6.305 2.105 6.435 2.235 ;
 RECT 6.82 0.88 6.95 1.01 ;
 RECT 14.275 1.9 14.405 2.03 ;
 RECT 19.745 1.705 19.875 1.835 ;
 RECT 18.39 0.91 18.52 1.04 ;
 RECT 16.7 0.765 16.83 0.895 ;
 RECT 13.75 0.875 13.88 1.005 ;
 RECT 6.8 2.07 6.93 2.2 ;
 RECT 2.59 1.6 2.72 1.73 ;
 RECT 19.27 1.705 19.4 1.835 ;
 RECT 1.285 2.275 1.415 2.405 ;
 RECT 7.75 1.825 7.88 1.955 ;
 RECT 3.665 1.75 3.795 1.88 ;
 RECT 21.115 0.5 21.245 0.63 ;
 RECT 0.815 0.735 0.945 0.865 ;
 RECT 26.25 1.49 26.38 1.62 ;
 RECT 24.8 0.435 24.93 0.565 ;
 RECT 11.95 0.89 12.08 1.02 ;
 RECT 20.625 0.975 20.755 1.105 ;
 RECT 4.64 2.05 4.77 2.18 ;
 RECT 7.425 0.53 7.555 0.66 ;
 RECT 4.17 0.74 4.3 0.87 ;
 RECT 12.65 2.225 12.78 2.355 ;
 RECT 4.17 2.115 4.3 2.245 ;
 RECT 24.02 1.475 24.15 1.605 ;
 RECT 25.235 0.12 25.365 0.25 ;
 RECT 17.77 1.835 17.9 1.965 ;
 RECT 27.195 1.465 27.325 1.595 ;
 RECT 15.675 2.38 15.805 2.51 ;
 RECT 5.89 1.825 6.02 1.955 ;
 RECT 21.63 0.975 21.76 1.105 ;
 RECT 9.71 2.235 9.84 2.365 ;
 RECT 1.29 1.51 1.42 1.64 ;
 RECT 23.55 1.425 23.68 1.555 ;
 RECT 25.88 1.405 26.01 1.535 ;
 RECT 18.8 1.705 18.93 1.835 ;
 RECT 11.505 0.905 11.635 1.035 ;
 RECT 11.025 2.015 11.155 2.145 ;
 RECT 3.665 0.735 3.795 0.865 ;
 RECT 24.02 0.135 24.15 0.265 ;
 RECT 7.1 1.525 7.23 1.655 ;
 RECT 1.285 0.735 1.415 0.865 ;
 RECT 6.07 1.49 6.2 1.62 ;
 RECT 2.23 0.735 2.36 0.865 ;
 RECT 3.195 2.31 3.325 2.44 ;
 RECT 14.78 1.87 14.91 2 ;
 RECT 0.315 0.59 0.445 0.72 ;
 RECT 2.425 2.075 2.555 2.205 ;
 RECT 13.015 1.28 13.145 1.41 ;
 RECT 6.705 0.525 6.835 0.655 ;
 RECT 11.95 1.995 12.08 2.125 ;
 RECT 1.285 2.015 1.415 2.145 ;
 RECT 4.76 1.55 4.89 1.68 ;
 RECT 8.22 2.11 8.35 2.24 ;
 RECT 2.41 1.19 2.54 1.32 ;
 RECT 3.195 2.05 3.325 2.18 ;
 RECT 11.505 2.07 11.635 2.2 ;
 RECT 5.295 1.495 5.425 1.625 ;
 RECT 5.245 0.745 5.375 0.875 ;
 RECT 0.315 2.085 0.445 2.215 ;
 RECT 23.3 0.505 23.43 0.635 ;
 RECT 1.89 1.155 2.02 1.285 ;
 RECT 3.665 2.01 3.795 2.14 ;
 RECT 24.8 1.485 24.93 1.615 ;
 RECT 8.035 0.32 8.165 0.45 ;
 LAYER M1 ;
 RECT 27.19 1.385 27.645 1.525 ;
 RECT 25.115 1.145 25.255 1.345 ;
 RECT 24.795 1.485 24.935 1.76 ;
 RECT 25.115 0.73 25.255 0.935 ;
 RECT 24.795 0.355 24.935 0.59 ;
 RECT 24.795 1.345 25.255 1.485 ;
 RECT 25.07 0.935 25.3 1.145 ;
 RECT 24.795 0.59 25.255 0.73 ;
 RECT 23.095 1.225 23.325 1.245 ;
 RECT 23.095 1.195 23.685 1.225 ;
 RECT 23.235 1.015 23.545 1.035 ;
 RECT 23.095 1.035 23.545 1.055 ;
 RECT 23.37 0.64 23.51 1.015 ;
 RECT 23.545 1.225 23.685 1.75 ;
 RECT 23.25 0.5 23.51 0.64 ;
 RECT 24.145 1.035 24.375 1.055 ;
 RECT 24.145 1.195 24.375 1.245 ;
 RECT 23.095 1.055 24.375 1.195 ;
 RECT 22.055 0.36 22.285 0.43 ;
 RECT 23.65 0.36 23.79 0.565 ;
 RECT 22.055 0.22 23.79 0.36 ;
 RECT 24.39 0.705 24.53 0.75 ;
 RECT 24.515 0.995 24.82 1.205 ;
 RECT 24.515 0.89 24.655 0.995 ;
 RECT 24.39 0.75 24.655 0.89 ;
 RECT 23.65 0.565 24.53 0.705 ;
 RECT 17.08 0.57 17.31 0.95 ;
 RECT 17.925 0.42 18.155 0.6 ;
 RECT 19.265 1.385 19.405 1.625 ;
 RECT 19.825 1.105 19.965 1.245 ;
 RECT 19.93 0.42 20.07 0.915 ;
 RECT 19.265 1.245 20.335 1.385 ;
 RECT 20.105 1.385 20.335 1.455 ;
 RECT 19.795 0.92 20.15 1.055 ;
 RECT 19.825 1.055 20.15 1.105 ;
 RECT 19.795 0.915 20.095 0.92 ;
 RECT 17.925 0.28 20.07 0.42 ;
 RECT 19.235 1.625 19.49 1.92 ;
 RECT 17.8 1.545 17.94 1.83 ;
 RECT 17.8 1.17 17.94 1.405 ;
 RECT 16.755 1.83 18.005 1.97 ;
 RECT 17.73 1.03 18.01 1.17 ;
 RECT 18.82 0.765 18.96 1.405 ;
 RECT 19.545 0.56 19.775 0.625 ;
 RECT 19.545 0.765 19.775 0.77 ;
 RECT 18.82 0.625 19.775 0.765 ;
 RECT 17.8 1.405 18.96 1.545 ;
 RECT 14.775 0.525 14.915 0.885 ;
 RECT 14.775 1.095 14.915 2.065 ;
 RECT 14.775 0.885 15.05 1.095 ;
 RECT 11.5 1.04 11.64 2.34 ;
 RECT 11.5 0.895 11.64 0.9 ;
 RECT 11.43 0.9 11.705 1.04 ;
 RECT 12.295 2.055 12.435 2.34 ;
 RECT 11.5 2.34 12.435 2.48 ;
 RECT 13.43 1.66 13.57 1.915 ;
 RECT 12.295 1.915 13.57 2.055 ;
 RECT 13.745 0.765 13.885 1.52 ;
 RECT 13.745 1.66 13.885 2.145 ;
 RECT 14.27 0.525 14.41 1.52 ;
 RECT 14.27 1.66 14.41 2.11 ;
 RECT 13.43 1.52 14.41 1.66 ;
 RECT 15.5 0.585 16.455 0.63 ;
 RECT 16.225 0.63 16.455 0.665 ;
 RECT 16.225 0.455 16.455 0.49 ;
 RECT 15.525 0.49 16.455 0.585 ;
 RECT 15.5 0.63 15.73 0.795 ;
 RECT 5.95 1.67 6.09 1.82 ;
 RECT 5.95 1.96 6.09 2.51 ;
 RECT 5.95 0.5 6.09 1.44 ;
 RECT 5.95 1.44 6.205 1.67 ;
 RECT 5.82 1.82 6.09 1.96 ;
 RECT 8.31 2.445 8.54 2.51 ;
 RECT 8.31 2.65 8.54 2.655 ;
 RECT 5.95 2.51 8.54 2.65 ;
 RECT 3.945 1.335 4.085 2.11 ;
 RECT 3.945 2.25 4.085 2.255 ;
 RECT 3.945 0.875 4.085 1.195 ;
 RECT 3.945 2.11 4.37 2.25 ;
 RECT 3.945 0.735 4.37 0.875 ;
 RECT 3.945 1.195 5.055 1.335 ;
 RECT 4.915 0.6 5.055 1.195 ;
 RECT 6.345 0.36 6.485 2.035 ;
 RECT 5.66 0.22 6.485 0.36 ;
 RECT 5.66 0.36 5.8 0.46 ;
 RECT 6.3 2.17 6.44 2.305 ;
 RECT 6.3 2.035 6.485 2.17 ;
 RECT 4.915 0.46 5.8 0.6 ;
 RECT 7.095 0.66 7.235 0.895 ;
 RECT 6.635 0.52 7.235 0.66 ;
 RECT 7.095 0.895 10.78 1.035 ;
 RECT 10.55 1.035 10.78 1.105 ;
 RECT 5.195 0.88 5.335 1.475 ;
 RECT 5.155 1.63 5.295 1.99 ;
 RECT 5.155 1.475 5.5 1.63 ;
 RECT 5.045 1.99 5.295 2.13 ;
 RECT 5.195 0.74 5.515 0.88 ;
 RECT 3.66 0.46 3.8 2.21 ;
 RECT 4.13 0.22 4.495 0.32 ;
 RECT 4.13 0.46 4.495 0.525 ;
 RECT 3.66 0.32 4.495 0.46 ;
 RECT 2.88 0.87 3.02 1.15 ;
 RECT 2.88 1.29 3.02 2.07 ;
 RECT 2.37 2.07 3.02 2.21 ;
 RECT 2.175 0.73 3.02 0.87 ;
 RECT 3.28 1.115 3.51 1.15 ;
 RECT 3.28 1.29 3.51 1.325 ;
 RECT 2.88 1.15 3.51 1.29 ;
 RECT 0.81 0.68 0.95 1.155 ;
 RECT 0.81 1.295 0.95 2.23 ;
 RECT 1.595 0.36 1.735 1.155 ;
 RECT 0.81 1.155 1.735 1.295 ;
 RECT 2.815 0.36 3.045 0.43 ;
 RECT 1.595 0.22 3.045 0.36 ;
 RECT 16.19 1.895 16.33 2.39 ;
 RECT 20.335 2.205 20.475 2.39 ;
 RECT 16.19 2.39 20.475 2.53 ;
 RECT 15.065 1.755 16.33 1.895 ;
 RECT 15.065 1.895 15.205 2.34 ;
 RECT 13.795 2.3 14.025 2.34 ;
 RECT 13.795 2.48 14.025 2.51 ;
 RECT 13.795 2.34 15.205 2.48 ;
 RECT 20.335 2.065 22.83 2.205 ;
 RECT 22.69 2.205 22.83 2.52 ;
 RECT 27.03 2.48 27.17 2.52 ;
 RECT 22.69 2.52 27.17 2.66 ;
 RECT 27.03 2.27 27.26 2.48 ;
 RECT 18.74 1.7 19.075 1.84 ;
 RECT 18.935 1.84 19.075 2.075 ;
 RECT 19.63 1.84 19.77 2.075 ;
 RECT 19.63 1.7 19.925 1.84 ;
 RECT 18.935 2.075 19.77 2.215 ;
 RECT 16.47 1.56 16.61 2.11 ;
 RECT 15.42 1.405 15.65 1.42 ;
 RECT 15.42 1.56 15.65 1.615 ;
 RECT 15.42 1.42 16.61 1.56 ;
 RECT 16.47 2.11 18.795 2.245 ;
 RECT 16.47 2.245 18.79 2.25 ;
 RECT 18.565 2.035 18.795 2.11 ;
 RECT 11.945 1.025 12.085 1.475 ;
 RECT 11.785 1.475 12.085 1.635 ;
 RECT 11.945 1.775 12.085 2.18 ;
 RECT 11.875 0.885 12.15 1.025 ;
 RECT 11.945 1.685 13.15 1.775 ;
 RECT 13.01 1.415 13.15 1.635 ;
 RECT 11.785 1.635 13.15 1.685 ;
 RECT 12.955 1.275 13.215 1.415 ;
 RECT 7.2 2.105 8.42 2.245 ;
 RECT 9.705 1.365 9.845 2.43 ;
 RECT 7.76 1.365 7.9 1.5 ;
 RECT 6.93 1.64 7.435 1.675 ;
 RECT 6.93 1.5 7.9 1.64 ;
 RECT 11.02 1.04 11.16 1.25 ;
 RECT 11.02 1.39 11.16 2.215 ;
 RECT 11.02 0.885 11.16 0.9 ;
 RECT 7.76 1.25 11.16 1.365 ;
 RECT 7.76 1.225 10.41 1.25 ;
 RECT 10.27 1.365 11.16 1.39 ;
 RECT 10.955 0.9 11.23 1.04 ;
 RECT 6.725 1.96 7.005 2.215 ;
 RECT 8.08 1.79 8.22 1.82 ;
 RECT 6.64 1.22 6.955 1.36 ;
 RECT 6.815 0.805 6.955 1.22 ;
 RECT 6.64 1.82 8.22 1.96 ;
 RECT 6.64 1.36 6.78 1.82 ;
 RECT 9.28 1.615 9.51 1.65 ;
 RECT 9.28 1.79 9.51 1.825 ;
 RECT 8.08 1.65 9.515 1.79 ;
 RECT 25.735 0.73 25.875 1.04 ;
 RECT 25.875 1.18 26.015 1.605 ;
 RECT 25.67 0.59 25.945 0.73 ;
 RECT 26.995 0.99 27.225 1.04 ;
 RECT 25.735 1.04 27.225 1.18 ;
 RECT 26.995 1.18 27.225 1.2 ;
 RECT 25.855 0.29 26.225 0.43 ;
 RECT 26.085 0.43 26.225 0.71 ;
 RECT 25.855 0.22 26.085 0.29 ;
 RECT 27.505 0.85 27.645 1.385 ;
 RECT 27.19 1.525 27.33 1.73 ;
 RECT 26.085 0.71 27.645 0.85 ;
 RECT 27.19 0.51 27.33 0.71 ;
 END
END RSDFFNSRASRNX1

MACRO RSDFFNSRASRNX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 29.44 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.615 0.59 22.985 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 27.845 1.435 28.185 1.8 ;
 RECT 26.165 1.99 28.03 2.13 ;
 RECT 23.935 2.22 26.305 2.36 ;
 RECT 26.165 1.435 26.305 1.99 ;
 RECT 27.89 1.8 28.03 1.99 ;
 RECT 23.935 1.39 24.075 2.22 ;
 RECT 25.32 1.37 25.46 2.22 ;
 RECT 26.165 2.13 26.305 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 29.44 0.08 ;
 RECT 5.155 0.08 5.435 0.295 ;
 RECT 26.285 0.08 26.525 0.26 ;
 RECT 9.085 0.31 9.375 0.45 ;
 RECT 12.77 0.59 13.045 0.73 ;
 RECT 16.695 0.275 17.72 0.415 ;
 RECT 21.055 0.335 21.32 0.495 ;
 RECT 17.58 0.75 18.525 0.89 ;
 RECT 1.28 0.08 1.42 0.93 ;
 RECT 0.31 0.08 0.45 0.775 ;
 RECT 3.19 0.08 3.33 0.74 ;
 RECT 4.635 0.08 4.775 0.97 ;
 RECT 7.98 0.08 8.215 0.46 ;
 RECT 23.935 0.08 24.075 0.36 ;
 RECT 25.15 0.08 25.29 0.35 ;
 RECT 9.165 0.08 9.305 0.31 ;
 RECT 12.835 0.08 12.975 0.59 ;
 RECT 16.695 0.415 16.835 0.945 ;
 RECT 16.695 0.08 16.835 0.275 ;
 RECT 21.11 0.08 21.25 0.335 ;
 RECT 18.385 0.89 18.525 1.11 ;
 RECT 17.58 0.415 17.72 0.75 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.62 1.205 20.9 1.445 ;
 RECT 20.62 0.595 20.76 1.205 ;
 RECT 21.625 1.84 21.765 1.885 ;
 RECT 21.625 0.62 21.765 1.7 ;
 RECT 20.62 1.84 20.76 1.885 ;
 RECT 20.62 1.7 21.765 1.84 ;
 RECT 20.62 1.445 20.76 1.7 ;
 END
 ANTENNADIFFAREA 1.089 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 12.58 2.215 12.855 2.355 ;
 RECT 21.04 2.345 21.305 2.545 ;
 RECT 0 2.8 29.44 2.96 ;
 RECT 1.28 1.965 1.42 2.8 ;
 RECT 0.31 1.74 0.45 2.8 ;
 RECT 5.31 2.34 5.56 2.8 ;
 RECT 3.19 1.99 3.33 2.8 ;
 RECT 4.635 1.98 4.775 2.8 ;
 RECT 8.685 2.07 8.825 2.8 ;
 RECT 10.195 2 10.335 2.8 ;
 RECT 9.165 1.98 9.305 2.8 ;
 RECT 15.605 2.335 15.875 2.8 ;
 RECT 12.645 2.355 12.785 2.8 ;
 RECT 12.645 2.195 12.785 2.215 ;
 RECT 21.115 2.545 21.255 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.685 1.475 5.015 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.225 1.155 12.6 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.055 0.44 12.435 0.58 ;
 RECT 7.375 0.485 7.785 0.605 ;
 RECT 7.375 0.605 10.195 0.745 ;
 RECT 10.055 0.58 10.195 0.605 ;
 RECT 13.21 1.015 13.35 1.02 ;
 RECT 12.295 0.875 13.35 1.015 ;
 RECT 13.21 0.245 15.355 0.255 ;
 RECT 13.21 0.255 15.36 0.385 ;
 RECT 15.22 1.09 17.21 1.23 ;
 RECT 17.415 1.56 17.645 1.6 ;
 RECT 17.07 1.42 17.645 1.56 ;
 RECT 17.415 1.39 17.645 1.42 ;
 RECT 12.295 0.58 12.435 0.875 ;
 RECT 13.21 0.385 13.35 0.875 ;
 RECT 15.22 0.385 15.36 1.09 ;
 RECT 17.07 1.23 17.21 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.985 1.51 10.425 1.855 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.1 1.435 1.625 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.79 1.59 2.735 1.75 ;
 RECT 1.885 1.09 2.025 1.44 ;
 RECT 1.79 1.44 2.035 1.59 ;
 RECT 2.585 1.75 2.725 1.805 ;
 RECT 2.585 1.53 2.725 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.25 1.115 2.67 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 OBS
 LAYER PO ;
 RECT 14.525 1.29 15.615 1.39 ;
 RECT 5.67 2.675 6.655 2.775 ;
 RECT 15.42 1.405 15.65 1.615 ;
 RECT 24.195 1.245 24.295 2.02 ;
 RECT 24.065 1.035 24.295 1.245 ;
 RECT 15.915 0.105 18.74 0.205 ;
 RECT 15.915 0.205 16.015 1.91 ;
 RECT 18.64 0.205 18.74 1.265 ;
 RECT 15.095 1.71 15.195 1.91 ;
 RECT 14.01 1.61 15.195 1.71 ;
 RECT 14.01 0.475 14.11 1.61 ;
 RECT 14.56 1.71 14.66 2.425 ;
 RECT 10.68 0.375 14.11 0.475 ;
 RECT 10.68 0.475 10.78 0.815 ;
 RECT 15.095 1.91 16.015 2.01 ;
 RECT 10.55 0.815 10.78 1.025 ;
 RECT 17.925 0.39 18.155 0.45 ;
 RECT 16.225 0.45 18.155 0.55 ;
 RECT 17.925 0.55 18.155 0.6 ;
 RECT 16.225 0.55 16.455 0.665 ;
 RECT 17.08 0.55 17.31 0.835 ;
 RECT 17.08 0.835 17.18 2.39 ;
 RECT 24.5 0.215 24.6 0.995 ;
 RECT 24.5 0.995 24.74 1.205 ;
 RECT 24.5 1.205 24.6 2 ;
 RECT 26.895 0.375 26.995 0.99 ;
 RECT 26.895 0.99 27.145 1.2 ;
 RECT 26.895 1.2 26.995 2.27 ;
 RECT 26.895 2.27 27.18 2.48 ;
 RECT 13.49 0.655 13.59 2.305 ;
 RECT 13.795 2.3 14.025 2.305 ;
 RECT 13.795 2.405 14.025 2.51 ;
 RECT 13.49 2.305 14.025 2.405 ;
 RECT 23.72 0.855 23.82 2.2 ;
 RECT 26.585 1.125 26.685 2.2 ;
 RECT 22.755 0.755 24.29 0.84 ;
 RECT 22.755 0.84 24.285 0.855 ;
 RECT 24.19 0.215 24.29 0.755 ;
 RECT 23.72 0.21 23.82 0.755 ;
 RECT 22.755 0.595 22.985 0.755 ;
 RECT 23.72 2.2 26.685 2.3 ;
 RECT 12.2 1.28 12.455 1.45 ;
 RECT 12.2 1.45 12.3 1.655 ;
 RECT 12.2 0.655 12.3 1.18 ;
 RECT 12.2 1.655 13.16 1.755 ;
 RECT 13.06 1.755 13.16 2.355 ;
 RECT 11.285 0.66 11.385 1.18 ;
 RECT 12.2 1.755 12.3 2.51 ;
 RECT 11.285 1.24 12.455 1.28 ;
 RECT 11.285 1.18 12.3 1.24 ;
 RECT 25.41 0.38 25.51 0.96 ;
 RECT 25.41 1.06 25.51 1.14 ;
 RECT 24.99 0.935 25.22 0.96 ;
 RECT 24.99 0.96 25.51 1.06 ;
 RECT 24.99 1.06 25.22 1.145 ;
 RECT 25.41 1.14 25.68 1.24 ;
 RECT 25.58 1.24 25.68 1.84 ;
 RECT 25.775 0.22 26.005 0.28 ;
 RECT 25.775 0.38 26.005 0.43 ;
 RECT 25.41 0.28 26.005 0.38 ;
 RECT 11.275 1.575 11.375 2.485 ;
 RECT 11.785 1.575 12.015 1.685 ;
 RECT 11.275 1.475 12.015 1.575 ;
 RECT 27.595 0.195 27.695 2.665 ;
 RECT 26.585 0.095 27.695 0.195 ;
 RECT 22.96 1.245 23.06 2.665 ;
 RECT 22.96 1.2 23.245 1.245 ;
 RECT 26.585 0.195 26.685 0.945 ;
 RECT 23.015 1.035 23.245 1.1 ;
 RECT 22.96 2.665 27.695 2.765 ;
 RECT 22.96 1.1 23.29 1.2 ;
 RECT 15.5 0.795 15.665 0.925 ;
 RECT 14.82 0.885 15.05 0.925 ;
 RECT 14.82 1.025 15.05 1.095 ;
 RECT 14.82 0.925 15.665 1.025 ;
 RECT 15.5 0.585 15.73 0.795 ;
 RECT 4.42 0.52 4.52 2.465 ;
 RECT 4.18 0.27 4.52 0.52 ;
 RECT 7.05 1.33 7.19 1.475 ;
 RECT 7.05 1.71 7.15 2.475 ;
 RECT 7.09 0.65 7.19 1.33 ;
 RECT 7.05 1.475 7.28 1.71 ;
 RECT 1.87 0.515 1.97 1.105 ;
 RECT 1.83 1.105 2.075 1.345 ;
 RECT 6.6 0.705 6.7 1.165 ;
 RECT 6.16 1.27 6.26 1.445 ;
 RECT 6.6 0.47 6.885 0.705 ;
 RECT 6.16 1.17 6.7 1.265 ;
 RECT 6.16 1.265 6.535 1.27 ;
 RECT 6.39 1.165 6.7 1.17 ;
 RECT 6.015 1.445 6.26 1.69 ;
 RECT 13.095 0.655 13.195 1.24 ;
 RECT 12.965 1.24 13.195 1.475 ;
 RECT 2.255 1.37 2.355 1.605 ;
 RECT 2.485 0.515 2.585 1.14 ;
 RECT 2.205 1.705 2.305 2.695 ;
 RECT 2.205 1.605 2.355 1.705 ;
 RECT 2.255 1.14 2.585 1.37 ;
 RECT 4.895 0.49 4.995 1.495 ;
 RECT 4.7 1.495 4.995 1.745 ;
 RECT 4.895 1.745 4.995 2.37 ;
 RECT 2.675 1.78 2.775 2.695 ;
 RECT 2.535 1.55 2.775 1.78 ;
 RECT 1.065 1.435 1.635 1.71 ;
 RECT 1.535 0.515 1.635 1.435 ;
 RECT 1.535 1.71 1.635 2.695 ;
 RECT 1.065 0.515 1.165 1.435 ;
 RECT 1.065 1.71 1.165 2.645 ;
 RECT 7.49 0.715 7.59 1.61 ;
 RECT 7.525 1.71 7.625 2.48 ;
 RECT 7.49 1.61 7.625 1.71 ;
 RECT 7.37 0.485 7.61 0.715 ;
 RECT 2.975 0.135 3.075 0.22 ;
 RECT 2.815 0.22 3.075 0.43 ;
 RECT 2.975 0.43 3.075 2.695 ;
 RECT 3.445 0.295 3.545 1.115 ;
 RECT 3.28 1.115 3.545 1.325 ;
 RECT 3.445 1.325 3.545 2.74 ;
 RECT 20.885 0.375 20.985 1.36 ;
 RECT 20.105 1.4 21.475 1.46 ;
 RECT 20.885 1.46 21.475 1.5 ;
 RECT 20.105 1.36 20.985 1.4 ;
 RECT 20.885 1.5 20.985 2.765 ;
 RECT 21.375 0.375 21.475 1.4 ;
 RECT 21.375 1.5 21.475 2.765 ;
 RECT 20.105 1.245 20.335 1.36 ;
 RECT 8.31 2.445 8.57 2.655 ;
 RECT 8.47 1.79 8.57 2.445 ;
 RECT 18.58 1.445 18.68 2.035 ;
 RECT 18.565 2.035 18.795 2.245 ;
 RECT 19.05 0.55 19.15 2.69 ;
 RECT 9.98 1.83 10.08 2.69 ;
 RECT 9.98 1.58 10.08 1.62 ;
 RECT 9.72 1.01 9.82 1.48 ;
 RECT 9.98 1.62 10.215 1.83 ;
 RECT 9.98 2.69 19.15 2.79 ;
 RECT 9.72 1.48 10.08 1.58 ;
 RECT 9.42 0.98 9.52 1.615 ;
 RECT 9.28 1.615 9.52 1.825 ;
 RECT 9.42 1.825 9.52 2.51 ;
 RECT 19.52 0.56 19.775 0.615 ;
 RECT 19.52 0.55 19.62 0.56 ;
 RECT 19.52 0.615 20.34 0.715 ;
 RECT 19.52 0.715 19.775 0.77 ;
 RECT 19.52 0.77 19.62 2.155 ;
 RECT 20.24 0.19 20.34 0.615 ;
 RECT 21.975 0.19 22.205 0.43 ;
 RECT 20.24 0.09 22.205 0.19 ;
 RECT 17.55 0.73 17.65 1.39 ;
 RECT 17.415 1.39 17.65 1.6 ;
 RECT 17.55 1.6 17.65 2.39 ;
 RECT 5.735 0.285 5.835 1.52 ;
 RECT 5.235 1.52 5.835 1.62 ;
 RECT 5.735 0.185 14.625 0.195 ;
 RECT 7.79 0.095 14.625 0.185 ;
 RECT 5.735 0.195 7.89 0.285 ;
 RECT 14.525 0.195 14.625 1.29 ;
 RECT 15.42 1.39 15.615 1.405 ;
 RECT 6.555 1.565 6.655 2.675 ;
 RECT 5.67 1.62 5.77 2.675 ;
 RECT 5.235 1.44 5.48 1.52 ;
 RECT 5.235 1.62 5.48 1.69 ;
 RECT 7.79 0.285 7.89 1.24 ;
 LAYER CO ;
 RECT 19.27 1.705 19.4 1.835 ;
 RECT 3.195 0.545 3.325 0.675 ;
 RECT 21.115 0.36 21.245 0.49 ;
 RECT 3.665 0.735 3.795 0.865 ;
 RECT 24.72 0.435 24.85 0.565 ;
 RECT 20.625 1.705 20.755 1.835 ;
 RECT 5.38 2.345 5.51 2.475 ;
 RECT 21.63 1.705 21.76 1.835 ;
 RECT 6.82 0.88 6.95 1.01 ;
 RECT 21.12 2.395 21.25 2.525 ;
 RECT 1.89 1.155 2.02 1.285 ;
 RECT 6.35 0.88 6.48 1.01 ;
 RECT 2.865 0.26 2.995 0.39 ;
 RECT 3.33 1.155 3.46 1.285 ;
 RECT 20.155 1.285 20.285 1.415 ;
 RECT 17.975 0.43 18.105 0.56 ;
 RECT 19.595 0.6 19.725 0.73 ;
 RECT 8.36 2.485 8.49 2.615 ;
 RECT 18.615 2.075 18.745 2.205 ;
 RECT 10.035 1.66 10.165 1.79 ;
 RECT 9.33 1.655 9.46 1.785 ;
 RECT 22.025 0.26 22.155 0.39 ;
 RECT 26.965 1.03 27.095 1.16 ;
 RECT 16.275 0.495 16.405 0.625 ;
 RECT 17.465 1.43 17.595 1.56 ;
 RECT 15.55 0.625 15.68 0.755 ;
 RECT 15.47 1.445 15.6 1.575 ;
 RECT 24.115 1.075 24.245 1.205 ;
 RECT 10.6 0.855 10.73 0.985 ;
 RECT 25.04 0.975 25.17 1.105 ;
 RECT 17.13 0.665 17.26 0.795 ;
 RECT 24.56 1.035 24.69 1.165 ;
 RECT 27 2.31 27.13 2.44 ;
 RECT 13.845 2.34 13.975 2.47 ;
 RECT 22.805 0.635 22.935 0.765 ;
 RECT 12.275 1.28 12.405 1.41 ;
 RECT 25.825 0.26 25.955 0.39 ;
 RECT 11.835 1.515 11.965 1.645 ;
 RECT 23.065 1.075 23.195 1.205 ;
 RECT 14.87 0.925 15 1.055 ;
 RECT 25.325 1.445 25.455 1.575 ;
 RECT 18.39 0.91 18.52 1.04 ;
 RECT 3.195 2.31 3.325 2.44 ;
 RECT 6.305 2.105 6.435 2.235 ;
 RECT 14.78 0.595 14.91 0.725 ;
 RECT 19.745 1.705 19.875 1.835 ;
 RECT 6.07 1.49 6.2 1.62 ;
 RECT 1.285 0.735 1.415 0.865 ;
 RECT 14.275 1.9 14.405 2.03 ;
 RECT 0.315 0.59 0.445 0.72 ;
 RECT 6.705 0.525 6.835 0.655 ;
 RECT 8.22 2.11 8.35 2.24 ;
 RECT 14.78 1.87 14.91 2 ;
 RECT 20.625 0.68 20.755 0.81 ;
 RECT 21.63 0.715 21.76 0.845 ;
 RECT 9.17 2.075 9.3 2.205 ;
 RECT 8.035 0.32 8.165 0.45 ;
 RECT 23.94 0.135 24.07 0.265 ;
 RECT 5.225 0.145 5.355 0.275 ;
 RECT 9.17 0.315 9.3 0.445 ;
 RECT 14.275 0.595 14.405 0.725 ;
 RECT 8.69 2.135 8.82 2.265 ;
 RECT 11.03 0.905 11.16 1.035 ;
 RECT 11.025 2.015 11.155 2.145 ;
 RECT 7.1 1.525 7.23 1.655 ;
 RECT 4.24 0.325 4.37 0.455 ;
 RECT 17.805 1.035 17.935 1.165 ;
 RECT 5.245 0.745 5.375 0.875 ;
 RECT 4.64 2.05 4.77 2.18 ;
 RECT 6.8 2.07 6.93 2.2 ;
 RECT 0.815 0.735 0.945 0.865 ;
 RECT 20.625 0.94 20.755 1.07 ;
 RECT 0.315 2.085 0.445 2.215 ;
 RECT 4.17 2.115 4.3 2.245 ;
 RECT 7.425 0.53 7.555 0.66 ;
 RECT 21.63 0.975 21.76 1.105 ;
 RECT 17.77 1.835 17.9 1.965 ;
 RECT 15.675 2.38 15.805 2.51 ;
 RECT 2.59 1.6 2.72 1.73 ;
 RECT 26.17 1.49 26.3 1.62 ;
 RECT 25.8 1.405 25.93 1.535 ;
 RECT 3.665 1.75 3.795 1.88 ;
 RECT 4.76 1.55 4.89 1.68 ;
 RECT 2.23 0.735 2.36 0.865 ;
 RECT 2.425 2.075 2.555 2.205 ;
 RECT 11.95 1.995 12.08 2.125 ;
 RECT 11.505 2.07 11.635 2.2 ;
 RECT 13.015 1.28 13.145 1.41 ;
 RECT 3.195 2.05 3.325 2.18 ;
 RECT 1.285 2.015 1.415 2.145 ;
 RECT 5.295 1.495 5.425 1.625 ;
 RECT 2.41 1.19 2.54 1.32 ;
 RECT 5.115 1.995 5.245 2.125 ;
 RECT 16.7 0.765 16.83 0.895 ;
 RECT 13.75 0.875 13.88 1.005 ;
 RECT 0.315 2.345 0.445 2.475 ;
 RECT 1.285 2.275 1.415 2.405 ;
 RECT 4.64 0.74 4.77 0.87 ;
 RECT 9.71 2.045 9.84 2.175 ;
 RECT 26.335 0.12 26.465 0.25 ;
 RECT 7.75 1.825 7.88 1.955 ;
 RECT 7.27 2.11 7.4 2.24 ;
 RECT 27.895 1.475 28.025 1.605 ;
 RECT 13.75 1.945 13.88 2.075 ;
 RECT 10.2 2.11 10.33 2.24 ;
 RECT 1.29 1.51 1.42 1.64 ;
 RECT 4.17 0.74 4.3 0.87 ;
 RECT 12.84 0.595 12.97 0.725 ;
 RECT 23.22 0.505 23.35 0.635 ;
 RECT 23.94 1.475 24.07 1.605 ;
 RECT 0.315 0.33 0.445 0.46 ;
 RECT 24.72 1.485 24.85 1.615 ;
 RECT 11.505 0.905 11.635 1.035 ;
 RECT 11.95 0.885 12.08 1.015 ;
 RECT 27.115 1.465 27.245 1.595 ;
 RECT 27.115 0.595 27.245 0.725 ;
 RECT 16.83 1.835 16.96 1.965 ;
 RECT 9.98 1.23 10.11 1.36 ;
 RECT 5.89 1.825 6.02 1.955 ;
 RECT 25.155 0.12 25.285 0.25 ;
 RECT 5.955 0.79 6.085 0.92 ;
 RECT 25.66 0.595 25.79 0.725 ;
 RECT 12.65 2.225 12.78 2.355 ;
 RECT 23.47 1.425 23.6 1.555 ;
 RECT 0.315 1.825 0.445 1.955 ;
 RECT 19.865 0.92 19.995 1.05 ;
 RECT 3.665 2.01 3.795 2.14 ;
 RECT 0.815 2.015 0.945 2.145 ;
 RECT 18.8 1.705 18.93 1.835 ;
 LAYER M1 ;
 RECT 25.655 0.73 25.795 1.04 ;
 RECT 25.795 1.18 25.935 1.605 ;
 RECT 25.59 0.59 25.865 0.73 ;
 RECT 26.915 0.99 27.145 1.04 ;
 RECT 25.655 1.04 27.145 1.18 ;
 RECT 26.915 1.18 27.145 1.2 ;
 RECT 25.775 0.29 26.145 0.43 ;
 RECT 26.005 0.43 26.145 0.71 ;
 RECT 25.775 0.22 26.005 0.29 ;
 RECT 27.425 0.85 27.565 1.385 ;
 RECT 27.11 1.525 27.25 1.73 ;
 RECT 26.005 0.71 27.565 0.85 ;
 RECT 27.11 0.51 27.25 0.71 ;
 RECT 27.11 1.385 27.565 1.525 ;
 RECT 25.035 1.145 25.175 1.345 ;
 RECT 24.715 1.485 24.855 1.76 ;
 RECT 25.035 0.73 25.175 0.935 ;
 RECT 24.715 0.355 24.855 0.59 ;
 RECT 24.715 1.345 25.175 1.485 ;
 RECT 24.99 0.935 25.22 1.145 ;
 RECT 24.715 0.59 25.175 0.73 ;
 RECT 23.015 1.225 23.245 1.245 ;
 RECT 23.015 1.195 23.605 1.225 ;
 RECT 23.155 1.015 23.465 1.035 ;
 RECT 23.015 1.035 23.465 1.055 ;
 RECT 23.29 0.64 23.43 1.015 ;
 RECT 23.465 1.225 23.605 1.75 ;
 RECT 23.17 0.5 23.43 0.64 ;
 RECT 24.065 1.035 24.295 1.055 ;
 RECT 24.065 1.195 24.295 1.245 ;
 RECT 23.015 1.055 24.295 1.195 ;
 RECT 21.975 0.36 22.205 0.43 ;
 RECT 23.57 0.36 23.71 0.565 ;
 RECT 21.975 0.22 23.71 0.36 ;
 RECT 24.31 0.705 24.45 0.75 ;
 RECT 24.435 0.995 24.74 1.205 ;
 RECT 24.435 0.89 24.575 0.995 ;
 RECT 24.31 0.75 24.575 0.89 ;
 RECT 23.57 0.565 24.45 0.705 ;
 RECT 17.08 0.57 17.31 0.95 ;
 RECT 17.925 0.42 18.155 0.6 ;
 RECT 19.265 1.385 19.405 1.625 ;
 RECT 19.825 1.055 19.965 1.245 ;
 RECT 19.915 0.42 20.055 0.915 ;
 RECT 19.265 1.245 20.335 1.385 ;
 RECT 20.105 1.385 20.335 1.455 ;
 RECT 17.925 0.28 20.055 0.42 ;
 RECT 19.235 1.625 19.49 1.92 ;
 RECT 19.795 0.915 20.08 1.055 ;
 RECT 17.8 1.545 17.94 1.83 ;
 RECT 17.8 1.17 17.94 1.405 ;
 RECT 16.755 1.83 18.005 1.97 ;
 RECT 17.73 1.03 18.01 1.17 ;
 RECT 18.82 0.765 18.96 1.405 ;
 RECT 19.545 0.56 19.775 0.625 ;
 RECT 19.545 0.765 19.775 0.77 ;
 RECT 18.82 0.625 19.775 0.765 ;
 RECT 17.8 1.405 18.96 1.545 ;
 RECT 11.5 1.04 11.64 2.34 ;
 RECT 11.5 0.895 11.64 0.9 ;
 RECT 11.43 0.9 11.705 1.04 ;
 RECT 12.295 2.055 12.435 2.34 ;
 RECT 11.5 2.34 12.435 2.48 ;
 RECT 13.43 1.66 13.57 1.915 ;
 RECT 12.295 1.915 13.57 2.055 ;
 RECT 13.745 0.765 13.885 1.52 ;
 RECT 13.745 1.66 13.885 2.145 ;
 RECT 14.27 0.525 14.41 1.52 ;
 RECT 14.27 1.66 14.41 2.11 ;
 RECT 13.43 1.52 14.41 1.66 ;
 RECT 14.775 0.525 14.915 0.885 ;
 RECT 14.775 1.095 14.915 2.065 ;
 RECT 14.775 0.885 15.05 1.095 ;
 RECT 15.5 0.585 16.455 0.63 ;
 RECT 16.225 0.63 16.455 0.665 ;
 RECT 16.225 0.455 16.455 0.49 ;
 RECT 15.525 0.49 16.455 0.585 ;
 RECT 15.5 0.63 15.73 0.795 ;
 RECT 5.95 1.67 6.09 1.82 ;
 RECT 5.95 1.96 6.09 2.51 ;
 RECT 5.95 0.5 6.09 1.44 ;
 RECT 5.95 1.44 6.205 1.67 ;
 RECT 5.82 1.82 6.09 1.96 ;
 RECT 8.31 2.445 8.54 2.51 ;
 RECT 8.31 2.65 8.54 2.655 ;
 RECT 5.95 2.51 8.54 2.65 ;
 RECT 7.095 0.66 7.235 0.885 ;
 RECT 7.095 1.025 7.235 1.035 ;
 RECT 6.635 0.52 7.235 0.66 ;
 RECT 10.55 0.815 10.78 0.885 ;
 RECT 7.095 0.885 10.78 1.025 ;
 RECT 3.945 1.335 4.085 2.11 ;
 RECT 3.945 2.25 4.085 2.255 ;
 RECT 3.945 0.875 4.085 1.195 ;
 RECT 3.945 2.11 4.37 2.25 ;
 RECT 3.945 0.735 4.37 0.875 ;
 RECT 3.945 1.195 5.055 1.335 ;
 RECT 4.915 0.6 5.055 1.195 ;
 RECT 6.345 0.36 6.485 2.035 ;
 RECT 5.66 0.22 6.485 0.36 ;
 RECT 5.66 0.36 5.8 0.46 ;
 RECT 6.3 2.17 6.44 2.305 ;
 RECT 6.3 2.035 6.485 2.17 ;
 RECT 4.915 0.46 5.8 0.6 ;
 RECT 3.66 0.46 3.8 2.21 ;
 RECT 4.13 0.22 4.495 0.32 ;
 RECT 4.13 0.46 4.495 0.525 ;
 RECT 3.66 0.32 4.495 0.46 ;
 RECT 0.81 0.68 0.95 1.155 ;
 RECT 0.81 1.295 0.95 2.23 ;
 RECT 1.595 0.36 1.735 1.155 ;
 RECT 0.81 1.155 1.735 1.295 ;
 RECT 2.815 0.36 3.045 0.43 ;
 RECT 1.595 0.22 3.045 0.36 ;
 RECT 16.19 1.895 16.33 2.39 ;
 RECT 20.335 2.205 20.475 2.39 ;
 RECT 16.19 2.39 20.475 2.53 ;
 RECT 15.065 1.755 16.33 1.895 ;
 RECT 15.065 1.895 15.205 2.34 ;
 RECT 13.795 2.3 14.025 2.34 ;
 RECT 13.795 2.48 14.025 2.51 ;
 RECT 13.795 2.34 15.205 2.48 ;
 RECT 20.335 2.065 22.75 2.205 ;
 RECT 22.61 2.205 22.75 2.52 ;
 RECT 26.95 2.48 27.09 2.52 ;
 RECT 22.61 2.52 27.09 2.66 ;
 RECT 26.95 2.27 27.18 2.48 ;
 RECT 18.74 1.7 19.075 1.84 ;
 RECT 18.935 1.84 19.075 2.075 ;
 RECT 19.63 1.7 19.925 1.84 ;
 RECT 19.63 1.84 19.77 2.075 ;
 RECT 18.935 2.075 19.77 2.215 ;
 RECT 16.47 1.56 16.61 2.11 ;
 RECT 15.42 1.405 15.65 1.42 ;
 RECT 15.42 1.56 15.65 1.615 ;
 RECT 15.42 1.42 16.61 1.56 ;
 RECT 16.47 2.11 18.795 2.245 ;
 RECT 16.47 2.245 18.79 2.25 ;
 RECT 18.565 2.035 18.795 2.11 ;
 RECT 11.945 1.02 12.085 1.475 ;
 RECT 11.785 1.475 12.085 1.635 ;
 RECT 11.945 1.775 12.085 2.18 ;
 RECT 11.875 0.88 12.15 1.02 ;
 RECT 11.945 1.685 13.15 1.775 ;
 RECT 13.01 1.415 13.15 1.635 ;
 RECT 11.785 1.635 13.15 1.685 ;
 RECT 12.96 1.275 13.215 1.415 ;
 RECT 7.2 2.105 8.42 2.245 ;
 RECT 9.705 1.365 9.845 2.25 ;
 RECT 7.755 1.365 7.895 1.5 ;
 RECT 6.93 1.5 7.895 1.64 ;
 RECT 6.93 1.64 7.435 1.675 ;
 RECT 11.02 0.885 11.16 0.9 ;
 RECT 11.02 1.04 11.16 1.225 ;
 RECT 11.02 1.365 11.16 2.215 ;
 RECT 10.955 0.9 11.23 1.04 ;
 RECT 7.755 1.225 11.16 1.365 ;
 RECT 5.195 0.88 5.335 1.475 ;
 RECT 5.155 1.63 5.295 1.99 ;
 RECT 5.155 1.475 5.5 1.63 ;
 RECT 5.195 0.74 5.515 0.88 ;
 RECT 5.045 1.99 5.295 2.13 ;
 RECT 6.64 1.82 8.22 1.96 ;
 RECT 8.08 1.79 8.22 1.82 ;
 RECT 6.64 1.22 6.955 1.36 ;
 RECT 6.815 0.805 6.955 1.22 ;
 RECT 6.725 1.96 7.005 2.215 ;
 RECT 6.64 1.36 6.78 1.82 ;
 RECT 9.28 1.615 9.51 1.65 ;
 RECT 9.28 1.79 9.51 1.825 ;
 RECT 8.08 1.65 9.515 1.79 ;
 RECT 2.88 0.87 3.02 1.15 ;
 RECT 2.88 1.29 3.02 2.07 ;
 RECT 2.175 0.73 3.02 0.87 ;
 RECT 2.37 2.07 3.02 2.21 ;
 RECT 3.28 1.115 3.51 1.15 ;
 RECT 3.28 1.29 3.51 1.325 ;
 RECT 2.88 1.15 3.51 1.29 ;
 END
END RSDFFNSRASRNX2

MACRO RSDFFNSRASRQX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 31.04 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 24.225 0.59 24.595 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 29.455 1.435 29.795 1.8 ;
 RECT 27.775 1.99 29.64 2.13 ;
 RECT 25.545 2.22 27.915 2.36 ;
 RECT 27.775 1.435 27.915 1.99 ;
 RECT 29.5 1.8 29.64 1.99 ;
 RECT 25.545 1.39 25.685 2.22 ;
 RECT 26.93 1.37 27.07 2.22 ;
 RECT 27.775 2.13 27.915 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 5.155 0.08 5.435 0.295 ;
 RECT 27.895 0.08 28.135 0.26 ;
 RECT 9.085 0.31 9.375 0.45 ;
 RECT 16.695 0.275 17.72 0.415 ;
 RECT 12.77 0.59 13.045 0.73 ;
 RECT 17.58 0.75 18.525 0.89 ;
 RECT 0 -0.08 31.04 0.08 ;
 RECT 3.19 0.08 3.33 0.74 ;
 RECT 0.31 0.08 0.45 0.775 ;
 RECT 1.28 0.08 1.42 0.93 ;
 RECT 7.98 0.08 8.215 0.46 ;
 RECT 4.635 0.08 4.775 0.97 ;
 RECT 16.695 0.415 16.835 0.945 ;
 RECT 21.66 0.08 21.8 0.82 ;
 RECT 25.545 0.08 25.685 0.36 ;
 RECT 26.76 0.08 26.9 0.35 ;
 RECT 18.385 0.89 18.525 1.11 ;
 RECT 17.58 0.415 17.72 0.75 ;
 RECT 9.165 0.08 9.305 0.31 ;
 RECT 16.695 0.08 16.835 0.275 ;
 RECT 12.835 0.08 12.975 0.59 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 21.595 2.6 21.86 2.8 ;
 RECT 22.555 2.6 22.82 2.8 ;
 RECT 12.58 2.215 12.855 2.355 ;
 RECT 0 2.8 31.04 2.96 ;
 RECT 1.28 1.965 1.42 2.8 ;
 RECT 3.19 1.99 3.33 2.8 ;
 RECT 0.31 1.74 0.45 2.8 ;
 RECT 5.31 2.34 5.56 2.8 ;
 RECT 4.635 1.98 4.775 2.8 ;
 RECT 8.685 2.07 8.825 2.8 ;
 RECT 9.165 2.195 9.305 2.8 ;
 RECT 10.195 2.225 10.335 2.8 ;
 RECT 15.605 2.335 15.875 2.8 ;
 RECT 12.645 2.355 12.785 2.8 ;
 RECT 12.645 2.195 12.785 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.685 1.475 5.015 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.14 1.095 22.52 1.335 ;
 RECT 21.185 1.765 23.405 1.905 ;
 RECT 22.14 0.51 22.28 1.095 ;
 RECT 21.185 1.905 21.325 1.915 ;
 RECT 21.185 0.51 21.325 1.765 ;
 RECT 23.2 1.905 23.34 1.91 ;
 RECT 23.2 1.64 23.34 1.765 ;
 RECT 22.14 1.905 22.28 1.915 ;
 RECT 22.14 1.335 22.28 1.765 ;
 END
 ANTENNADIFFAREA 0.871 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.225 1.16 12.63 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.375 0.485 7.69 0.605 ;
 RECT 7.375 0.715 11.57 0.745 ;
 RECT 11.43 0.575 12.435 0.605 ;
 RECT 7.375 0.605 12.435 0.715 ;
 RECT 12.295 0.87 13.35 1.01 ;
 RECT 15.22 1.09 17.21 1.23 ;
 RECT 17.415 1.56 17.645 1.6 ;
 RECT 17.07 1.42 17.645 1.56 ;
 RECT 17.415 1.39 17.645 1.42 ;
 RECT 12.295 0.715 12.435 0.87 ;
 RECT 13.21 0.385 13.35 0.87 ;
 RECT 15.22 0.385 15.36 1.09 ;
 RECT 13.21 0.245 15.355 0.255 ;
 RECT 13.21 0.255 15.36 0.385 ;
 RECT 17.07 1.23 17.21 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.985 1.72 10.425 2.04 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.1 1.435 1.625 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.79 1.59 2.735 1.75 ;
 RECT 1.885 1.09 2.025 1.44 ;
 RECT 1.79 1.44 2.105 1.59 ;
 RECT 2.585 1.75 2.725 1.805 ;
 RECT 2.585 1.53 2.725 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.25 1.115 2.67 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 OBS
 LAYER PO ;
 RECT 25.675 1.035 25.905 1.245 ;
 RECT 15.915 0.105 18.74 0.205 ;
 RECT 15.915 0.205 16.015 1.91 ;
 RECT 18.64 0.205 18.74 1.265 ;
 RECT 15.095 1.71 15.195 1.91 ;
 RECT 14.01 1.61 15.195 1.71 ;
 RECT 14.01 0.475 14.11 1.61 ;
 RECT 14.56 1.71 14.66 2.425 ;
 RECT 10.675 0.475 10.775 0.895 ;
 RECT 15.095 1.91 16.015 2.01 ;
 RECT 10.675 0.375 14.11 0.475 ;
 RECT 10.55 0.895 10.78 1.105 ;
 RECT 16.225 0.455 18.155 0.535 ;
 RECT 17.925 0.535 18.155 0.6 ;
 RECT 17.925 0.39 18.155 0.435 ;
 RECT 16.305 0.435 18.155 0.455 ;
 RECT 16.225 0.535 16.455 0.665 ;
 RECT 17.08 0.535 17.31 0.835 ;
 RECT 17.08 0.835 17.18 2.39 ;
 RECT 26.11 0.215 26.21 0.995 ;
 RECT 26.11 0.995 26.35 1.205 ;
 RECT 26.11 1.205 26.21 2 ;
 RECT 28.505 0.375 28.605 0.99 ;
 RECT 28.505 0.99 28.755 1.2 ;
 RECT 28.505 1.2 28.605 2.27 ;
 RECT 28.505 2.27 28.79 2.48 ;
 RECT 13.49 0.655 13.59 2.305 ;
 RECT 13.795 2.3 14.025 2.305 ;
 RECT 13.795 2.405 14.025 2.51 ;
 RECT 13.49 2.305 14.025 2.405 ;
 RECT 25.33 0.21 25.43 0.755 ;
 RECT 25.33 0.855 25.43 2.2 ;
 RECT 28.195 1.125 28.295 2.2 ;
 RECT 24.365 0.755 25.9 0.84 ;
 RECT 24.365 0.84 25.895 0.855 ;
 RECT 25.8 0.215 25.9 0.755 ;
 RECT 24.365 0.595 24.595 0.755 ;
 RECT 25.33 2.2 28.295 2.3 ;
 RECT 12.2 1.28 12.455 1.45 ;
 RECT 12.2 1.45 12.3 1.655 ;
 RECT 12.2 0.655 12.3 1.18 ;
 RECT 12.2 1.655 13.16 1.755 ;
 RECT 13.06 1.755 13.16 2.355 ;
 RECT 11.285 0.66 11.385 1.18 ;
 RECT 12.2 1.755 12.3 2.51 ;
 RECT 11.285 1.24 12.455 1.28 ;
 RECT 11.285 1.18 12.3 1.24 ;
 RECT 27.02 0.38 27.12 0.96 ;
 RECT 27.02 1.06 27.12 1.14 ;
 RECT 26.6 0.935 26.83 0.96 ;
 RECT 26.6 0.96 27.12 1.06 ;
 RECT 26.6 1.06 26.83 1.145 ;
 RECT 27.02 1.14 27.29 1.24 ;
 RECT 27.19 1.24 27.29 1.84 ;
 RECT 27.385 0.22 27.615 0.28 ;
 RECT 27.385 0.38 27.615 0.43 ;
 RECT 27.02 0.28 27.615 0.38 ;
 RECT 11.275 1.575 11.375 2.485 ;
 RECT 11.785 1.575 12.015 1.685 ;
 RECT 11.275 1.475 12.015 1.575 ;
 RECT 29.205 0.195 29.305 2.665 ;
 RECT 28.195 0.095 29.305 0.195 ;
 RECT 24.57 1.245 24.67 2.665 ;
 RECT 28.195 0.195 28.295 0.945 ;
 RECT 24.57 1.2 24.855 1.245 ;
 RECT 24.625 1.035 24.855 1.1 ;
 RECT 24.57 2.665 29.305 2.765 ;
 RECT 24.57 1.1 24.9 1.2 ;
 RECT 15.5 0.795 15.665 0.925 ;
 RECT 14.82 0.885 15.05 0.925 ;
 RECT 14.82 1.025 15.05 1.095 ;
 RECT 14.82 0.925 15.665 1.025 ;
 RECT 15.5 0.585 15.73 0.795 ;
 RECT 2.535 1.55 2.775 1.78 ;
 RECT 2.675 1.78 2.775 2.695 ;
 RECT 1.065 1.435 1.635 1.71 ;
 RECT 1.065 0.515 1.165 1.435 ;
 RECT 1.065 1.71 1.165 2.645 ;
 RECT 1.535 0.515 1.635 1.435 ;
 RECT 1.535 1.71 1.635 2.695 ;
 RECT 2.255 1.37 2.355 1.605 ;
 RECT 2.485 0.515 2.585 1.14 ;
 RECT 2.205 1.705 2.305 2.695 ;
 RECT 2.205 1.605 2.355 1.705 ;
 RECT 2.255 1.14 2.585 1.37 ;
 RECT 1.87 0.515 1.97 1.105 ;
 RECT 1.83 1.105 2.075 1.345 ;
 RECT 4.42 0.52 4.52 2.465 ;
 RECT 4.18 0.27 4.52 0.52 ;
 RECT 7.05 1.33 7.19 1.475 ;
 RECT 7.05 1.71 7.15 2.475 ;
 RECT 7.09 0.65 7.19 1.33 ;
 RECT 7.05 1.475 7.28 1.71 ;
 RECT 6.6 0.705 6.7 1.165 ;
 RECT 6.16 1.27 6.26 1.445 ;
 RECT 6.6 0.47 6.885 0.705 ;
 RECT 6.16 1.17 6.7 1.265 ;
 RECT 6.16 1.265 6.535 1.27 ;
 RECT 6.39 1.165 6.7 1.17 ;
 RECT 6.015 1.445 6.26 1.69 ;
 RECT 7.49 0.715 7.59 1.61 ;
 RECT 7.525 1.71 7.625 2.48 ;
 RECT 7.49 1.61 7.625 1.71 ;
 RECT 7.37 0.485 7.61 0.715 ;
 RECT 13.095 0.655 13.195 1.24 ;
 RECT 12.965 1.24 13.195 1.475 ;
 RECT 4.895 0.49 4.995 1.495 ;
 RECT 4.7 1.495 4.995 1.745 ;
 RECT 4.895 1.745 4.995 2.37 ;
 RECT 2.975 0.135 3.075 0.22 ;
 RECT 2.815 0.22 3.075 0.43 ;
 RECT 2.975 0.43 3.075 2.695 ;
 RECT 3.445 0.295 3.545 1.115 ;
 RECT 3.28 1.115 3.545 1.325 ;
 RECT 3.445 1.325 3.545 2.74 ;
 RECT 19.52 0.77 19.62 2.155 ;
 RECT 19.52 0.55 19.62 0.56 ;
 RECT 19.52 0.56 19.775 0.77 ;
 RECT 20.155 0.43 20.255 1.245 ;
 RECT 20.105 1.245 20.335 1.455 ;
 RECT 20.09 0.22 20.32 0.43 ;
 RECT 8.31 2.445 8.57 2.655 ;
 RECT 8.47 1.79 8.57 2.445 ;
 RECT 18.58 1.445 18.68 2.035 ;
 RECT 18.565 2.035 18.795 2.245 ;
 RECT 19.05 0.55 19.15 2.69 ;
 RECT 9.98 1.58 10.08 1.72 ;
 RECT 9.72 1.01 9.82 1.48 ;
 RECT 9.98 1.93 10.08 2.69 ;
 RECT 9.98 1.72 10.215 1.93 ;
 RECT 9.72 1.48 10.08 1.58 ;
 RECT 9.98 2.69 19.15 2.79 ;
 RECT 9.42 0.98 9.52 1.615 ;
 RECT 9.28 1.615 9.52 1.825 ;
 RECT 9.42 1.825 9.52 2.68 ;
 RECT 21.92 0.355 22.02 1.33 ;
 RECT 20.73 1.33 23.08 1.43 ;
 RECT 22.98 1.43 23.08 2.695 ;
 RECT 22.4 1.43 22.5 2.69 ;
 RECT 21.44 0.385 21.54 1.33 ;
 RECT 21.44 1.43 21.54 2.69 ;
 RECT 20.73 1.25 20.96 1.33 ;
 RECT 20.73 1.43 20.96 1.46 ;
 RECT 21.92 1.43 22.02 2.69 ;
 RECT 21.92 0.255 23.815 0.355 ;
 RECT 23.585 0.22 23.815 0.255 ;
 RECT 23.585 0.355 23.815 0.43 ;
 RECT 17.55 0.73 17.65 1.39 ;
 RECT 17.415 1.39 17.65 1.6 ;
 RECT 17.55 1.6 17.65 2.39 ;
 RECT 5.735 0.285 5.835 1.52 ;
 RECT 5.235 1.52 5.835 1.62 ;
 RECT 5.735 0.185 14.625 0.195 ;
 RECT 7.79 0.095 14.625 0.185 ;
 RECT 5.735 0.195 7.89 0.285 ;
 RECT 14.525 0.195 14.625 1.29 ;
 RECT 15.42 1.39 15.615 1.405 ;
 RECT 6.555 1.565 6.655 2.675 ;
 RECT 5.67 1.62 5.77 2.675 ;
 RECT 5.235 1.44 5.48 1.52 ;
 RECT 5.235 1.62 5.48 1.69 ;
 RECT 7.79 0.285 7.89 1.24 ;
 RECT 14.525 1.29 15.615 1.39 ;
 RECT 5.67 2.675 6.655 2.775 ;
 RECT 15.42 1.405 15.65 1.615 ;
 RECT 25.805 1.245 25.905 2.02 ;
 LAYER CO ;
 RECT 0.315 1.825 0.445 1.955 ;
 RECT 17.805 1.035 17.935 1.165 ;
 RECT 18.39 0.91 18.52 1.04 ;
 RECT 10.2 2.3 10.33 2.43 ;
 RECT 2.865 0.26 2.995 0.39 ;
 RECT 3.33 1.155 3.46 1.285 ;
 RECT 20.78 1.29 20.91 1.42 ;
 RECT 20.155 1.285 20.285 1.415 ;
 RECT 17.975 0.43 18.105 0.56 ;
 RECT 19.595 0.6 19.725 0.73 ;
 RECT 20.14 0.26 20.27 0.39 ;
 RECT 8.36 2.485 8.49 2.615 ;
 RECT 18.615 2.075 18.745 2.205 ;
 RECT 10.035 1.76 10.165 1.89 ;
 RECT 9.33 1.655 9.46 1.785 ;
 RECT 23.635 0.26 23.765 0.39 ;
 RECT 28.575 1.03 28.705 1.16 ;
 RECT 16.275 0.495 16.405 0.625 ;
 RECT 17.465 1.43 17.595 1.56 ;
 RECT 15.55 0.625 15.68 0.755 ;
 RECT 15.47 1.445 15.6 1.575 ;
 RECT 25.725 1.075 25.855 1.205 ;
 RECT 10.6 0.935 10.73 1.065 ;
 RECT 26.65 0.975 26.78 1.105 ;
 RECT 17.13 0.665 17.26 0.795 ;
 RECT 26.17 1.035 26.3 1.165 ;
 RECT 28.61 2.31 28.74 2.44 ;
 RECT 13.845 2.34 13.975 2.47 ;
 RECT 24.415 0.635 24.545 0.765 ;
 RECT 12.275 1.28 12.405 1.41 ;
 RECT 27.435 0.26 27.565 0.39 ;
 RECT 11.835 1.515 11.965 1.645 ;
 RECT 24.675 1.075 24.805 1.205 ;
 RECT 14.87 0.925 15 1.055 ;
 RECT 4.76 1.55 4.89 1.68 ;
 RECT 21.66 2.64 21.79 2.77 ;
 RECT 21.19 0.655 21.32 0.785 ;
 RECT 21.19 1.725 21.32 1.855 ;
 RECT 1.285 0.735 1.415 0.865 ;
 RECT 1.29 1.51 1.42 1.64 ;
 RECT 0.815 0.735 0.945 0.865 ;
 RECT 3.195 2.31 3.325 2.44 ;
 RECT 1.285 2.015 1.415 2.145 ;
 RECT 1.89 1.155 2.02 1.285 ;
 RECT 3.195 2.05 3.325 2.18 ;
 RECT 2.59 1.6 2.72 1.73 ;
 RECT 3.665 2.01 3.795 2.14 ;
 RECT 3.665 0.735 3.795 0.865 ;
 RECT 2.425 2.075 2.555 2.205 ;
 RECT 1.285 2.275 1.415 2.405 ;
 RECT 3.195 0.545 3.325 0.675 ;
 RECT 3.665 1.75 3.795 1.88 ;
 RECT 0.815 2.015 0.945 2.145 ;
 RECT 2.23 0.735 2.36 0.865 ;
 RECT 2.41 1.19 2.54 1.32 ;
 RECT 28.725 0.595 28.855 0.725 ;
 RECT 7.1 1.525 7.23 1.655 ;
 RECT 12.65 2.225 12.78 2.355 ;
 RECT 22.62 2.64 22.75 2.77 ;
 RECT 4.17 2.115 4.3 2.245 ;
 RECT 27.27 0.595 27.4 0.725 ;
 RECT 6.705 0.525 6.835 0.655 ;
 RECT 7.75 1.825 7.88 1.955 ;
 RECT 27.78 1.49 27.91 1.62 ;
 RECT 6.35 0.88 6.48 1.01 ;
 RECT 14.78 1.87 14.91 2 ;
 RECT 8.22 2.11 8.35 2.24 ;
 RECT 8.035 0.32 8.165 0.45 ;
 RECT 25.55 0.135 25.68 0.265 ;
 RECT 5.295 1.495 5.425 1.625 ;
 RECT 5.245 0.745 5.375 0.875 ;
 RECT 5.115 1.995 5.245 2.125 ;
 RECT 11.95 1.995 12.08 2.125 ;
 RECT 0.315 0.59 0.445 0.72 ;
 RECT 11.505 2.07 11.635 2.2 ;
 RECT 14.275 0.595 14.405 0.725 ;
 RECT 6.07 1.49 6.2 1.62 ;
 RECT 13.015 1.28 13.145 1.41 ;
 RECT 22.145 1.725 22.275 1.855 ;
 RECT 0.315 2.085 0.445 2.215 ;
 RECT 9.71 2.235 9.84 2.365 ;
 RECT 21.665 0.62 21.795 0.75 ;
 RECT 8.69 2.135 8.82 2.265 ;
 RECT 6.305 2.105 6.435 2.235 ;
 RECT 7.27 2.11 7.4 2.24 ;
 RECT 5.225 0.145 5.355 0.275 ;
 RECT 14.275 1.9 14.405 2.03 ;
 RECT 0.315 2.345 0.445 2.475 ;
 RECT 5.38 2.345 5.51 2.475 ;
 RECT 26.33 0.435 26.46 0.565 ;
 RECT 9.98 1.23 10.11 1.36 ;
 RECT 18.8 1.705 18.93 1.835 ;
 RECT 9.17 2.265 9.3 2.395 ;
 RECT 6.82 0.88 6.95 1.01 ;
 RECT 16.83 1.835 16.96 1.965 ;
 RECT 16.7 0.765 16.83 0.895 ;
 RECT 4.64 0.74 4.77 0.87 ;
 RECT 27.945 0.12 28.075 0.25 ;
 RECT 7.425 0.53 7.555 0.66 ;
 RECT 22.145 0.62 22.275 0.75 ;
 RECT 15.675 2.38 15.805 2.51 ;
 RECT 11.95 0.885 12.08 1.015 ;
 RECT 25.08 1.425 25.21 1.555 ;
 RECT 0.315 0.33 0.445 0.46 ;
 RECT 19.865 0.92 19.995 1.05 ;
 RECT 25.55 1.475 25.68 1.605 ;
 RECT 13.75 0.875 13.88 1.005 ;
 RECT 5.955 0.79 6.085 0.92 ;
 RECT 17.77 1.835 17.9 1.965 ;
 RECT 6.8 2.07 6.93 2.2 ;
 RECT 29.505 1.475 29.635 1.605 ;
 RECT 23.205 1.71 23.335 1.84 ;
 RECT 4.17 0.74 4.3 0.87 ;
 RECT 5.89 1.825 6.02 1.955 ;
 RECT 13.75 1.945 13.88 2.075 ;
 RECT 4.64 2.05 4.77 2.18 ;
 RECT 24.83 0.505 24.96 0.635 ;
 RECT 11.025 2.015 11.155 2.145 ;
 RECT 26.765 0.12 26.895 0.25 ;
 RECT 26.33 1.485 26.46 1.615 ;
 RECT 28.725 1.465 28.855 1.595 ;
 RECT 19.27 1.705 19.4 1.835 ;
 RECT 19.745 1.705 19.875 1.835 ;
 RECT 27.41 1.405 27.54 1.535 ;
 RECT 11.03 0.905 11.16 1.035 ;
 RECT 4.24 0.325 4.37 0.455 ;
 RECT 9.17 0.315 9.3 0.445 ;
 RECT 11.505 0.905 11.635 1.035 ;
 RECT 14.78 0.595 14.91 0.725 ;
 RECT 12.84 0.595 12.97 0.725 ;
 RECT 26.935 1.445 27.065 1.575 ;
 LAYER M1 ;
 RECT 6.815 0.805 6.955 1.22 ;
 RECT 6.64 1.22 6.955 1.36 ;
 RECT 6.64 1.36 6.78 1.82 ;
 RECT 9.28 1.615 9.51 1.65 ;
 RECT 9.28 1.79 9.51 1.825 ;
 RECT 8.08 1.65 9.515 1.79 ;
 RECT 27.265 0.73 27.405 1.04 ;
 RECT 27.405 1.18 27.545 1.605 ;
 RECT 27.2 0.59 27.475 0.73 ;
 RECT 28.525 0.99 28.755 1.04 ;
 RECT 27.265 1.04 28.755 1.18 ;
 RECT 28.525 1.18 28.755 1.2 ;
 RECT 27.385 0.29 27.755 0.43 ;
 RECT 27.615 0.43 27.755 0.71 ;
 RECT 27.385 0.22 27.615 0.29 ;
 RECT 29.035 0.85 29.175 1.385 ;
 RECT 28.72 1.525 28.86 1.73 ;
 RECT 27.615 0.71 29.175 0.85 ;
 RECT 28.72 0.51 28.86 0.71 ;
 RECT 28.72 1.385 29.175 1.525 ;
 RECT 24.625 1.225 24.855 1.245 ;
 RECT 24.625 1.195 25.215 1.225 ;
 RECT 24.765 1.015 25.075 1.035 ;
 RECT 24.625 1.035 25.075 1.055 ;
 RECT 24.9 0.64 25.04 1.015 ;
 RECT 25.075 1.225 25.215 1.75 ;
 RECT 24.78 0.5 25.04 0.64 ;
 RECT 25.675 1.035 25.905 1.055 ;
 RECT 25.675 1.195 25.905 1.245 ;
 RECT 24.625 1.055 25.905 1.195 ;
 RECT 26.645 1.145 26.785 1.345 ;
 RECT 26.325 1.485 26.465 1.76 ;
 RECT 26.645 0.73 26.785 0.935 ;
 RECT 26.325 0.355 26.465 0.59 ;
 RECT 26.325 1.345 26.785 1.485 ;
 RECT 26.6 0.935 26.83 1.145 ;
 RECT 26.325 0.59 26.785 0.73 ;
 RECT 23.585 0.36 23.815 0.43 ;
 RECT 25.18 0.36 25.32 0.565 ;
 RECT 23.585 0.22 25.32 0.36 ;
 RECT 25.92 0.705 26.06 0.75 ;
 RECT 26.045 0.995 26.35 1.205 ;
 RECT 26.045 0.89 26.185 0.995 ;
 RECT 25.92 0.75 26.185 0.89 ;
 RECT 25.18 0.565 26.06 0.705 ;
 RECT 17.8 1.545 17.94 1.83 ;
 RECT 17.8 1.17 17.94 1.405 ;
 RECT 16.755 1.83 18.005 1.97 ;
 RECT 17.73 1.03 18.01 1.17 ;
 RECT 20.79 0.775 20.93 1.25 ;
 RECT 18.82 0.775 18.96 1.405 ;
 RECT 19.545 0.56 19.775 0.635 ;
 RECT 20.73 1.25 20.96 1.46 ;
 RECT 17.8 1.405 18.96 1.545 ;
 RECT 18.82 0.635 20.93 0.775 ;
 RECT 17.925 0.28 20.32 0.42 ;
 RECT 17.925 0.42 18.155 0.6 ;
 RECT 20.09 0.22 20.32 0.28 ;
 RECT 20.09 0.42 20.32 0.43 ;
 RECT 11.5 1.04 11.64 2.34 ;
 RECT 11.5 0.895 11.64 0.9 ;
 RECT 11.43 0.9 11.705 1.04 ;
 RECT 12.295 2.055 12.435 2.34 ;
 RECT 11.5 2.34 12.435 2.48 ;
 RECT 13.43 1.66 13.57 1.915 ;
 RECT 12.295 1.915 13.57 2.055 ;
 RECT 13.745 0.765 13.885 1.52 ;
 RECT 13.745 1.66 13.885 2.145 ;
 RECT 14.27 0.525 14.41 1.52 ;
 RECT 14.27 1.66 14.41 2.11 ;
 RECT 13.43 1.52 14.41 1.66 ;
 RECT 14.775 0.525 14.915 0.885 ;
 RECT 14.775 1.095 14.915 2.065 ;
 RECT 14.775 0.885 15.05 1.095 ;
 RECT 17.08 0.57 17.31 0.95 ;
 RECT 15.5 0.585 16.455 0.63 ;
 RECT 16.225 0.63 16.455 0.665 ;
 RECT 16.225 0.455 16.455 0.49 ;
 RECT 15.525 0.49 16.455 0.585 ;
 RECT 15.5 0.63 15.73 0.795 ;
 RECT 5.95 1.67 6.09 1.82 ;
 RECT 5.95 1.96 6.09 2.51 ;
 RECT 5.95 0.5 6.09 1.44 ;
 RECT 5.95 1.44 6.205 1.67 ;
 RECT 5.82 1.82 6.09 1.96 ;
 RECT 8.31 2.445 8.54 2.51 ;
 RECT 8.31 2.65 8.54 2.655 ;
 RECT 5.95 2.51 8.54 2.65 ;
 RECT 3.945 1.335 4.085 2.11 ;
 RECT 3.945 2.25 4.085 2.255 ;
 RECT 3.945 0.875 4.085 1.195 ;
 RECT 3.945 2.11 4.37 2.25 ;
 RECT 3.945 0.735 4.37 0.875 ;
 RECT 3.945 1.195 5.055 1.335 ;
 RECT 4.915 0.6 5.055 1.195 ;
 RECT 6.345 0.36 6.485 2.035 ;
 RECT 5.66 0.36 5.8 0.46 ;
 RECT 5.66 0.22 6.485 0.36 ;
 RECT 6.3 2.17 6.44 2.305 ;
 RECT 4.915 0.46 5.8 0.6 ;
 RECT 6.3 2.035 6.485 2.17 ;
 RECT 7.095 0.66 7.235 0.895 ;
 RECT 6.635 0.52 7.235 0.66 ;
 RECT 7.095 0.895 10.78 1.035 ;
 RECT 10.55 1.035 10.78 1.105 ;
 RECT 5.195 0.88 5.335 1.475 ;
 RECT 5.155 1.63 5.295 1.99 ;
 RECT 5.155 1.475 5.5 1.63 ;
 RECT 5.045 1.99 5.295 2.13 ;
 RECT 5.195 0.74 5.515 0.88 ;
 RECT 2.88 0.87 3.02 1.15 ;
 RECT 2.88 1.29 3.02 2.07 ;
 RECT 2.37 2.07 3.02 2.21 ;
 RECT 2.175 0.73 3.02 0.87 ;
 RECT 3.28 1.115 3.51 1.15 ;
 RECT 3.28 1.29 3.51 1.325 ;
 RECT 2.88 1.15 3.51 1.29 ;
 RECT 4.13 0.22 4.495 0.32 ;
 RECT 3.66 0.32 4.495 0.46 ;
 RECT 4.13 0.46 4.495 0.525 ;
 RECT 3.66 0.46 3.8 2.21 ;
 RECT 0.81 0.68 0.95 1.155 ;
 RECT 0.81 1.295 0.95 2.23 ;
 RECT 1.595 0.36 1.735 1.155 ;
 RECT 0.81 1.155 1.735 1.295 ;
 RECT 2.815 0.36 3.045 0.43 ;
 RECT 1.595 0.22 3.045 0.36 ;
 RECT 19.63 1.7 19.925 1.84 ;
 RECT 19.63 1.84 19.77 2.075 ;
 RECT 18.935 1.84 19.075 2.075 ;
 RECT 18.74 1.7 19.075 1.84 ;
 RECT 18.935 2.075 19.77 2.215 ;
 RECT 19.825 1.055 19.965 1.245 ;
 RECT 19.265 1.385 19.405 1.625 ;
 RECT 20.105 1.385 20.335 1.455 ;
 RECT 19.265 1.245 20.335 1.385 ;
 RECT 19.795 0.915 20.095 1.055 ;
 RECT 19.235 1.625 19.49 1.92 ;
 RECT 20.335 2.205 20.475 2.39 ;
 RECT 16.19 1.895 16.33 2.39 ;
 RECT 16.19 2.39 20.475 2.53 ;
 RECT 15.065 1.755 16.33 1.895 ;
 RECT 15.065 1.895 15.205 2.34 ;
 RECT 13.795 2.3 14.025 2.34 ;
 RECT 13.795 2.48 14.025 2.51 ;
 RECT 13.795 2.34 15.205 2.48 ;
 RECT 20.335 2.065 24.36 2.205 ;
 RECT 24.22 2.205 24.36 2.52 ;
 RECT 28.56 2.48 28.7 2.52 ;
 RECT 24.22 2.52 28.7 2.66 ;
 RECT 28.56 2.27 28.79 2.48 ;
 RECT 16.47 1.56 16.61 2.11 ;
 RECT 15.42 1.405 15.65 1.42 ;
 RECT 15.42 1.56 15.65 1.615 ;
 RECT 15.42 1.42 16.61 1.56 ;
 RECT 16.47 2.11 18.795 2.245 ;
 RECT 16.47 2.245 18.79 2.25 ;
 RECT 18.565 2.035 18.795 2.11 ;
 RECT 11.785 1.475 12.085 1.635 ;
 RECT 11.945 1.02 12.085 1.475 ;
 RECT 11.945 1.775 12.085 2.18 ;
 RECT 11.875 0.88 12.15 1.02 ;
 RECT 11.785 1.635 13.15 1.685 ;
 RECT 13.005 1.415 13.145 1.635 ;
 RECT 11.945 1.685 13.15 1.775 ;
 RECT 12.95 1.275 13.215 1.415 ;
 RECT 7.2 2.105 8.42 2.245 ;
 RECT 9.705 1.365 9.845 2.43 ;
 RECT 7.76 1.365 7.9 1.5 ;
 RECT 6.93 1.64 7.435 1.675 ;
 RECT 6.93 1.5 7.9 1.64 ;
 RECT 11.02 1.04 11.16 1.25 ;
 RECT 11.02 1.39 11.16 2.215 ;
 RECT 11.02 0.885 11.16 0.9 ;
 RECT 7.76 1.25 11.16 1.365 ;
 RECT 7.76 1.225 10.41 1.25 ;
 RECT 10.27 1.365 11.16 1.39 ;
 RECT 10.955 0.9 11.23 1.04 ;
 RECT 6.64 1.82 8.22 1.96 ;
 RECT 8.08 1.79 8.22 1.82 ;
 RECT 6.725 1.96 7.005 2.215 ;
 END
END RSDFFNSRASRQX1

MACRO RSDFFNSRASRQX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 32.64 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 25.92 0.59 26.29 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 31.15 1.435 31.49 1.8 ;
 RECT 29.47 1.99 31.335 2.13 ;
 RECT 27.24 2.22 29.61 2.36 ;
 RECT 29.47 1.435 29.61 1.99 ;
 RECT 31.195 1.8 31.335 1.99 ;
 RECT 27.24 1.39 27.38 2.22 ;
 RECT 28.625 1.37 28.765 2.22 ;
 RECT 29.47 2.13 29.61 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 5.145 0.08 5.425 0.295 ;
 RECT 29.59 0.08 29.83 0.26 ;
 RECT 9.075 0.31 9.365 0.45 ;
 RECT 12.76 0.59 13.03 0.73 ;
 RECT 16.685 0.275 17.71 0.415 ;
 RECT 17.57 0.75 18.515 0.89 ;
 RECT 0 -0.08 32.64 0.08 ;
 RECT 3.18 0.08 3.32 0.74 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 0.93 ;
 RECT 7.97 0.08 8.205 0.46 ;
 RECT 4.625 0.08 4.765 0.97 ;
 RECT 16.685 0.415 16.825 0.945 ;
 RECT 21.52 0.08 21.66 0.92 ;
 RECT 22.515 0.08 22.655 0.92 ;
 RECT 27.24 0.08 27.38 0.36 ;
 RECT 28.455 0.08 28.595 0.35 ;
 RECT 18.375 0.89 18.515 1.11 ;
 RECT 17.57 0.415 17.71 0.75 ;
 RECT 9.155 0.08 9.295 0.31 ;
 RECT 12.825 0.08 12.965 0.59 ;
 RECT 16.685 0.08 16.825 0.275 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 12.57 2.215 12.845 2.355 ;
 RECT 0 2.8 32.64 2.96 ;
 RECT 1.27 1.965 1.41 2.8 ;
 RECT 3.18 1.99 3.32 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 5.3 2.34 5.55 2.8 ;
 RECT 8.675 2.07 8.815 2.8 ;
 RECT 4.625 1.98 4.765 2.8 ;
 RECT 9.155 2.205 9.295 2.8 ;
 RECT 10.185 2.235 10.325 2.8 ;
 RECT 15.595 2.335 15.865 2.8 ;
 RECT 22.515 2.57 22.655 2.8 ;
 RECT 21.505 2.57 21.645 2.8 ;
 RECT 24.515 2.57 24.655 2.8 ;
 RECT 23.46 2.57 23.6 2.8 ;
 RECT 12.635 2.355 12.775 2.8 ;
 RECT 12.635 2.195 12.775 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.675 1.475 5.005 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.215 1.24 12.65 1.45 ;
 RECT 12.28 1.45 12.65 1.49 ;
 RECT 12.28 1.15 12.65 1.24 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.365 0.485 7.68 0.605 ;
 RECT 12.475 0.87 13.34 1.01 ;
 RECT 12.475 0.745 12.615 0.87 ;
 RECT 13.2 0.245 15.345 0.255 ;
 RECT 13.2 0.255 15.35 0.385 ;
 RECT 15.21 1.09 17.2 1.23 ;
 RECT 17.405 1.56 17.635 1.6 ;
 RECT 17.06 1.42 17.635 1.56 ;
 RECT 17.405 1.39 17.635 1.42 ;
 RECT 7.365 0.605 12.615 0.745 ;
 RECT 13.2 0.385 13.34 0.87 ;
 RECT 15.21 0.385 15.35 1.09 ;
 RECT 17.06 1.23 17.2 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.975 1.75 10.415 2.07 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.435 1.615 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.78 1.59 2.725 1.75 ;
 RECT 1.875 1.09 2.015 1.44 ;
 RECT 1.78 1.44 2.025 1.59 ;
 RECT 2.575 1.75 2.715 1.805 ;
 RECT 2.575 1.53 2.715 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.24 1.115 2.66 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.985 1.17 23.23 1.41 ;
 RECT 20.92 1.775 25.19 1.915 ;
 RECT 22.985 0.645 23.125 1.17 ;
 RECT 22.04 1.915 22.18 1.925 ;
 RECT 22.04 0.645 22.18 1.775 ;
 RECT 20.99 1.915 21.13 1.98 ;
 RECT 20.99 0.645 21.13 1.775 ;
 RECT 24.045 1.915 24.185 1.98 ;
 RECT 24.045 1.685 24.185 1.775 ;
 RECT 24.985 1.915 25.125 1.98 ;
 RECT 24.985 1.66 25.125 1.775 ;
 RECT 22.985 1.915 23.125 1.925 ;
 RECT 22.985 1.41 23.125 1.775 ;
 END
 ANTENNADIFFAREA 1.322 ;
 END Q

 OBS
 LAYER PO ;
 RECT 15.905 0.105 18.73 0.205 ;
 RECT 15.905 0.205 16.005 1.91 ;
 RECT 18.63 0.205 18.73 1.265 ;
 RECT 15.085 1.71 15.185 1.91 ;
 RECT 14 1.61 15.185 1.71 ;
 RECT 14 0.475 14.1 1.61 ;
 RECT 14.55 1.71 14.65 2.425 ;
 RECT 10.665 0.475 10.765 0.895 ;
 RECT 15.085 1.91 16.005 2.01 ;
 RECT 10.665 0.375 14.1 0.475 ;
 RECT 10.54 0.895 10.77 1.105 ;
 RECT 16.215 0.455 18.145 0.535 ;
 RECT 17.915 0.535 18.145 0.6 ;
 RECT 17.915 0.39 18.145 0.435 ;
 RECT 16.295 0.435 18.145 0.455 ;
 RECT 16.215 0.535 16.445 0.665 ;
 RECT 17.07 0.535 17.3 0.835 ;
 RECT 17.07 0.835 17.17 2.39 ;
 RECT 27.805 0.215 27.905 0.995 ;
 RECT 27.805 0.995 28.045 1.205 ;
 RECT 27.805 1.205 27.905 2 ;
 RECT 30.2 0.375 30.3 0.99 ;
 RECT 30.2 0.99 30.45 1.2 ;
 RECT 30.2 1.2 30.3 2.27 ;
 RECT 30.2 2.27 30.485 2.48 ;
 RECT 13.48 0.655 13.58 2.305 ;
 RECT 13.785 2.3 14.015 2.305 ;
 RECT 13.785 2.405 14.015 2.51 ;
 RECT 13.48 2.305 14.015 2.405 ;
 RECT 27.025 0.855 27.125 2.2 ;
 RECT 29.89 1.125 29.99 2.2 ;
 RECT 26.06 0.755 27.595 0.84 ;
 RECT 26.06 0.84 27.59 0.855 ;
 RECT 27.495 0.215 27.595 0.755 ;
 RECT 27.025 0.21 27.125 0.755 ;
 RECT 26.06 0.595 26.29 0.755 ;
 RECT 27.025 2.2 29.99 2.3 ;
 RECT 12.19 1.28 12.445 1.45 ;
 RECT 12.19 1.45 12.29 1.655 ;
 RECT 12.19 0.655 12.29 1.18 ;
 RECT 12.19 1.655 13.15 1.755 ;
 RECT 13.05 1.755 13.15 2.355 ;
 RECT 11.275 0.66 11.375 1.18 ;
 RECT 12.19 1.755 12.29 2.51 ;
 RECT 11.275 1.24 12.445 1.28 ;
 RECT 11.275 1.18 12.29 1.24 ;
 RECT 28.715 0.38 28.815 0.96 ;
 RECT 28.715 1.06 28.815 1.14 ;
 RECT 28.295 0.935 28.525 0.96 ;
 RECT 28.295 0.96 28.815 1.06 ;
 RECT 28.295 1.06 28.525 1.145 ;
 RECT 28.715 1.14 28.985 1.24 ;
 RECT 28.885 1.24 28.985 1.84 ;
 RECT 29.08 0.22 29.31 0.28 ;
 RECT 29.08 0.38 29.31 0.43 ;
 RECT 28.715 0.28 29.31 0.38 ;
 RECT 11.265 1.575 11.365 2.485 ;
 RECT 11.775 1.575 12.005 1.685 ;
 RECT 11.265 1.475 12.005 1.575 ;
 RECT 30.9 0.195 31 2.665 ;
 RECT 29.89 0.095 31 0.195 ;
 RECT 26.265 1.245 26.365 2.665 ;
 RECT 29.89 0.195 29.99 0.945 ;
 RECT 26.265 1.2 26.55 1.245 ;
 RECT 26.32 1.035 26.55 1.1 ;
 RECT 26.265 2.665 31 2.765 ;
 RECT 26.265 1.1 26.595 1.2 ;
 RECT 15.49 0.795 15.655 0.925 ;
 RECT 14.81 0.885 15.04 0.925 ;
 RECT 14.81 1.025 15.04 1.095 ;
 RECT 14.81 0.925 15.655 1.025 ;
 RECT 15.49 0.585 15.72 0.795 ;
 RECT 2.525 1.55 2.765 1.78 ;
 RECT 2.665 1.78 2.765 2.695 ;
 RECT 1.055 1.435 1.625 1.71 ;
 RECT 1.055 0.515 1.155 1.435 ;
 RECT 1.055 1.71 1.155 2.645 ;
 RECT 1.525 0.515 1.625 1.435 ;
 RECT 1.525 1.71 1.625 2.695 ;
 RECT 2.245 1.37 2.345 1.605 ;
 RECT 2.475 0.515 2.575 1.14 ;
 RECT 2.195 1.705 2.295 2.695 ;
 RECT 2.195 1.605 2.345 1.705 ;
 RECT 2.245 1.14 2.575 1.37 ;
 RECT 1.86 0.515 1.96 1.105 ;
 RECT 1.82 1.105 2.065 1.345 ;
 RECT 4.41 0.52 4.51 2.465 ;
 RECT 4.17 0.27 4.51 0.52 ;
 RECT 7.04 1.33 7.18 1.475 ;
 RECT 7.04 1.71 7.14 2.475 ;
 RECT 7.08 0.65 7.18 1.33 ;
 RECT 7.04 1.475 7.27 1.71 ;
 RECT 6.59 0.705 6.69 1.165 ;
 RECT 6.15 1.27 6.25 1.445 ;
 RECT 6.59 0.47 6.875 0.705 ;
 RECT 6.15 1.17 6.69 1.265 ;
 RECT 6.15 1.265 6.525 1.27 ;
 RECT 6.38 1.165 6.69 1.17 ;
 RECT 6.005 1.445 6.25 1.69 ;
 RECT 7.48 0.715 7.58 1.61 ;
 RECT 7.515 1.71 7.615 2.48 ;
 RECT 7.48 1.61 7.615 1.71 ;
 RECT 7.36 0.485 7.6 0.715 ;
 RECT 13.085 0.655 13.185 1.24 ;
 RECT 12.955 1.24 13.185 1.475 ;
 RECT 4.885 0.49 4.985 1.495 ;
 RECT 4.69 1.495 4.985 1.745 ;
 RECT 4.885 1.745 4.985 2.37 ;
 RECT 2.8 0.245 3.065 0.455 ;
 RECT 2.965 0.455 3.065 2.695 ;
 RECT 3.435 0.295 3.535 1.115 ;
 RECT 3.245 1.115 3.535 1.325 ;
 RECT 3.435 1.325 3.535 2.765 ;
 RECT 19.51 0.77 19.61 2.155 ;
 RECT 19.51 0.55 19.61 0.56 ;
 RECT 19.51 0.56 19.765 0.77 ;
 RECT 20.145 0.43 20.245 1.245 ;
 RECT 20.095 1.245 20.325 1.455 ;
 RECT 20.145 0.22 20.375 0.43 ;
 RECT 8.3 2.445 8.56 2.655 ;
 RECT 8.46 1.79 8.56 2.445 ;
 RECT 18.57 1.445 18.67 2.035 ;
 RECT 18.555 2.035 18.785 2.245 ;
 RECT 19.04 0.55 19.14 2.69 ;
 RECT 9.97 1.58 10.07 1.76 ;
 RECT 9.71 1.01 9.81 1.48 ;
 RECT 9.97 1.97 10.07 2.69 ;
 RECT 9.97 1.76 10.205 1.97 ;
 RECT 9.71 1.48 10.07 1.58 ;
 RECT 9.97 2.69 19.14 2.79 ;
 RECT 9.41 0.98 9.51 1.615 ;
 RECT 9.27 1.615 9.51 1.825 ;
 RECT 9.41 1.825 9.51 2.695 ;
 RECT 20.595 1.295 24.87 1.395 ;
 RECT 21.825 0.375 21.925 1.295 ;
 RECT 21.825 1.395 21.925 2.715 ;
 RECT 22.77 0.325 22.87 1.295 ;
 RECT 21.245 0.375 21.345 1.295 ;
 RECT 21.245 1.395 21.345 2.69 ;
 RECT 24.77 1.395 24.87 2.685 ;
 RECT 20.595 1.26 20.825 1.295 ;
 RECT 20.595 1.395 20.825 1.47 ;
 RECT 22.3 0.405 22.4 1.295 ;
 RECT 22.3 1.395 22.4 2.69 ;
 RECT 23.825 1.395 23.925 2.715 ;
 RECT 23.245 1.395 23.345 2.69 ;
 RECT 24.3 1.395 24.4 2.69 ;
 RECT 22.77 1.395 22.87 2.685 ;
 RECT 22.77 0.225 25.51 0.325 ;
 RECT 25.28 0.22 25.51 0.225 ;
 RECT 25.28 0.325 25.51 0.43 ;
 RECT 17.54 0.73 17.64 1.39 ;
 RECT 17.405 1.39 17.64 1.6 ;
 RECT 17.54 1.6 17.64 2.39 ;
 RECT 5.725 0.285 5.825 1.52 ;
 RECT 5.225 1.52 5.825 1.62 ;
 RECT 5.725 0.185 14.615 0.195 ;
 RECT 7.78 0.095 14.615 0.185 ;
 RECT 5.725 0.195 7.88 0.285 ;
 RECT 14.515 0.195 14.615 1.29 ;
 RECT 15.41 1.39 15.605 1.405 ;
 RECT 6.545 1.565 6.645 2.675 ;
 RECT 5.66 1.62 5.76 2.675 ;
 RECT 5.225 1.44 5.47 1.52 ;
 RECT 5.225 1.62 5.47 1.69 ;
 RECT 7.78 0.285 7.88 1.24 ;
 RECT 14.515 1.29 15.605 1.39 ;
 RECT 5.66 2.675 6.645 2.775 ;
 RECT 15.41 1.405 15.64 1.615 ;
 RECT 27.5 1.245 27.6 2.02 ;
 RECT 27.37 1.035 27.6 1.245 ;
 LAYER CO ;
 RECT 20.645 1.3 20.775 1.43 ;
 RECT 20.145 1.285 20.275 1.415 ;
 RECT 17.965 0.43 18.095 0.56 ;
 RECT 19.585 0.6 19.715 0.73 ;
 RECT 20.195 0.26 20.325 0.39 ;
 RECT 8.35 2.485 8.48 2.615 ;
 RECT 18.605 2.075 18.735 2.205 ;
 RECT 10.025 1.8 10.155 1.93 ;
 RECT 9.32 1.655 9.45 1.785 ;
 RECT 25.33 0.26 25.46 0.39 ;
 RECT 30.27 1.03 30.4 1.16 ;
 RECT 16.265 0.495 16.395 0.625 ;
 RECT 17.455 1.43 17.585 1.56 ;
 RECT 15.54 0.625 15.67 0.755 ;
 RECT 15.46 1.445 15.59 1.575 ;
 RECT 27.42 1.075 27.55 1.205 ;
 RECT 10.59 0.935 10.72 1.065 ;
 RECT 28.345 0.975 28.475 1.105 ;
 RECT 17.12 0.665 17.25 0.795 ;
 RECT 27.865 1.035 27.995 1.165 ;
 RECT 30.305 2.31 30.435 2.44 ;
 RECT 13.835 2.34 13.965 2.47 ;
 RECT 26.11 0.635 26.24 0.765 ;
 RECT 12.265 1.28 12.395 1.41 ;
 RECT 29.13 0.26 29.26 0.39 ;
 RECT 11.825 1.515 11.955 1.645 ;
 RECT 26.37 1.075 26.5 1.205 ;
 RECT 14.86 0.925 14.99 1.055 ;
 RECT 4.75 1.55 4.88 1.68 ;
 RECT 21.51 2.64 21.64 2.77 ;
 RECT 22.52 2.64 22.65 2.77 ;
 RECT 22.52 0.72 22.65 0.85 ;
 RECT 21.525 0.72 21.655 0.85 ;
 RECT 22.045 0.72 22.175 0.85 ;
 RECT 20.995 0.72 21.125 0.85 ;
 RECT 20.995 1.78 21.125 1.91 ;
 RECT 22.045 1.78 22.175 1.91 ;
 RECT 1.275 0.735 1.405 0.865 ;
 RECT 1.28 1.51 1.41 1.64 ;
 RECT 0.805 0.735 0.935 0.865 ;
 RECT 3.185 2.31 3.315 2.44 ;
 RECT 1.275 2.015 1.405 2.145 ;
 RECT 1.88 1.155 2.01 1.285 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 2.58 1.6 2.71 1.73 ;
 RECT 3.655 2.01 3.785 2.14 ;
 RECT 3.655 0.735 3.785 0.865 ;
 RECT 2.415 2.075 2.545 2.205 ;
 RECT 1.275 2.275 1.405 2.405 ;
 RECT 3.185 0.545 3.315 0.675 ;
 RECT 3.655 1.75 3.785 1.88 ;
 RECT 0.805 2.015 0.935 2.145 ;
 RECT 2.22 0.735 2.35 0.865 ;
 RECT 2.4 1.19 2.53 1.32 ;
 RECT 28.965 0.595 29.095 0.725 ;
 RECT 6.695 0.525 6.825 0.655 ;
 RECT 7.74 1.825 7.87 1.955 ;
 RECT 29.475 1.49 29.605 1.62 ;
 RECT 6.34 0.88 6.47 1.01 ;
 RECT 14.77 1.87 14.9 2 ;
 RECT 8.21 2.11 8.34 2.24 ;
 RECT 8.025 0.32 8.155 0.45 ;
 RECT 27.245 0.135 27.375 0.265 ;
 RECT 5.285 1.495 5.415 1.625 ;
 RECT 5.235 0.745 5.365 0.875 ;
 RECT 5.105 1.995 5.235 2.125 ;
 RECT 11.94 1.995 12.07 2.125 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 11.495 2.07 11.625 2.2 ;
 RECT 14.265 0.595 14.395 0.725 ;
 RECT 6.06 1.49 6.19 1.62 ;
 RECT 13.005 1.28 13.135 1.41 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 24.52 2.64 24.65 2.77 ;
 RECT 24.05 1.78 24.18 1.91 ;
 RECT 22.99 1.735 23.12 1.865 ;
 RECT 23.465 2.64 23.595 2.77 ;
 RECT 24.99 1.78 25.12 1.91 ;
 RECT 22.99 0.72 23.12 0.85 ;
 RECT 9.7 2.24 9.83 2.37 ;
 RECT 8.68 2.135 8.81 2.265 ;
 RECT 6.295 2.105 6.425 2.235 ;
 RECT 7.26 2.11 7.39 2.24 ;
 RECT 5.215 0.145 5.345 0.275 ;
 RECT 14.265 1.9 14.395 2.03 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 5.37 2.345 5.5 2.475 ;
 RECT 28.025 0.435 28.155 0.565 ;
 RECT 9.97 1.23 10.1 1.36 ;
 RECT 18.79 1.705 18.92 1.835 ;
 RECT 9.16 2.27 9.29 2.4 ;
 RECT 6.81 0.88 6.94 1.01 ;
 RECT 16.82 1.835 16.95 1.965 ;
 RECT 16.69 0.765 16.82 0.895 ;
 RECT 4.63 0.74 4.76 0.87 ;
 RECT 29.64 0.12 29.77 0.25 ;
 RECT 7.415 0.53 7.545 0.66 ;
 RECT 15.665 2.38 15.795 2.51 ;
 RECT 11.94 0.905 12.07 1.035 ;
 RECT 26.775 1.425 26.905 1.555 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 19.855 0.92 19.985 1.05 ;
 RECT 27.245 1.475 27.375 1.605 ;
 RECT 13.74 0.875 13.87 1.005 ;
 RECT 5.945 0.79 6.075 0.92 ;
 RECT 17.76 1.835 17.89 1.965 ;
 RECT 6.79 2.07 6.92 2.2 ;
 RECT 31.2 1.475 31.33 1.605 ;
 RECT 4.16 0.74 4.29 0.87 ;
 RECT 5.88 1.825 6.01 1.955 ;
 RECT 13.74 1.945 13.87 2.075 ;
 RECT 4.63 2.05 4.76 2.18 ;
 RECT 26.525 0.505 26.655 0.635 ;
 RECT 11.015 2.015 11.145 2.145 ;
 RECT 28.46 0.12 28.59 0.25 ;
 RECT 28.025 1.485 28.155 1.615 ;
 RECT 30.42 1.465 30.55 1.595 ;
 RECT 19.26 1.705 19.39 1.835 ;
 RECT 30.42 0.595 30.55 0.725 ;
 RECT 7.09 1.525 7.22 1.655 ;
 RECT 12.64 2.225 12.77 2.355 ;
 RECT 4.16 2.115 4.29 2.245 ;
 RECT 19.735 1.705 19.865 1.835 ;
 RECT 29.105 1.405 29.235 1.535 ;
 RECT 11.02 0.905 11.15 1.035 ;
 RECT 4.23 0.325 4.36 0.455 ;
 RECT 9.16 0.315 9.29 0.445 ;
 RECT 11.495 0.905 11.625 1.035 ;
 RECT 14.77 0.595 14.9 0.725 ;
 RECT 12.83 0.595 12.96 0.725 ;
 RECT 28.63 1.445 28.76 1.575 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 17.795 1.035 17.925 1.165 ;
 RECT 18.38 0.91 18.51 1.04 ;
 RECT 10.19 2.305 10.32 2.435 ;
 RECT 2.85 0.285 2.98 0.415 ;
 RECT 3.295 1.155 3.425 1.285 ;
 LAYER M1 ;
 RECT 28.02 0.355 28.16 0.59 ;
 RECT 28.02 1.345 28.48 1.485 ;
 RECT 28.295 0.935 28.525 1.145 ;
 RECT 28.02 0.59 28.48 0.73 ;
 RECT 28.96 0.73 29.1 1.04 ;
 RECT 29.1 1.18 29.24 1.605 ;
 RECT 28.895 0.59 29.17 0.73 ;
 RECT 30.22 0.99 30.45 1.04 ;
 RECT 28.96 1.04 30.45 1.18 ;
 RECT 30.22 1.18 30.45 1.2 ;
 RECT 29.08 0.29 29.45 0.43 ;
 RECT 29.31 0.43 29.45 0.71 ;
 RECT 29.08 0.22 29.31 0.29 ;
 RECT 30.73 0.85 30.87 1.385 ;
 RECT 30.415 1.525 30.555 1.73 ;
 RECT 29.31 0.71 30.87 0.85 ;
 RECT 30.415 0.51 30.555 0.71 ;
 RECT 30.415 1.385 30.87 1.525 ;
 RECT 26.32 1.225 26.55 1.245 ;
 RECT 26.32 1.195 26.91 1.225 ;
 RECT 26.46 1.015 26.77 1.035 ;
 RECT 26.32 1.035 26.77 1.055 ;
 RECT 26.595 0.64 26.735 1.015 ;
 RECT 26.77 1.225 26.91 1.75 ;
 RECT 26.475 0.5 26.735 0.64 ;
 RECT 27.37 1.035 27.6 1.055 ;
 RECT 27.37 1.195 27.6 1.245 ;
 RECT 26.32 1.055 27.6 1.195 ;
 RECT 25.28 0.36 25.51 0.43 ;
 RECT 26.875 0.36 27.015 0.565 ;
 RECT 25.28 0.22 27.015 0.36 ;
 RECT 27.615 0.705 27.755 0.75 ;
 RECT 27.74 0.995 28.045 1.205 ;
 RECT 27.74 0.89 27.88 0.995 ;
 RECT 27.615 0.75 27.88 0.89 ;
 RECT 26.875 0.565 27.755 0.705 ;
 RECT 17.79 1.545 17.93 1.83 ;
 RECT 16.745 1.83 17.995 1.97 ;
 RECT 17.79 1.17 17.93 1.405 ;
 RECT 17.72 1.03 18 1.17 ;
 RECT 20.51 1.26 20.825 1.42 ;
 RECT 20.51 0.775 20.65 1.26 ;
 RECT 20.595 1.42 20.825 1.47 ;
 RECT 18.81 0.775 18.95 1.405 ;
 RECT 19.535 0.56 19.765 0.635 ;
 RECT 17.79 1.405 18.95 1.545 ;
 RECT 18.81 0.635 20.65 0.775 ;
 RECT 11.49 1.04 11.63 2.34 ;
 RECT 11.49 0.895 11.63 0.9 ;
 RECT 11.42 0.9 11.695 1.04 ;
 RECT 12.285 2.055 12.425 2.34 ;
 RECT 11.49 2.34 12.425 2.48 ;
 RECT 13.42 1.66 13.56 1.915 ;
 RECT 12.285 1.915 13.56 2.055 ;
 RECT 13.735 0.765 13.875 1.52 ;
 RECT 13.735 1.66 13.875 2.145 ;
 RECT 14.26 0.525 14.4 1.52 ;
 RECT 14.26 1.66 14.4 2.11 ;
 RECT 13.42 1.52 14.4 1.66 ;
 RECT 14.765 0.525 14.905 0.885 ;
 RECT 14.765 1.095 14.905 2.065 ;
 RECT 14.765 0.885 15.04 1.095 ;
 RECT 17.07 0.57 17.3 0.95 ;
 RECT 20.145 0.22 20.375 0.28 ;
 RECT 20.145 0.42 20.375 0.43 ;
 RECT 17.915 0.28 20.375 0.42 ;
 RECT 17.915 0.42 18.145 0.6 ;
 RECT 15.49 0.585 16.445 0.63 ;
 RECT 16.215 0.63 16.445 0.665 ;
 RECT 16.215 0.455 16.445 0.49 ;
 RECT 15.515 0.49 16.445 0.585 ;
 RECT 15.49 0.63 15.72 0.795 ;
 RECT 5.94 1.67 6.08 1.82 ;
 RECT 5.94 1.96 6.08 2.51 ;
 RECT 5.94 0.5 6.08 1.44 ;
 RECT 5.94 1.44 6.195 1.67 ;
 RECT 5.81 1.82 6.08 1.96 ;
 RECT 8.3 2.445 8.53 2.51 ;
 RECT 8.3 2.65 8.53 2.655 ;
 RECT 5.94 2.51 8.53 2.65 ;
 RECT 3.935 0.875 4.075 1.195 ;
 RECT 3.935 1.335 4.075 2.11 ;
 RECT 3.935 2.25 4.075 2.255 ;
 RECT 3.935 0.735 4.36 0.875 ;
 RECT 3.935 2.11 4.36 2.25 ;
 RECT 3.935 1.195 5.045 1.335 ;
 RECT 4.905 0.6 5.045 1.195 ;
 RECT 6.335 0.36 6.475 2.035 ;
 RECT 5.65 0.36 5.79 0.46 ;
 RECT 5.65 0.22 6.475 0.36 ;
 RECT 6.29 2.17 6.43 2.305 ;
 RECT 4.905 0.46 5.79 0.6 ;
 RECT 6.29 2.035 6.475 2.17 ;
 RECT 7.085 0.66 7.225 0.895 ;
 RECT 6.625 0.52 7.225 0.66 ;
 RECT 7.085 0.895 10.77 1.035 ;
 RECT 10.54 1.035 10.77 1.105 ;
 RECT 2.87 0.87 3.01 1.15 ;
 RECT 2.87 1.29 3.01 2.07 ;
 RECT 2.36 2.07 3.01 2.21 ;
 RECT 2.165 0.73 3.01 0.87 ;
 RECT 3.245 1.115 3.475 1.15 ;
 RECT 3.245 1.29 3.475 1.325 ;
 RECT 2.87 1.15 3.475 1.29 ;
 RECT 4.12 0.22 4.485 0.32 ;
 RECT 3.65 0.32 4.485 0.46 ;
 RECT 4.12 0.46 4.485 0.525 ;
 RECT 3.65 0.46 3.79 2.21 ;
 RECT 0.8 0.68 0.94 1.155 ;
 RECT 0.8 1.295 0.94 2.23 ;
 RECT 1.585 0.385 1.725 1.155 ;
 RECT 0.8 1.155 1.725 1.295 ;
 RECT 2.8 0.385 3.03 0.455 ;
 RECT 1.585 0.245 3.03 0.385 ;
 RECT 16.18 1.895 16.32 2.39 ;
 RECT 16.18 2.415 20.465 2.53 ;
 RECT 15.055 1.755 16.32 1.895 ;
 RECT 15.055 1.895 15.195 2.34 ;
 RECT 13.785 2.3 14.015 2.34 ;
 RECT 13.785 2.48 14.015 2.51 ;
 RECT 13.785 2.34 15.195 2.48 ;
 RECT 25.915 2.415 26.055 2.52 ;
 RECT 16.18 2.39 26.055 2.415 ;
 RECT 20.325 2.275 26.055 2.39 ;
 RECT 30.255 2.48 30.395 2.52 ;
 RECT 25.915 2.52 30.395 2.66 ;
 RECT 30.255 2.27 30.485 2.48 ;
 RECT 19.62 1.7 19.915 1.84 ;
 RECT 19.62 1.84 19.76 2.075 ;
 RECT 18.925 1.84 19.065 2.075 ;
 RECT 18.73 1.7 19.065 1.84 ;
 RECT 18.925 2.075 19.76 2.215 ;
 RECT 19.815 1.055 19.955 1.245 ;
 RECT 19.255 1.385 19.395 1.625 ;
 RECT 20.095 1.385 20.325 1.455 ;
 RECT 19.255 1.245 20.325 1.385 ;
 RECT 19.785 0.915 20.085 1.055 ;
 RECT 19.225 1.625 19.48 1.92 ;
 RECT 16.46 1.56 16.6 2.11 ;
 RECT 15.41 1.405 15.64 1.42 ;
 RECT 15.41 1.56 15.64 1.615 ;
 RECT 15.41 1.42 16.6 1.56 ;
 RECT 16.46 2.11 18.785 2.245 ;
 RECT 16.46 2.245 18.78 2.25 ;
 RECT 18.555 2.035 18.785 2.11 ;
 RECT 11.935 1.04 12.075 1.475 ;
 RECT 11.775 1.475 12.075 1.635 ;
 RECT 11.935 1.775 12.075 2.18 ;
 RECT 11.865 0.9 12.14 1.04 ;
 RECT 11.935 1.685 13.15 1.775 ;
 RECT 13.01 1.415 13.15 1.635 ;
 RECT 11.775 1.635 13.15 1.685 ;
 RECT 12.945 1.275 13.205 1.415 ;
 RECT 7.19 2.105 8.41 2.245 ;
 RECT 9.695 1.365 9.835 2.435 ;
 RECT 7.75 1.365 7.89 1.5 ;
 RECT 6.92 1.64 7.425 1.675 ;
 RECT 6.92 1.5 7.89 1.64 ;
 RECT 11.01 1.04 11.15 1.25 ;
 RECT 11.01 1.39 11.15 2.215 ;
 RECT 11.01 0.885 11.15 0.9 ;
 RECT 7.75 1.25 11.15 1.365 ;
 RECT 7.75 1.225 10.4 1.25 ;
 RECT 10.26 1.365 11.15 1.39 ;
 RECT 10.945 0.9 11.22 1.04 ;
 RECT 5.145 1.475 5.49 1.63 ;
 RECT 5.145 1.63 5.285 1.99 ;
 RECT 5.185 0.88 5.325 1.475 ;
 RECT 5.035 1.99 5.285 2.13 ;
 RECT 5.185 0.74 5.505 0.88 ;
 RECT 6.63 1.82 8.21 1.96 ;
 RECT 8.07 1.79 8.21 1.82 ;
 RECT 6.715 1.96 6.995 2.215 ;
 RECT 6.805 0.805 6.945 1.22 ;
 RECT 6.63 1.22 6.945 1.36 ;
 RECT 6.63 1.36 6.77 1.82 ;
 RECT 9.27 1.615 9.5 1.65 ;
 RECT 9.27 1.79 9.5 1.825 ;
 RECT 8.07 1.65 9.505 1.79 ;
 RECT 28.34 1.145 28.48 1.345 ;
 RECT 28.02 1.485 28.16 1.76 ;
 RECT 28.34 0.73 28.48 0.935 ;
 END
END RSDFFNSRASRQX2

MACRO RSDFFNSRASRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 31.04 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 24.225 0.59 24.595 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 29.455 1.435 29.795 1.8 ;
 RECT 27.775 1.99 29.64 2.13 ;
 RECT 25.545 2.22 27.915 2.36 ;
 RECT 27.775 1.435 27.915 1.99 ;
 RECT 29.5 1.8 29.64 1.99 ;
 RECT 25.545 1.39 25.685 2.22 ;
 RECT 26.93 1.37 27.07 2.22 ;
 RECT 27.775 2.13 27.915 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 5.155 0.08 5.435 0.295 ;
 RECT 27.895 0.08 28.135 0.26 ;
 RECT 12.765 0.595 13.04 0.735 ;
 RECT 9.085 0.31 9.375 0.45 ;
 RECT 16.695 0.275 17.72 0.415 ;
 RECT 21.055 0.335 21.32 0.495 ;
 RECT 17.58 0.75 18.525 0.89 ;
 RECT 0 -0.08 31.04 0.08 ;
 RECT 3.19 0.08 3.33 0.74 ;
 RECT 0.31 0.08 0.45 0.775 ;
 RECT 1.28 0.08 1.42 0.93 ;
 RECT 7.98 0.08 8.215 0.46 ;
 RECT 4.635 0.08 4.775 0.97 ;
 RECT 16.695 0.415 16.835 0.945 ;
 RECT 22.7 0.08 22.84 0.82 ;
 RECT 25.545 0.08 25.685 0.36 ;
 RECT 26.76 0.08 26.9 0.35 ;
 RECT 18.385 0.89 18.525 1.11 ;
 RECT 17.58 0.415 17.72 0.75 ;
 RECT 12.835 0.08 12.975 0.595 ;
 RECT 9.165 0.08 9.305 0.31 ;
 RECT 16.695 0.08 16.835 0.275 ;
 RECT 21.11 0.08 21.25 0.335 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.51 1.205 20.845 1.445 ;
 RECT 20.62 0.915 20.76 1.205 ;
 RECT 21.625 1.84 21.765 1.885 ;
 RECT 21.625 0.915 21.765 1.7 ;
 RECT 20.62 1.84 20.76 1.885 ;
 RECT 20.62 1.7 21.765 1.84 ;
 RECT 20.62 1.445 20.76 1.7 ;
 END
 ANTENNADIFFAREA 0.433 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 20.965 2.6 21.23 2.8 ;
 RECT 22.555 2.6 22.82 2.8 ;
 RECT 12.58 2.215 12.855 2.355 ;
 RECT 0 2.8 31.04 2.96 ;
 RECT 1.28 1.965 1.42 2.8 ;
 RECT 3.19 1.99 3.33 2.8 ;
 RECT 0.31 1.74 0.45 2.8 ;
 RECT 5.31 2.34 5.56 2.8 ;
 RECT 4.635 1.98 4.775 2.8 ;
 RECT 12.645 2.195 12.785 2.215 ;
 RECT 8.685 2.07 8.825 2.8 ;
 RECT 9.165 1.98 9.305 2.8 ;
 RECT 10.195 2.35 10.335 2.8 ;
 RECT 15.605 2.335 15.875 2.8 ;
 RECT 12.645 2.355 12.785 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.685 1.475 5.015 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.02 1.095 22.28 1.335 ;
 RECT 22.14 0.51 22.28 1.095 ;
 RECT 23.2 1.905 23.34 1.91 ;
 RECT 22.14 1.765 23.34 1.905 ;
 RECT 23.2 0.56 23.34 1.765 ;
 RECT 22.14 1.905 22.28 1.915 ;
 RECT 22.14 1.335 22.28 1.765 ;
 END
 ANTENNADIFFAREA 0.73 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.245 1.16 12.61 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.375 0.485 7.69 0.6 ;
 RECT 12.485 0.875 13.35 1.015 ;
 RECT 13.21 0.245 15.355 0.255 ;
 RECT 13.21 0.255 15.36 0.385 ;
 RECT 15.22 1.09 17.21 1.23 ;
 RECT 17.415 1.56 17.645 1.6 ;
 RECT 17.07 1.42 17.645 1.56 ;
 RECT 17.415 1.39 17.645 1.42 ;
 RECT 11.585 0.535 12.625 0.6 ;
 RECT 7.375 0.675 11.725 0.74 ;
 RECT 7.375 0.6 12.625 0.675 ;
 RECT 12.485 0.675 12.625 0.875 ;
 RECT 13.21 0.385 13.35 0.875 ;
 RECT 15.22 0.385 15.36 1.09 ;
 RECT 17.07 1.23 17.21 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.985 1.615 10.355 2.03 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.1 1.435 1.625 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.79 1.59 2.735 1.75 ;
 RECT 1.885 1.09 2.025 1.44 ;
 RECT 1.79 1.44 2.035 1.59 ;
 RECT 2.585 1.75 2.725 1.805 ;
 RECT 2.585 1.53 2.725 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.25 1.115 2.67 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 OBS
 LAYER PO ;
 RECT 25.805 1.245 25.905 2.02 ;
 RECT 25.675 1.035 25.905 1.245 ;
 RECT 15.915 0.105 18.74 0.205 ;
 RECT 15.915 0.205 16.015 1.91 ;
 RECT 18.64 0.205 18.74 1.265 ;
 RECT 15.095 1.71 15.195 1.91 ;
 RECT 14.01 1.61 15.195 1.71 ;
 RECT 14.01 0.475 14.11 1.61 ;
 RECT 14.56 1.71 14.66 2.425 ;
 RECT 10.675 0.475 10.775 0.88 ;
 RECT 15.095 1.91 16.015 2.01 ;
 RECT 10.675 0.375 14.11 0.475 ;
 RECT 10.585 0.88 10.815 1.09 ;
 RECT 16.225 0.455 18.155 0.535 ;
 RECT 17.925 0.535 18.155 0.6 ;
 RECT 17.925 0.39 18.155 0.435 ;
 RECT 16.305 0.435 18.155 0.455 ;
 RECT 16.225 0.535 16.455 0.665 ;
 RECT 17.08 0.535 17.31 0.835 ;
 RECT 17.08 0.835 17.18 2.39 ;
 RECT 26.11 0.215 26.21 0.995 ;
 RECT 26.11 0.995 26.35 1.205 ;
 RECT 26.11 1.205 26.21 2 ;
 RECT 28.505 0.375 28.605 0.99 ;
 RECT 28.505 0.99 28.755 1.2 ;
 RECT 28.505 1.2 28.605 2.27 ;
 RECT 28.505 2.27 28.79 2.48 ;
 RECT 13.49 0.655 13.59 2.305 ;
 RECT 13.795 2.3 14.025 2.305 ;
 RECT 13.795 2.405 14.025 2.51 ;
 RECT 13.49 2.305 14.025 2.405 ;
 RECT 25.33 0.21 25.43 0.755 ;
 RECT 25.33 0.855 25.43 2.2 ;
 RECT 28.195 1.125 28.295 2.2 ;
 RECT 24.365 0.755 25.9 0.84 ;
 RECT 24.365 0.84 25.895 0.855 ;
 RECT 25.8 0.215 25.9 0.755 ;
 RECT 24.365 0.595 24.595 0.755 ;
 RECT 25.33 2.2 28.295 2.3 ;
 RECT 12.2 1.28 12.48 1.45 ;
 RECT 12.2 1.45 12.3 1.655 ;
 RECT 12.2 0.655 12.3 1.18 ;
 RECT 12.2 1.655 13.16 1.755 ;
 RECT 13.06 1.755 13.16 2.355 ;
 RECT 11.285 0.66 11.385 1.18 ;
 RECT 12.2 1.755 12.3 2.51 ;
 RECT 11.285 1.24 12.48 1.28 ;
 RECT 11.285 1.18 12.3 1.24 ;
 RECT 27.02 0.38 27.12 0.96 ;
 RECT 27.02 1.06 27.12 1.14 ;
 RECT 26.6 0.935 26.83 0.96 ;
 RECT 26.6 0.96 27.12 1.06 ;
 RECT 26.6 1.06 26.83 1.145 ;
 RECT 27.02 1.14 27.29 1.24 ;
 RECT 27.19 1.24 27.29 1.84 ;
 RECT 27.385 0.22 27.615 0.28 ;
 RECT 27.385 0.38 27.615 0.43 ;
 RECT 27.02 0.28 27.615 0.38 ;
 RECT 11.275 1.575 11.375 2.485 ;
 RECT 11.785 1.575 12.015 1.685 ;
 RECT 11.275 1.475 12.015 1.575 ;
 RECT 29.205 0.195 29.305 2.665 ;
 RECT 28.195 0.095 29.305 0.195 ;
 RECT 24.57 1.245 24.67 2.665 ;
 RECT 28.195 0.195 28.295 0.945 ;
 RECT 24.57 1.2 24.855 1.245 ;
 RECT 24.625 1.035 24.855 1.1 ;
 RECT 24.57 2.665 29.305 2.765 ;
 RECT 24.57 1.1 24.9 1.2 ;
 RECT 15.5 0.795 15.665 0.925 ;
 RECT 14.82 0.885 15.05 0.925 ;
 RECT 14.82 1.025 15.05 1.095 ;
 RECT 14.82 0.925 15.665 1.025 ;
 RECT 15.5 0.585 15.73 0.795 ;
 RECT 2.535 1.55 2.775 1.78 ;
 RECT 2.675 1.78 2.775 2.695 ;
 RECT 1.065 1.435 1.635 1.71 ;
 RECT 1.065 0.515 1.165 1.435 ;
 RECT 1.065 1.71 1.165 2.645 ;
 RECT 1.535 0.515 1.635 1.435 ;
 RECT 1.535 1.71 1.635 2.695 ;
 RECT 2.255 1.37 2.355 1.605 ;
 RECT 2.485 0.515 2.585 1.14 ;
 RECT 2.205 1.705 2.305 2.695 ;
 RECT 2.205 1.605 2.355 1.705 ;
 RECT 2.255 1.14 2.585 1.37 ;
 RECT 1.87 0.515 1.97 1.105 ;
 RECT 1.83 1.105 2.075 1.345 ;
 RECT 4.42 0.52 4.52 2.465 ;
 RECT 4.18 0.27 4.52 0.52 ;
 RECT 7.05 1.33 7.19 1.475 ;
 RECT 7.05 1.71 7.15 2.475 ;
 RECT 7.09 0.65 7.19 1.33 ;
 RECT 7.05 1.475 7.28 1.71 ;
 RECT 6.6 0.705 6.7 1.165 ;
 RECT 6.16 1.27 6.26 1.445 ;
 RECT 6.6 0.47 6.885 0.705 ;
 RECT 6.16 1.17 6.7 1.265 ;
 RECT 6.16 1.265 6.535 1.27 ;
 RECT 6.39 1.165 6.7 1.17 ;
 RECT 6.015 1.445 6.26 1.69 ;
 RECT 7.49 0.715 7.59 1.61 ;
 RECT 7.525 1.71 7.625 2.48 ;
 RECT 7.49 1.61 7.625 1.71 ;
 RECT 7.37 0.485 7.61 0.715 ;
 RECT 13.095 0.655 13.195 1.24 ;
 RECT 12.965 1.24 13.195 1.475 ;
 RECT 4.895 0.49 4.995 1.495 ;
 RECT 4.7 1.495 4.995 1.745 ;
 RECT 4.895 1.745 4.995 2.37 ;
 RECT 2.975 0.135 3.075 0.22 ;
 RECT 2.815 0.22 3.075 0.43 ;
 RECT 2.975 0.43 3.075 2.695 ;
 RECT 3.445 0.295 3.545 1.115 ;
 RECT 3.28 1.115 3.545 1.325 ;
 RECT 3.445 1.325 3.545 2.74 ;
 RECT 19.52 0.77 19.62 2.155 ;
 RECT 19.52 0.55 19.62 0.56 ;
 RECT 19.52 0.56 19.775 0.77 ;
 RECT 20.885 0.39 20.985 1.4 ;
 RECT 20.155 0.43 20.255 1.245 ;
 RECT 21.375 0.51 21.475 1.4 ;
 RECT 21.375 1.5 21.475 2.26 ;
 RECT 20.885 1.5 20.985 2.235 ;
 RECT 20.09 0.22 20.32 0.29 ;
 RECT 20.09 0.39 20.32 0.43 ;
 RECT 20.09 0.29 20.985 0.39 ;
 RECT 20.885 1.4 21.475 1.5 ;
 RECT 20.105 1.245 20.335 1.455 ;
 RECT 8.31 2.445 8.57 2.655 ;
 RECT 8.47 1.79 8.57 2.445 ;
 RECT 18.58 1.445 18.68 2.035 ;
 RECT 18.565 2.035 18.795 2.245 ;
 RECT 19.05 0.55 19.15 2.69 ;
 RECT 9.98 1.58 10.08 1.615 ;
 RECT 9.72 1.01 9.82 1.48 ;
 RECT 9.98 1.825 10.08 2.69 ;
 RECT 9.98 1.615 10.215 1.825 ;
 RECT 9.72 1.48 10.08 1.58 ;
 RECT 9.98 2.69 19.15 2.79 ;
 RECT 9.42 1.01 9.52 1.615 ;
 RECT 9.28 1.615 9.52 1.825 ;
 RECT 9.42 1.825 9.52 2.51 ;
 RECT 22.98 0.375 23.08 1.33 ;
 RECT 22.4 1.25 22.65 1.33 ;
 RECT 22.4 1.33 23.08 1.43 ;
 RECT 22.4 1.43 22.65 1.46 ;
 RECT 22.4 0.385 22.5 1.25 ;
 RECT 22.4 1.46 22.5 2.69 ;
 RECT 22.98 1.43 23.08 2.695 ;
 RECT 23.585 0.22 23.815 0.275 ;
 RECT 23.585 0.375 23.815 0.43 ;
 RECT 22.98 0.275 23.815 0.375 ;
 RECT 17.55 0.73 17.65 1.39 ;
 RECT 17.415 1.39 17.65 1.6 ;
 RECT 17.55 1.6 17.65 2.39 ;
 RECT 5.67 1.62 5.77 2.675 ;
 RECT 5.735 0.185 14.625 0.19 ;
 RECT 14.525 0.19 14.625 1.29 ;
 RECT 5.735 0.19 7.89 0.285 ;
 RECT 5.735 0.285 5.835 1.52 ;
 RECT 15.42 1.39 15.615 1.405 ;
 RECT 6.555 1.565 6.655 2.675 ;
 RECT 5.235 1.44 5.48 1.52 ;
 RECT 5.235 1.62 5.48 1.69 ;
 RECT 5.235 1.52 5.835 1.62 ;
 RECT 7.79 0.285 7.89 1.24 ;
 RECT 7.79 0.09 14.625 0.185 ;
 RECT 14.525 1.29 15.615 1.39 ;
 RECT 5.67 2.675 6.655 2.775 ;
 RECT 15.42 1.405 15.65 1.615 ;
 LAYER CO ;
 RECT 2.865 0.26 2.995 0.39 ;
 RECT 3.33 1.155 3.46 1.285 ;
 RECT 22.47 1.29 22.6 1.42 ;
 RECT 20.155 1.285 20.285 1.415 ;
 RECT 17.975 0.43 18.105 0.56 ;
 RECT 19.595 0.6 19.725 0.73 ;
 RECT 20.14 0.26 20.27 0.39 ;
 RECT 8.36 2.485 8.49 2.615 ;
 RECT 18.615 2.075 18.745 2.205 ;
 RECT 10.035 1.655 10.165 1.785 ;
 RECT 9.33 1.655 9.46 1.785 ;
 RECT 23.635 0.26 23.765 0.39 ;
 RECT 28.575 1.03 28.705 1.16 ;
 RECT 16.275 0.495 16.405 0.625 ;
 RECT 17.465 1.43 17.595 1.56 ;
 RECT 15.55 0.625 15.68 0.755 ;
 RECT 15.47 1.445 15.6 1.575 ;
 RECT 25.725 1.075 25.855 1.205 ;
 RECT 10.635 0.92 10.765 1.05 ;
 RECT 26.65 0.975 26.78 1.105 ;
 RECT 17.13 0.665 17.26 0.795 ;
 RECT 26.17 1.035 26.3 1.165 ;
 RECT 28.61 2.31 28.74 2.44 ;
 RECT 13.845 2.34 13.975 2.47 ;
 RECT 24.415 0.635 24.545 0.765 ;
 RECT 12.3 1.28 12.43 1.41 ;
 RECT 27.435 0.26 27.565 0.39 ;
 RECT 11.835 1.515 11.965 1.645 ;
 RECT 24.675 1.075 24.805 1.205 ;
 RECT 14.87 0.925 15 1.055 ;
 RECT 4.76 1.55 4.89 1.68 ;
 RECT 1.285 0.735 1.415 0.865 ;
 RECT 1.29 1.51 1.42 1.64 ;
 RECT 0.815 0.735 0.945 0.865 ;
 RECT 3.195 2.31 3.325 2.44 ;
 RECT 1.285 2.015 1.415 2.145 ;
 RECT 1.89 1.155 2.02 1.285 ;
 RECT 3.195 2.05 3.325 2.18 ;
 RECT 2.59 1.6 2.72 1.73 ;
 RECT 3.665 2.01 3.795 2.14 ;
 RECT 3.665 0.735 3.795 0.865 ;
 RECT 2.425 2.075 2.555 2.205 ;
 RECT 1.285 2.275 1.415 2.405 ;
 RECT 3.195 0.545 3.325 0.675 ;
 RECT 3.665 1.75 3.795 1.88 ;
 RECT 0.815 2.015 0.945 2.145 ;
 RECT 2.23 0.735 2.36 0.865 ;
 RECT 2.41 1.19 2.54 1.32 ;
 RECT 12.65 2.225 12.78 2.355 ;
 RECT 21.63 0.975 21.76 1.105 ;
 RECT 22.62 2.64 22.75 2.77 ;
 RECT 4.17 2.115 4.3 2.245 ;
 RECT 21.115 0.36 21.245 0.49 ;
 RECT 23.205 0.63 23.335 0.76 ;
 RECT 27.27 0.595 27.4 0.725 ;
 RECT 6.705 0.525 6.835 0.655 ;
 RECT 7.75 1.825 7.88 1.955 ;
 RECT 27.78 1.49 27.91 1.62 ;
 RECT 6.35 0.88 6.48 1.01 ;
 RECT 14.78 1.87 14.91 2 ;
 RECT 8.22 2.11 8.35 2.24 ;
 RECT 8.035 0.31 8.165 0.44 ;
 RECT 25.55 0.135 25.68 0.265 ;
 RECT 5.295 1.495 5.425 1.625 ;
 RECT 5.245 0.745 5.375 0.875 ;
 RECT 5.115 1.995 5.245 2.125 ;
 RECT 11.95 1.995 12.08 2.125 ;
 RECT 0.315 0.59 0.445 0.72 ;
 RECT 11.505 2.07 11.635 2.2 ;
 RECT 14.275 0.595 14.405 0.725 ;
 RECT 6.07 1.49 6.2 1.62 ;
 RECT 13.015 1.28 13.145 1.41 ;
 RECT 22.145 1.725 22.275 1.855 ;
 RECT 0.315 2.085 0.445 2.215 ;
 RECT 9.71 2.045 9.84 2.175 ;
 RECT 5.225 0.145 5.355 0.275 ;
 RECT 14.275 1.9 14.405 2.03 ;
 RECT 0.315 2.345 0.445 2.475 ;
 RECT 5.38 2.345 5.51 2.475 ;
 RECT 26.33 0.435 26.46 0.565 ;
 RECT 20.625 1.705 20.755 1.835 ;
 RECT 9.94 1.23 10.07 1.36 ;
 RECT 18.8 1.705 18.93 1.835 ;
 RECT 9.17 2.075 9.3 2.205 ;
 RECT 6.82 0.88 6.95 1.01 ;
 RECT 16.83 1.835 16.96 1.965 ;
 RECT 16.7 0.765 16.83 0.895 ;
 RECT 4.64 0.74 4.77 0.87 ;
 RECT 27.945 0.12 28.075 0.25 ;
 RECT 7.425 0.53 7.555 0.66 ;
 RECT 22.145 0.62 22.275 0.75 ;
 RECT 15.675 2.38 15.805 2.51 ;
 RECT 11.95 0.895 12.08 1.025 ;
 RECT 25.08 1.425 25.21 1.555 ;
 RECT 0.315 0.33 0.445 0.46 ;
 RECT 19.865 0.92 19.995 1.05 ;
 RECT 25.55 1.475 25.68 1.605 ;
 RECT 13.75 0.875 13.88 1.005 ;
 RECT 5.955 0.79 6.085 0.92 ;
 RECT 17.77 1.835 17.9 1.965 ;
 RECT 6.8 2.07 6.93 2.2 ;
 RECT 29.505 1.475 29.635 1.605 ;
 RECT 21.63 1.705 21.76 1.835 ;
 RECT 23.205 1.71 23.335 1.84 ;
 RECT 20.625 0.975 20.755 1.105 ;
 RECT 4.17 0.74 4.3 0.87 ;
 RECT 5.89 1.825 6.02 1.955 ;
 RECT 13.75 1.945 13.88 2.075 ;
 RECT 4.64 2.05 4.77 2.18 ;
 RECT 24.83 0.505 24.96 0.635 ;
 RECT 11.025 2.015 11.155 2.145 ;
 RECT 26.765 0.12 26.895 0.25 ;
 RECT 26.33 1.485 26.46 1.615 ;
 RECT 28.725 1.465 28.855 1.595 ;
 RECT 19.27 1.705 19.4 1.835 ;
 RECT 28.725 0.595 28.855 0.725 ;
 RECT 7.1 1.525 7.23 1.655 ;
 RECT 19.745 1.705 19.875 1.835 ;
 RECT 21.03 2.64 21.16 2.77 ;
 RECT 27.41 1.405 27.54 1.535 ;
 RECT 11.03 0.905 11.16 1.035 ;
 RECT 4.24 0.325 4.37 0.455 ;
 RECT 9.17 0.31 9.3 0.44 ;
 RECT 11.505 0.905 11.635 1.035 ;
 RECT 14.78 0.595 14.91 0.725 ;
 RECT 12.84 0.6 12.97 0.73 ;
 RECT 26.935 1.445 27.065 1.575 ;
 RECT 0.315 1.825 0.445 1.955 ;
 RECT 17.805 1.035 17.935 1.165 ;
 RECT 18.39 0.91 18.52 1.04 ;
 RECT 10.2 2.42 10.33 2.55 ;
 RECT 22.705 0.62 22.835 0.75 ;
 RECT 8.69 2.135 8.82 2.265 ;
 RECT 6.305 2.105 6.435 2.235 ;
 RECT 7.27 2.11 7.4 2.24 ;
 LAYER M1 ;
 RECT 6.815 0.805 6.955 1.22 ;
 RECT 6.64 1.22 6.955 1.36 ;
 RECT 6.64 1.36 6.78 1.82 ;
 RECT 9.28 1.615 9.51 1.65 ;
 RECT 9.28 1.79 9.51 1.825 ;
 RECT 8.08 1.65 9.515 1.79 ;
 RECT 27.265 0.73 27.405 1.04 ;
 RECT 27.405 1.18 27.545 1.605 ;
 RECT 27.2 0.59 27.475 0.73 ;
 RECT 28.525 0.99 28.755 1.04 ;
 RECT 27.265 1.04 28.755 1.18 ;
 RECT 28.525 1.18 28.755 1.2 ;
 RECT 27.385 0.29 27.755 0.43 ;
 RECT 27.615 0.43 27.755 0.71 ;
 RECT 27.385 0.22 27.615 0.29 ;
 RECT 29.035 0.85 29.175 1.385 ;
 RECT 28.72 1.525 28.86 1.73 ;
 RECT 27.615 0.71 29.175 0.85 ;
 RECT 28.72 0.51 28.86 0.71 ;
 RECT 28.72 1.385 29.175 1.525 ;
 RECT 26.645 1.145 26.785 1.345 ;
 RECT 26.325 1.485 26.465 1.76 ;
 RECT 26.645 0.73 26.785 0.935 ;
 RECT 26.325 0.355 26.465 0.59 ;
 RECT 26.325 1.345 26.785 1.485 ;
 RECT 26.6 0.935 26.83 1.145 ;
 RECT 26.325 0.59 26.785 0.73 ;
 RECT 24.625 1.225 24.855 1.245 ;
 RECT 24.625 1.195 25.215 1.225 ;
 RECT 24.765 1.015 25.075 1.035 ;
 RECT 24.625 1.035 25.075 1.055 ;
 RECT 24.9 0.64 25.04 1.015 ;
 RECT 25.075 1.225 25.215 1.75 ;
 RECT 24.78 0.5 25.04 0.64 ;
 RECT 25.675 1.035 25.905 1.055 ;
 RECT 25.675 1.195 25.905 1.245 ;
 RECT 24.625 1.055 25.905 1.195 ;
 RECT 23.585 0.36 23.815 0.43 ;
 RECT 25.18 0.36 25.32 0.565 ;
 RECT 23.585 0.22 25.32 0.36 ;
 RECT 25.92 0.705 26.06 0.75 ;
 RECT 26.045 0.995 26.35 1.205 ;
 RECT 26.045 0.89 26.185 0.995 ;
 RECT 25.92 0.75 26.185 0.89 ;
 RECT 25.18 0.565 26.06 0.705 ;
 RECT 18.82 0.775 18.96 1.405 ;
 RECT 19.545 0.56 19.775 0.635 ;
 RECT 17.8 1.405 18.96 1.545 ;
 RECT 17.8 1.545 17.94 1.83 ;
 RECT 17.8 1.17 17.94 1.405 ;
 RECT 16.755 1.83 18.005 1.97 ;
 RECT 17.73 1.03 18.01 1.17 ;
 RECT 21.74 0.36 21.88 0.635 ;
 RECT 18.82 0.635 21.88 0.775 ;
 RECT 22.42 0.36 22.56 1.25 ;
 RECT 22.42 1.25 22.65 1.46 ;
 RECT 21.74 0.22 22.56 0.36 ;
 RECT 17.925 0.28 20.32 0.42 ;
 RECT 17.925 0.42 18.155 0.6 ;
 RECT 20.09 0.22 20.32 0.28 ;
 RECT 20.09 0.42 20.32 0.43 ;
 RECT 11.5 1.04 11.64 2.34 ;
 RECT 11.43 0.9 11.685 1.04 ;
 RECT 12.295 2.055 12.435 2.34 ;
 RECT 11.5 2.34 12.435 2.48 ;
 RECT 13.745 0.765 13.885 1.915 ;
 RECT 13.745 2.055 13.885 2.145 ;
 RECT 12.295 1.915 14.41 2.055 ;
 RECT 14.27 0.525 14.41 1.915 ;
 RECT 14.27 2.055 14.41 2.11 ;
 RECT 14.775 0.525 14.915 0.885 ;
 RECT 14.775 1.095 14.915 2.065 ;
 RECT 14.775 0.885 15.05 1.095 ;
 RECT 17.08 0.57 17.31 0.95 ;
 RECT 15.5 0.585 16.455 0.63 ;
 RECT 16.225 0.63 16.455 0.665 ;
 RECT 16.225 0.455 16.455 0.49 ;
 RECT 15.525 0.49 16.455 0.585 ;
 RECT 15.5 0.63 15.73 0.795 ;
 RECT 5.95 1.67 6.09 1.82 ;
 RECT 5.95 1.96 6.09 2.51 ;
 RECT 5.95 0.5 6.09 1.44 ;
 RECT 5.95 1.44 6.205 1.67 ;
 RECT 5.82 1.82 6.09 1.96 ;
 RECT 8.31 2.445 8.54 2.51 ;
 RECT 8.31 2.65 8.54 2.655 ;
 RECT 5.95 2.51 8.54 2.65 ;
 RECT 7.095 0.66 7.235 0.895 ;
 RECT 6.635 0.52 7.235 0.66 ;
 RECT 7.095 0.895 10.815 1.035 ;
 RECT 10.585 0.88 10.815 0.895 ;
 RECT 10.585 1.035 10.815 1.09 ;
 RECT 5.195 0.88 5.335 1.475 ;
 RECT 5.155 1.63 5.295 1.99 ;
 RECT 5.155 1.475 5.5 1.63 ;
 RECT 5.045 1.99 5.295 2.13 ;
 RECT 5.195 0.74 5.515 0.88 ;
 RECT 2.88 0.87 3.02 1.15 ;
 RECT 2.88 1.29 3.02 2.07 ;
 RECT 2.37 2.07 3.02 2.21 ;
 RECT 2.175 0.73 3.02 0.87 ;
 RECT 3.28 1.115 3.51 1.15 ;
 RECT 3.28 1.29 3.51 1.325 ;
 RECT 2.88 1.15 3.51 1.29 ;
 RECT 3.945 0.875 4.085 1.195 ;
 RECT 3.945 1.335 4.085 2.11 ;
 RECT 3.945 2.25 4.085 2.255 ;
 RECT 3.945 2.11 4.37 2.25 ;
 RECT 3.945 0.735 4.37 0.875 ;
 RECT 4.915 0.6 5.055 1.195 ;
 RECT 3.945 1.195 5.055 1.335 ;
 RECT 6.345 0.36 6.485 2.035 ;
 RECT 5.66 0.22 6.485 0.36 ;
 RECT 5.66 0.36 5.8 0.46 ;
 RECT 6.3 2.17 6.44 2.305 ;
 RECT 6.3 2.035 6.485 2.17 ;
 RECT 4.915 0.46 5.8 0.6 ;
 RECT 3.66 0.46 3.8 2.21 ;
 RECT 4.13 0.22 4.495 0.32 ;
 RECT 4.13 0.46 4.495 0.525 ;
 RECT 3.66 0.32 4.495 0.46 ;
 RECT 0.81 0.68 0.95 1.155 ;
 RECT 0.81 1.295 0.95 2.23 ;
 RECT 1.595 0.36 1.735 1.155 ;
 RECT 0.81 1.155 1.735 1.295 ;
 RECT 2.815 0.36 3.045 0.43 ;
 RECT 1.595 0.22 3.045 0.36 ;
 RECT 19.63 1.7 19.925 1.84 ;
 RECT 19.63 1.84 19.77 2.075 ;
 RECT 18.935 1.84 19.075 2.075 ;
 RECT 18.74 1.7 19.075 1.84 ;
 RECT 18.935 2.075 19.77 2.215 ;
 RECT 19.825 1.055 19.965 1.245 ;
 RECT 19.265 1.385 19.405 1.625 ;
 RECT 20.105 1.385 20.335 1.455 ;
 RECT 19.265 1.245 20.335 1.385 ;
 RECT 19.795 0.915 20.095 1.055 ;
 RECT 19.235 1.625 19.49 1.92 ;
 RECT 20.335 2.205 20.475 2.39 ;
 RECT 16.19 1.895 16.33 2.39 ;
 RECT 16.19 2.39 20.475 2.53 ;
 RECT 15.065 1.755 16.33 1.895 ;
 RECT 15.065 1.895 15.205 2.34 ;
 RECT 13.795 2.3 14.025 2.34 ;
 RECT 13.795 2.48 14.025 2.51 ;
 RECT 13.795 2.34 15.205 2.48 ;
 RECT 20.335 2.065 24.36 2.205 ;
 RECT 24.22 2.205 24.36 2.52 ;
 RECT 28.56 2.48 28.7 2.52 ;
 RECT 24.22 2.52 28.7 2.66 ;
 RECT 28.56 2.27 28.79 2.48 ;
 RECT 16.47 1.56 16.61 2.11 ;
 RECT 15.42 1.405 15.65 1.42 ;
 RECT 15.42 1.56 15.65 1.615 ;
 RECT 15.42 1.42 16.61 1.56 ;
 RECT 16.47 2.11 18.795 2.245 ;
 RECT 16.47 2.245 18.79 2.25 ;
 RECT 18.565 2.035 18.795 2.11 ;
 RECT 11.785 1.475 12.085 1.635 ;
 RECT 11.945 1.775 12.085 2.18 ;
 RECT 11.945 0.825 12.085 1.475 ;
 RECT 11.785 1.635 13.145 1.685 ;
 RECT 13.005 1.415 13.145 1.635 ;
 RECT 11.945 1.685 13.145 1.775 ;
 RECT 12.96 1.275 13.215 1.415 ;
 RECT 7.2 2.105 8.42 2.245 ;
 RECT 7.76 1.365 7.9 1.5 ;
 RECT 6.93 1.64 7.435 1.675 ;
 RECT 6.93 1.5 7.9 1.64 ;
 RECT 9.705 1.365 9.845 2.25 ;
 RECT 11.02 1.04 11.16 1.23 ;
 RECT 11.02 1.37 11.16 2.215 ;
 RECT 11.02 0.885 11.16 0.9 ;
 RECT 7.76 1.23 11.16 1.365 ;
 RECT 7.76 1.225 10.41 1.23 ;
 RECT 10.15 1.365 11.16 1.37 ;
 RECT 10.955 0.9 11.23 1.04 ;
 RECT 6.64 1.82 8.22 1.96 ;
 RECT 8.08 1.79 8.22 1.82 ;
 RECT 6.725 1.96 7.005 2.215 ;
 END
END RSDFFNSRASRX1

MACRO RSDFFNSRASRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 32.64 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 25.92 0.59 26.29 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 31.15 1.435 31.49 1.8 ;
 RECT 29.47 1.99 31.335 2.13 ;
 RECT 27.24 2.22 29.61 2.36 ;
 RECT 29.47 1.435 29.61 1.99 ;
 RECT 31.195 1.8 31.335 1.99 ;
 RECT 27.24 1.39 27.38 2.22 ;
 RECT 28.625 1.37 28.765 2.22 ;
 RECT 29.47 2.13 29.61 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 5.145 0.08 5.425 0.295 ;
 RECT 29.59 0.08 29.83 0.26 ;
 RECT 9.075 0.31 9.365 0.45 ;
 RECT 12.755 0.595 13.035 0.735 ;
 RECT 16.685 0.275 17.71 0.415 ;
 RECT 21.22 0.29 21.485 0.45 ;
 RECT 17.57 0.75 18.515 0.89 ;
 RECT 0 -0.08 32.64 0.08 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.625 0.08 4.765 0.97 ;
 RECT 3.18 0.08 3.32 0.74 ;
 RECT 1.27 0.08 1.41 0.93 ;
 RECT 7.97 0.08 8.205 0.46 ;
 RECT 16.685 0.415 16.825 0.945 ;
 RECT 22.855 0.08 22.995 0.92 ;
 RECT 27.24 0.08 27.38 0.36 ;
 RECT 28.455 0.08 28.595 0.35 ;
 RECT 18.375 0.89 18.515 1.11 ;
 RECT 17.57 0.415 17.71 0.75 ;
 RECT 9.155 0.08 9.295 0.31 ;
 RECT 12.825 0.08 12.965 0.595 ;
 RECT 16.685 0.08 16.825 0.275 ;
 RECT 21.275 0.08 21.415 0.29 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 32.64 2.96 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.27 1.965 1.41 2.8 ;
 RECT 3.18 1.99 3.32 2.8 ;
 RECT 4.625 1.98 4.765 2.8 ;
 RECT 5.3 2.34 5.55 2.8 ;
 RECT 8.675 2.07 8.815 2.8 ;
 RECT 9.155 1.98 9.295 2.8 ;
 RECT 12.635 2.37 12.775 2.8 ;
 RECT 10.185 2.365 10.325 2.8 ;
 RECT 15.595 2.335 15.865 2.8 ;
 RECT 21.265 2.54 21.405 2.8 ;
 RECT 22.77 2.57 22.91 2.8 ;
 RECT 23.825 2.57 23.965 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.675 1.475 5.005 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.215 1.16 12.67 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.365 0.485 7.68 0.605 ;
 RECT 11.42 0.545 12.615 0.605 ;
 RECT 7.365 0.605 12.615 0.685 ;
 RECT 12.475 0.685 12.615 0.875 ;
 RECT 12.475 0.875 13.34 1.015 ;
 RECT 13.2 0.245 15.345 0.255 ;
 RECT 13.2 0.255 15.35 0.385 ;
 RECT 15.21 1.09 17.2 1.23 ;
 RECT 17.405 1.56 17.635 1.6 ;
 RECT 17.06 1.42 17.635 1.56 ;
 RECT 17.405 1.39 17.635 1.42 ;
 RECT 7.365 0.685 11.56 0.745 ;
 RECT 13.2 0.385 13.34 0.875 ;
 RECT 15.21 0.385 15.35 1.09 ;
 RECT 17.06 1.23 17.2 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.975 1.61 10.415 2.04 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.435 1.615 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.78 1.59 2.725 1.75 ;
 RECT 1.875 1.09 2.015 1.44 ;
 RECT 1.78 1.44 2.025 1.59 ;
 RECT 2.575 1.75 2.715 1.805 ;
 RECT 2.575 1.53 2.715 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.24 1.115 2.66 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.58 1.27 20.925 1.545 ;
 RECT 20.715 0.93 21.04 1.07 ;
 RECT 21.7 0.93 22.025 1.07 ;
 RECT 20.785 1.71 21.93 1.85 ;
 RECT 20.785 1.85 20.925 1.895 ;
 RECT 20.785 1.545 20.925 1.71 ;
 RECT 20.785 1.07 20.925 1.27 ;
 RECT 20.785 0.915 20.925 0.93 ;
 RECT 21.79 0.925 21.93 0.93 ;
 RECT 21.79 1.85 21.93 1.895 ;
 RECT 21.79 1.07 21.93 1.71 ;
 END
 ANTENNADIFFAREA 0.805 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.195 1.285 22.435 1.525 ;
 RECT 22.295 1.775 24.5 1.915 ;
 RECT 22.295 0.645 22.435 1.285 ;
 RECT 23.355 1.915 23.495 1.92 ;
 RECT 23.355 0.66 23.495 1.775 ;
 RECT 22.295 1.915 22.435 1.925 ;
 RECT 22.295 1.525 22.435 1.775 ;
 END
 ANTENNADIFFAREA 1.186 ;
 END Q

 OBS
 LAYER PO ;
 RECT 27.37 1.035 27.6 1.245 ;
 RECT 15.905 0.105 18.73 0.205 ;
 RECT 15.905 0.205 16.005 1.91 ;
 RECT 18.63 0.205 18.73 1.265 ;
 RECT 15.085 1.71 15.185 1.91 ;
 RECT 14 1.61 15.185 1.71 ;
 RECT 14 0.475 14.1 1.61 ;
 RECT 14.55 1.71 14.65 2.425 ;
 RECT 10.665 0.475 10.765 0.895 ;
 RECT 15.085 1.91 16.005 2.01 ;
 RECT 10.665 0.375 14.1 0.475 ;
 RECT 10.54 0.895 10.77 1.105 ;
 RECT 16.215 0.455 18.145 0.535 ;
 RECT 17.915 0.535 18.145 0.6 ;
 RECT 17.915 0.39 18.145 0.435 ;
 RECT 16.295 0.435 18.145 0.455 ;
 RECT 16.215 0.535 16.445 0.665 ;
 RECT 17.07 0.535 17.3 0.835 ;
 RECT 17.07 0.835 17.17 2.39 ;
 RECT 27.805 0.215 27.905 0.995 ;
 RECT 27.805 0.995 28.045 1.205 ;
 RECT 27.805 1.205 27.905 2 ;
 RECT 30.2 0.375 30.3 0.99 ;
 RECT 30.2 0.99 30.45 1.2 ;
 RECT 30.2 1.2 30.3 2.27 ;
 RECT 30.2 2.27 30.485 2.48 ;
 RECT 13.48 0.655 13.58 2.305 ;
 RECT 13.785 2.3 14.015 2.305 ;
 RECT 13.785 2.405 14.015 2.51 ;
 RECT 13.48 2.305 14.015 2.405 ;
 RECT 27.025 0.21 27.125 0.755 ;
 RECT 27.025 0.855 27.125 2.2 ;
 RECT 29.89 1.125 29.99 2.2 ;
 RECT 26.06 0.755 27.595 0.84 ;
 RECT 26.06 0.84 27.59 0.855 ;
 RECT 27.495 0.215 27.595 0.755 ;
 RECT 26.06 0.595 26.29 0.755 ;
 RECT 27.025 2.2 29.99 2.3 ;
 RECT 12.19 1.28 12.445 1.47 ;
 RECT 12.19 1.47 12.29 1.655 ;
 RECT 12.19 0.655 12.29 1.18 ;
 RECT 12.19 1.655 13.15 1.755 ;
 RECT 13.05 1.755 13.15 2.355 ;
 RECT 11.275 0.66 11.375 1.18 ;
 RECT 12.19 1.755 12.29 2.51 ;
 RECT 11.275 1.26 12.445 1.28 ;
 RECT 11.275 1.18 12.29 1.26 ;
 RECT 28.715 0.38 28.815 0.96 ;
 RECT 28.715 1.06 28.815 1.14 ;
 RECT 28.295 0.935 28.525 0.96 ;
 RECT 28.295 0.96 28.815 1.06 ;
 RECT 28.295 1.06 28.525 1.145 ;
 RECT 28.715 1.14 28.985 1.24 ;
 RECT 28.885 1.24 28.985 1.84 ;
 RECT 29.08 0.22 29.31 0.28 ;
 RECT 29.08 0.38 29.31 0.43 ;
 RECT 28.715 0.28 29.31 0.38 ;
 RECT 11.265 1.575 11.365 2.485 ;
 RECT 11.775 1.575 12.005 1.685 ;
 RECT 11.265 1.475 12.005 1.575 ;
 RECT 30.9 0.195 31 2.665 ;
 RECT 29.89 0.095 31 0.195 ;
 RECT 26.265 1.245 26.365 2.665 ;
 RECT 29.89 0.195 29.99 0.945 ;
 RECT 26.265 1.2 26.55 1.245 ;
 RECT 26.32 1.035 26.55 1.1 ;
 RECT 26.265 2.665 31 2.765 ;
 RECT 26.265 1.1 26.595 1.2 ;
 RECT 15.49 0.795 15.655 0.925 ;
 RECT 14.81 0.885 15.04 0.925 ;
 RECT 14.81 1.025 15.04 1.095 ;
 RECT 14.81 0.925 15.655 1.025 ;
 RECT 15.49 0.585 15.72 0.795 ;
 RECT 2.525 1.55 2.765 1.78 ;
 RECT 2.665 1.78 2.765 2.695 ;
 RECT 1.055 1.435 1.625 1.71 ;
 RECT 1.055 0.515 1.155 1.435 ;
 RECT 1.055 1.71 1.155 2.645 ;
 RECT 1.525 0.515 1.625 1.435 ;
 RECT 1.525 1.71 1.625 2.695 ;
 RECT 2.245 1.37 2.345 1.605 ;
 RECT 2.475 0.515 2.575 1.14 ;
 RECT 2.195 1.705 2.295 2.695 ;
 RECT 2.195 1.605 2.345 1.705 ;
 RECT 2.245 1.14 2.575 1.37 ;
 RECT 1.86 0.515 1.96 1.105 ;
 RECT 1.82 1.105 2.065 1.345 ;
 RECT 4.41 0.52 4.51 2.465 ;
 RECT 4.17 0.27 4.51 0.52 ;
 RECT 7.04 1.33 7.18 1.475 ;
 RECT 7.04 1.71 7.14 2.475 ;
 RECT 7.08 0.65 7.18 1.33 ;
 RECT 7.04 1.475 7.27 1.71 ;
 RECT 6.59 0.705 6.69 1.165 ;
 RECT 6.15 1.27 6.25 1.445 ;
 RECT 6.59 0.47 6.875 0.705 ;
 RECT 6.15 1.17 6.69 1.265 ;
 RECT 6.15 1.265 6.525 1.27 ;
 RECT 6.38 1.165 6.69 1.17 ;
 RECT 6.005 1.445 6.25 1.69 ;
 RECT 7.48 0.715 7.58 1.61 ;
 RECT 7.515 1.71 7.615 2.48 ;
 RECT 7.48 1.61 7.615 1.71 ;
 RECT 7.36 0.485 7.6 0.715 ;
 RECT 13.085 0.655 13.185 1.24 ;
 RECT 12.955 1.24 13.185 1.475 ;
 RECT 4.885 0.49 4.985 1.495 ;
 RECT 4.69 1.495 4.985 1.745 ;
 RECT 4.885 1.745 4.985 2.37 ;
 RECT 2.8 0.245 3.065 0.455 ;
 RECT 2.965 0.455 3.065 2.695 ;
 RECT 3.435 0.295 3.535 1.115 ;
 RECT 3.245 1.115 3.535 1.325 ;
 RECT 3.435 1.325 3.535 2.765 ;
 RECT 19.51 0.77 19.61 2.155 ;
 RECT 19.51 0.55 19.61 0.56 ;
 RECT 19.51 0.56 19.765 0.77 ;
 RECT 21.05 0.375 21.15 1.41 ;
 RECT 20.145 0.215 20.245 0.22 ;
 RECT 20.145 0.43 20.245 1.245 ;
 RECT 21.54 0.445 21.64 1.41 ;
 RECT 21.54 1.51 21.64 2.645 ;
 RECT 21.05 1.51 21.15 2.57 ;
 RECT 20.145 0.22 20.375 0.275 ;
 RECT 20.145 0.375 20.375 0.43 ;
 RECT 20.145 0.275 21.15 0.375 ;
 RECT 21.05 1.41 21.64 1.51 ;
 RECT 20.095 1.245 20.325 1.455 ;
 RECT 8.3 2.445 8.56 2.655 ;
 RECT 8.46 1.79 8.56 2.445 ;
 RECT 18.57 1.445 18.67 2.035 ;
 RECT 18.555 2.035 18.785 2.245 ;
 RECT 19.04 0.55 19.14 2.69 ;
 RECT 9.97 1.58 10.07 1.615 ;
 RECT 9.71 1.01 9.81 1.48 ;
 RECT 9.97 1.825 10.07 2.69 ;
 RECT 9.97 1.615 10.205 1.825 ;
 RECT 9.71 1.48 10.07 1.58 ;
 RECT 9.97 2.69 19.14 2.79 ;
 RECT 9.41 0.98 9.51 1.615 ;
 RECT 9.27 1.615 9.51 1.825 ;
 RECT 9.41 1.825 9.51 2.51 ;
 RECT 23.135 0.375 23.235 1.295 ;
 RECT 22.555 1.295 24.18 1.395 ;
 RECT 22.555 1.26 22.805 1.295 ;
 RECT 22.555 0.375 22.655 1.26 ;
 RECT 24.08 1.395 24.18 2.685 ;
 RECT 23.61 1.395 23.71 2.69 ;
 RECT 22.555 1.47 22.655 2.69 ;
 RECT 22.555 1.395 22.805 1.47 ;
 RECT 23.135 1.395 23.235 2.715 ;
 RECT 25.28 0.22 25.51 0.275 ;
 RECT 25.28 0.375 25.51 0.43 ;
 RECT 23.135 0.275 25.51 0.375 ;
 RECT 17.54 0.73 17.64 1.39 ;
 RECT 17.405 1.39 17.64 1.6 ;
 RECT 17.54 1.6 17.64 2.39 ;
 RECT 5.725 0.285 5.825 1.52 ;
 RECT 5.225 1.52 5.825 1.62 ;
 RECT 5.725 0.185 14.615 0.195 ;
 RECT 7.78 0.095 14.615 0.185 ;
 RECT 5.725 0.195 7.88 0.285 ;
 RECT 14.515 0.195 14.615 1.29 ;
 RECT 15.41 1.39 15.605 1.405 ;
 RECT 6.545 1.565 6.645 2.675 ;
 RECT 5.66 1.62 5.76 2.675 ;
 RECT 5.225 1.44 5.47 1.52 ;
 RECT 5.225 1.62 5.47 1.69 ;
 RECT 7.78 0.285 7.88 1.24 ;
 RECT 14.515 1.29 15.605 1.39 ;
 RECT 5.66 2.675 6.645 2.775 ;
 RECT 15.41 1.405 15.64 1.615 ;
 RECT 27.5 1.245 27.6 2.02 ;
 LAYER CO ;
 RECT 20.145 1.285 20.275 1.415 ;
 RECT 17.965 0.43 18.095 0.56 ;
 RECT 19.585 0.6 19.715 0.73 ;
 RECT 20.195 0.26 20.325 0.39 ;
 RECT 8.35 2.485 8.48 2.615 ;
 RECT 18.605 2.075 18.735 2.205 ;
 RECT 10.025 1.655 10.155 1.785 ;
 RECT 9.32 1.655 9.45 1.785 ;
 RECT 25.33 0.26 25.46 0.39 ;
 RECT 30.27 1.03 30.4 1.16 ;
 RECT 16.265 0.495 16.395 0.625 ;
 RECT 17.455 1.43 17.585 1.56 ;
 RECT 15.54 0.625 15.67 0.755 ;
 RECT 15.46 1.445 15.59 1.575 ;
 RECT 27.42 1.075 27.55 1.205 ;
 RECT 10.59 0.935 10.72 1.065 ;
 RECT 28.345 0.975 28.475 1.105 ;
 RECT 17.12 0.665 17.25 0.795 ;
 RECT 27.865 1.035 27.995 1.165 ;
 RECT 30.305 2.31 30.435 2.44 ;
 RECT 13.835 2.34 13.965 2.47 ;
 RECT 26.11 0.635 26.24 0.765 ;
 RECT 12.265 1.3 12.395 1.43 ;
 RECT 29.13 0.26 29.26 0.39 ;
 RECT 11.825 1.515 11.955 1.645 ;
 RECT 26.37 1.075 26.5 1.205 ;
 RECT 14.86 0.925 14.99 1.055 ;
 RECT 4.75 1.55 4.88 1.68 ;
 RECT 20.79 1.715 20.92 1.845 ;
 RECT 22.86 0.72 22.99 0.85 ;
 RECT 21.795 0.935 21.925 1.065 ;
 RECT 1.275 0.735 1.405 0.865 ;
 RECT 1.28 1.51 1.41 1.64 ;
 RECT 0.805 0.735 0.935 0.865 ;
 RECT 3.185 2.31 3.315 2.44 ;
 RECT 1.275 2.015 1.405 2.145 ;
 RECT 1.88 1.155 2.01 1.285 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 2.58 1.6 2.71 1.73 ;
 RECT 3.655 2.01 3.785 2.14 ;
 RECT 3.655 0.735 3.785 0.865 ;
 RECT 2.415 2.075 2.545 2.205 ;
 RECT 1.275 2.275 1.405 2.405 ;
 RECT 3.185 0.545 3.315 0.675 ;
 RECT 3.655 1.75 3.785 1.88 ;
 RECT 0.805 2.015 0.935 2.145 ;
 RECT 2.22 0.735 2.35 0.865 ;
 RECT 2.4 1.19 2.53 1.32 ;
 RECT 28.965 0.595 29.095 0.725 ;
 RECT 6.695 0.525 6.825 0.655 ;
 RECT 7.74 1.825 7.87 1.955 ;
 RECT 29.475 1.49 29.605 1.62 ;
 RECT 6.34 0.88 6.47 1.01 ;
 RECT 14.77 1.87 14.9 2 ;
 RECT 8.21 2.11 8.34 2.24 ;
 RECT 8.025 0.32 8.155 0.45 ;
 RECT 27.245 0.135 27.375 0.265 ;
 RECT 5.285 1.495 5.415 1.625 ;
 RECT 5.235 0.745 5.365 0.875 ;
 RECT 5.105 1.995 5.235 2.125 ;
 RECT 11.94 1.995 12.07 2.125 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 11.495 2.07 11.625 2.2 ;
 RECT 14.265 0.595 14.395 0.725 ;
 RECT 6.06 1.49 6.19 1.62 ;
 RECT 13.005 1.28 13.135 1.41 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 23.83 2.64 23.96 2.77 ;
 RECT 23.36 1.72 23.49 1.85 ;
 RECT 23.36 0.73 23.49 0.86 ;
 RECT 20.79 0.935 20.92 1.065 ;
 RECT 21.28 0.315 21.41 0.445 ;
 RECT 22.3 1.735 22.43 1.865 ;
 RECT 22.775 2.64 22.905 2.77 ;
 RECT 21.795 1.715 21.925 1.845 ;
 RECT 21.27 2.64 21.4 2.77 ;
 RECT 24.3 1.78 24.43 1.91 ;
 RECT 22.3 0.72 22.43 0.85 ;
 RECT 9.7 2.045 9.83 2.175 ;
 RECT 5.215 0.145 5.345 0.275 ;
 RECT 14.265 1.9 14.395 2.03 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 5.37 2.345 5.5 2.475 ;
 RECT 28.025 0.435 28.155 0.565 ;
 RECT 9.97 1.23 10.1 1.36 ;
 RECT 18.79 1.705 18.92 1.835 ;
 RECT 9.16 2.075 9.29 2.205 ;
 RECT 6.81 0.88 6.94 1.01 ;
 RECT 16.82 1.835 16.95 1.965 ;
 RECT 16.69 0.765 16.82 0.895 ;
 RECT 4.63 0.74 4.76 0.87 ;
 RECT 29.64 0.12 29.77 0.25 ;
 RECT 7.415 0.53 7.545 0.66 ;
 RECT 15.665 2.38 15.795 2.51 ;
 RECT 11.94 0.905 12.07 1.035 ;
 RECT 26.775 1.425 26.905 1.555 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 19.855 0.92 19.985 1.05 ;
 RECT 27.245 1.475 27.375 1.605 ;
 RECT 13.74 0.875 13.87 1.005 ;
 RECT 5.945 0.79 6.075 0.92 ;
 RECT 17.76 1.835 17.89 1.965 ;
 RECT 6.79 2.07 6.92 2.2 ;
 RECT 31.2 1.475 31.33 1.605 ;
 RECT 4.16 0.74 4.29 0.87 ;
 RECT 5.88 1.825 6.01 1.955 ;
 RECT 13.74 1.945 13.87 2.075 ;
 RECT 4.63 2.05 4.76 2.18 ;
 RECT 26.525 0.505 26.655 0.635 ;
 RECT 11.015 2.015 11.145 2.145 ;
 RECT 28.46 0.12 28.59 0.25 ;
 RECT 28.025 1.485 28.155 1.615 ;
 RECT 30.42 1.465 30.55 1.595 ;
 RECT 19.26 1.705 19.39 1.835 ;
 RECT 30.42 0.595 30.55 0.725 ;
 RECT 7.09 1.525 7.22 1.655 ;
 RECT 12.64 2.44 12.77 2.57 ;
 RECT 4.16 2.115 4.29 2.245 ;
 RECT 19.735 1.705 19.865 1.835 ;
 RECT 29.105 1.405 29.235 1.535 ;
 RECT 11.02 0.905 11.15 1.035 ;
 RECT 4.23 0.325 4.36 0.455 ;
 RECT 9.16 0.315 9.29 0.445 ;
 RECT 11.495 0.905 11.625 1.035 ;
 RECT 14.77 0.595 14.9 0.725 ;
 RECT 12.83 0.6 12.96 0.73 ;
 RECT 28.63 1.445 28.76 1.575 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 17.795 1.035 17.925 1.165 ;
 RECT 18.38 0.91 18.51 1.04 ;
 RECT 10.19 2.435 10.32 2.565 ;
 RECT 8.68 2.135 8.81 2.265 ;
 RECT 6.295 2.105 6.425 2.235 ;
 RECT 7.26 2.11 7.39 2.24 ;
 RECT 2.85 0.285 2.98 0.415 ;
 RECT 3.295 1.155 3.425 1.285 ;
 RECT 22.625 1.3 22.755 1.43 ;
 LAYER M1 ;
 RECT 29.08 0.22 29.31 0.29 ;
 RECT 30.73 0.85 30.87 1.385 ;
 RECT 30.415 1.525 30.555 1.73 ;
 RECT 29.31 0.71 30.87 0.85 ;
 RECT 30.415 0.51 30.555 0.71 ;
 RECT 30.415 1.385 30.87 1.525 ;
 RECT 26.32 1.225 26.55 1.245 ;
 RECT 26.32 1.195 26.91 1.225 ;
 RECT 26.46 1.015 26.77 1.035 ;
 RECT 26.32 1.035 26.77 1.055 ;
 RECT 26.595 0.64 26.735 1.015 ;
 RECT 26.77 1.225 26.91 1.75 ;
 RECT 26.475 0.5 26.735 0.64 ;
 RECT 27.37 1.035 27.6 1.055 ;
 RECT 27.37 1.195 27.6 1.245 ;
 RECT 26.32 1.055 27.6 1.195 ;
 RECT 28.34 1.145 28.48 1.345 ;
 RECT 28.02 1.485 28.16 1.76 ;
 RECT 28.34 0.73 28.48 0.935 ;
 RECT 28.02 0.355 28.16 0.59 ;
 RECT 28.02 1.345 28.48 1.485 ;
 RECT 28.295 0.935 28.525 1.145 ;
 RECT 28.02 0.59 28.48 0.73 ;
 RECT 25.28 0.36 25.51 0.43 ;
 RECT 26.875 0.36 27.015 0.565 ;
 RECT 25.28 0.22 27.015 0.36 ;
 RECT 27.615 0.705 27.755 0.75 ;
 RECT 27.74 0.995 28.045 1.205 ;
 RECT 27.74 0.89 27.88 0.995 ;
 RECT 27.615 0.75 27.88 0.89 ;
 RECT 26.875 0.565 27.755 0.705 ;
 RECT 14.765 0.525 14.905 0.885 ;
 RECT 14.765 1.095 14.905 2.065 ;
 RECT 14.765 0.885 15.04 1.095 ;
 RECT 18.81 0.775 18.95 1.405 ;
 RECT 19.535 0.56 19.765 0.635 ;
 RECT 17.79 1.405 18.95 1.545 ;
 RECT 17.79 1.545 17.93 1.83 ;
 RECT 16.745 1.83 17.995 1.97 ;
 RECT 17.79 1.17 17.93 1.405 ;
 RECT 17.72 1.03 18 1.17 ;
 RECT 21.685 0.38 21.825 0.635 ;
 RECT 18.81 0.635 21.825 0.775 ;
 RECT 22.575 0.38 22.715 1.26 ;
 RECT 21.685 0.24 22.715 0.38 ;
 RECT 22.575 1.26 22.805 1.47 ;
 RECT 17.07 0.57 17.3 0.95 ;
 RECT 20.145 0.22 20.375 0.28 ;
 RECT 20.145 0.42 20.375 0.43 ;
 RECT 17.915 0.28 20.375 0.42 ;
 RECT 17.915 0.42 18.145 0.6 ;
 RECT 15.49 0.585 16.445 0.63 ;
 RECT 16.215 0.63 16.445 0.665 ;
 RECT 16.215 0.455 16.445 0.49 ;
 RECT 15.515 0.49 16.445 0.585 ;
 RECT 15.49 0.63 15.72 0.795 ;
 RECT 11.49 1.04 11.63 2.34 ;
 RECT 11.49 0.895 11.63 0.9 ;
 RECT 11.42 0.9 11.695 1.04 ;
 RECT 12.285 2.16 12.425 2.34 ;
 RECT 11.49 2.34 12.425 2.48 ;
 RECT 14.26 2.055 14.4 2.11 ;
 RECT 13.735 0.765 13.875 1.915 ;
 RECT 14.26 0.525 14.4 1.915 ;
 RECT 12.285 2.02 14.41 2.055 ;
 RECT 12.285 2.055 13.875 2.16 ;
 RECT 13.735 1.915 14.41 2.02 ;
 RECT 5.94 1.67 6.08 1.82 ;
 RECT 5.94 1.96 6.08 2.51 ;
 RECT 5.94 0.5 6.08 1.44 ;
 RECT 5.94 1.44 6.195 1.67 ;
 RECT 5.81 1.82 6.08 1.96 ;
 RECT 8.3 2.445 8.53 2.51 ;
 RECT 8.3 2.65 8.53 2.655 ;
 RECT 5.94 2.51 8.53 2.65 ;
 RECT 7.085 0.66 7.225 0.895 ;
 RECT 6.625 0.52 7.225 0.66 ;
 RECT 7.085 0.895 10.77 1.035 ;
 RECT 10.54 1.035 10.77 1.105 ;
 RECT 5.185 0.88 5.325 1.475 ;
 RECT 5.145 1.63 5.285 1.99 ;
 RECT 5.145 1.475 5.49 1.63 ;
 RECT 5.035 1.99 5.285 2.13 ;
 RECT 5.185 0.74 5.505 0.88 ;
 RECT 2.87 0.87 3.01 1.15 ;
 RECT 2.87 1.29 3.01 2.07 ;
 RECT 2.36 2.07 3.01 2.21 ;
 RECT 2.165 0.73 3.01 0.87 ;
 RECT 3.245 1.115 3.475 1.15 ;
 RECT 3.245 1.29 3.475 1.325 ;
 RECT 2.87 1.15 3.475 1.29 ;
 RECT 3.935 1.335 4.075 2.11 ;
 RECT 3.935 2.25 4.075 2.255 ;
 RECT 3.935 0.875 4.075 1.195 ;
 RECT 3.935 2.11 4.36 2.25 ;
 RECT 3.935 0.735 4.36 0.875 ;
 RECT 3.935 1.195 5.045 1.335 ;
 RECT 4.905 0.6 5.045 1.195 ;
 RECT 6.335 0.36 6.475 2.035 ;
 RECT 5.65 0.22 6.475 0.36 ;
 RECT 5.65 0.36 5.79 0.46 ;
 RECT 6.29 2.17 6.43 2.305 ;
 RECT 6.29 2.035 6.475 2.17 ;
 RECT 4.905 0.46 5.79 0.6 ;
 RECT 3.65 0.46 3.79 2.21 ;
 RECT 4.12 0.22 4.485 0.32 ;
 RECT 4.12 0.46 4.485 0.525 ;
 RECT 3.65 0.32 4.485 0.46 ;
 RECT 0.8 0.68 0.94 1.155 ;
 RECT 0.8 1.295 0.94 2.23 ;
 RECT 1.585 0.385 1.725 1.155 ;
 RECT 0.8 1.155 1.725 1.295 ;
 RECT 2.8 0.385 3.03 0.455 ;
 RECT 1.585 0.245 3.03 0.385 ;
 RECT 16.18 1.895 16.32 2.39 ;
 RECT 20.325 2.205 20.465 2.39 ;
 RECT 16.18 2.39 20.465 2.53 ;
 RECT 15.055 1.755 16.32 1.895 ;
 RECT 15.055 1.895 15.195 2.34 ;
 RECT 13.785 2.3 14.015 2.34 ;
 RECT 13.785 2.48 14.015 2.51 ;
 RECT 13.785 2.34 15.195 2.48 ;
 RECT 20.325 2.065 26.055 2.205 ;
 RECT 25.915 2.205 26.055 2.52 ;
 RECT 30.255 2.48 30.395 2.52 ;
 RECT 25.915 2.52 30.395 2.66 ;
 RECT 30.255 2.27 30.485 2.48 ;
 RECT 19.815 1.055 19.955 1.245 ;
 RECT 19.255 1.385 19.395 1.625 ;
 RECT 20.095 1.385 20.325 1.455 ;
 RECT 19.255 1.245 20.325 1.385 ;
 RECT 19.785 0.915 20.085 1.055 ;
 RECT 19.225 1.625 19.48 1.92 ;
 RECT 19.62 1.7 19.915 1.84 ;
 RECT 19.62 1.84 19.76 2.075 ;
 RECT 18.925 1.84 19.065 2.075 ;
 RECT 18.73 1.7 19.065 1.84 ;
 RECT 18.925 2.075 19.76 2.215 ;
 RECT 16.46 1.56 16.6 2.11 ;
 RECT 15.41 1.405 15.64 1.42 ;
 RECT 15.41 1.56 15.64 1.615 ;
 RECT 15.41 1.42 16.6 1.56 ;
 RECT 16.46 2.11 18.785 2.245 ;
 RECT 16.46 2.245 18.78 2.25 ;
 RECT 18.555 2.035 18.785 2.11 ;
 RECT 11.935 1.685 12.075 1.71 ;
 RECT 11.935 1.85 12.075 2.18 ;
 RECT 11.935 0.83 12.075 1.475 ;
 RECT 11.775 1.475 12.075 1.685 ;
 RECT 11.935 1.71 13.14 1.85 ;
 RECT 13 1.415 13.14 1.71 ;
 RECT 12.93 1.275 13.205 1.415 ;
 RECT 7.19 2.105 8.41 2.245 ;
 RECT 7.75 1.365 7.89 1.5 ;
 RECT 6.92 1.64 7.425 1.675 ;
 RECT 6.92 1.5 7.89 1.64 ;
 RECT 9.695 1.365 9.835 2.25 ;
 RECT 11.01 1.04 11.15 1.25 ;
 RECT 11.01 1.39 11.15 2.215 ;
 RECT 11.01 0.885 11.15 0.9 ;
 RECT 7.75 1.25 11.15 1.365 ;
 RECT 7.75 1.225 10.4 1.25 ;
 RECT 10.26 1.365 11.15 1.39 ;
 RECT 10.945 0.9 11.22 1.04 ;
 RECT 6.63 1.82 8.21 1.96 ;
 RECT 8.07 1.79 8.21 1.82 ;
 RECT 6.63 1.22 6.945 1.36 ;
 RECT 6.805 0.805 6.945 1.22 ;
 RECT 6.715 1.96 6.995 2.215 ;
 RECT 6.63 1.36 6.77 1.82 ;
 RECT 9.27 1.615 9.5 1.65 ;
 RECT 9.27 1.79 9.5 1.825 ;
 RECT 8.07 1.65 9.505 1.79 ;
 RECT 28.96 0.73 29.1 1.04 ;
 RECT 29.1 1.18 29.24 1.605 ;
 RECT 28.895 0.59 29.17 0.73 ;
 RECT 30.22 0.99 30.45 1.04 ;
 RECT 28.96 1.04 30.45 1.18 ;
 RECT 30.22 1.18 30.45 1.2 ;
 RECT 29.08 0.29 29.45 0.43 ;
 RECT 29.31 0.43 29.45 0.71 ;
 END
END RSDFFNSRASRX2

MACRO RSDFFNSRASX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 31.04 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 24.225 0.59 24.595 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 29.455 1.435 29.795 1.8 ;
 RECT 27.775 1.99 29.64 2.13 ;
 RECT 25.545 2.22 27.915 2.36 ;
 RECT 27.775 1.435 27.915 1.99 ;
 RECT 29.5 1.8 29.64 1.99 ;
 RECT 25.545 1.39 25.685 2.22 ;
 RECT 26.93 1.37 27.07 2.22 ;
 RECT 27.775 2.13 27.915 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 5.155 0.08 5.435 0.295 ;
 RECT 27.895 0.08 28.135 0.26 ;
 RECT 12.765 0.59 13.04 0.73 ;
 RECT 9.085 0.31 9.375 0.45 ;
 RECT 16.695 0.275 17.72 0.415 ;
 RECT 21.055 0.335 21.32 0.495 ;
 RECT 17.58 0.75 18.525 0.89 ;
 RECT 0 -0.08 31.04 0.08 ;
 RECT 3.19 0.08 3.33 0.74 ;
 RECT 0.31 0.08 0.45 0.775 ;
 RECT 1.28 0.08 1.42 0.93 ;
 RECT 7.98 0.08 8.215 0.46 ;
 RECT 4.635 0.08 4.775 0.97 ;
 RECT 16.695 0.415 16.835 0.945 ;
 RECT 22.7 0.08 22.84 0.82 ;
 RECT 25.545 0.08 25.685 0.36 ;
 RECT 26.76 0.08 26.9 0.35 ;
 RECT 18.385 0.89 18.525 1.11 ;
 RECT 17.58 0.415 17.72 0.75 ;
 RECT 12.835 0.08 12.975 0.59 ;
 RECT 9.165 0.08 9.305 0.31 ;
 RECT 16.695 0.08 16.835 0.275 ;
 RECT 21.11 0.08 21.25 0.335 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.51 1.205 20.845 1.445 ;
 RECT 20.62 0.915 20.76 1.205 ;
 RECT 21.625 1.84 21.765 1.885 ;
 RECT 21.625 0.915 21.765 1.7 ;
 RECT 20.62 1.84 20.76 1.885 ;
 RECT 20.62 1.7 21.765 1.84 ;
 RECT 20.62 1.445 20.76 1.7 ;
 END
 ANTENNADIFFAREA 0.433 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 20.965 2.6 21.23 2.8 ;
 RECT 22.555 2.6 22.82 2.8 ;
 RECT 12.58 2.215 12.855 2.355 ;
 RECT 0 2.8 31.04 2.96 ;
 RECT 1.28 1.965 1.42 2.8 ;
 RECT 3.19 1.99 3.33 2.8 ;
 RECT 0.31 1.74 0.45 2.8 ;
 RECT 5.31 2.34 5.56 2.8 ;
 RECT 4.635 1.98 4.775 2.8 ;
 RECT 9.165 2.195 9.305 2.8 ;
 RECT 10.195 2.23 10.335 2.8 ;
 RECT 15.605 2.335 15.875 2.8 ;
 RECT 12.645 2.355 12.785 2.8 ;
 RECT 12.645 2.195 12.785 2.215 ;
 RECT 8.685 2.645 8.825 2.8 ;
 RECT 8.685 2.435 9.015 2.645 ;
 RECT 8.685 2.07 8.825 2.435 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.685 1.475 5.015 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.02 1.095 22.28 1.335 ;
 RECT 22.14 0.51 22.28 1.095 ;
 RECT 23.2 1.905 23.34 1.91 ;
 RECT 22.14 1.765 23.34 1.905 ;
 RECT 23.2 0.56 23.34 1.765 ;
 RECT 22.14 1.905 22.28 1.915 ;
 RECT 22.14 1.335 22.28 1.765 ;
 END
 ANTENNADIFFAREA 0.73 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.225 1.16 12.6 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.985 1.79 10.36 2.04 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.1 1.435 1.625 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.79 1.59 2.735 1.75 ;
 RECT 1.885 1.09 2.025 1.44 ;
 RECT 1.79 1.44 2.035 1.59 ;
 RECT 2.585 1.75 2.725 1.805 ;
 RECT 2.585 1.53 2.725 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.25 1.115 2.67 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 OBS
 LAYER PO ;
 RECT 16.225 0.535 16.455 0.665 ;
 RECT 17.08 0.535 17.31 0.835 ;
 RECT 17.08 0.835 17.18 2.39 ;
 RECT 26.11 0.215 26.21 0.995 ;
 RECT 26.11 0.995 26.35 1.205 ;
 RECT 26.11 1.205 26.21 2 ;
 RECT 28.505 0.375 28.605 0.99 ;
 RECT 28.505 0.99 28.755 1.2 ;
 RECT 28.505 1.2 28.605 2.27 ;
 RECT 28.505 2.27 28.79 2.48 ;
 RECT 13.49 0.655 13.59 2.305 ;
 RECT 13.795 2.3 14.025 2.305 ;
 RECT 13.795 2.405 14.025 2.51 ;
 RECT 13.49 2.305 14.025 2.405 ;
 RECT 25.33 0.21 25.43 0.755 ;
 RECT 25.33 0.855 25.43 2.2 ;
 RECT 28.195 1.125 28.295 2.2 ;
 RECT 24.365 0.755 25.9 0.84 ;
 RECT 24.365 0.84 25.895 0.855 ;
 RECT 25.8 0.215 25.9 0.755 ;
 RECT 24.365 0.595 24.595 0.755 ;
 RECT 25.33 2.2 28.295 2.3 ;
 RECT 12.2 1.28 12.455 1.45 ;
 RECT 12.2 1.45 12.3 1.655 ;
 RECT 12.2 0.655 12.3 1.18 ;
 RECT 12.2 1.655 13.16 1.755 ;
 RECT 13.06 1.755 13.16 2.355 ;
 RECT 11.285 0.66 11.385 1.18 ;
 RECT 12.2 1.755 12.3 2.51 ;
 RECT 11.285 1.24 12.455 1.28 ;
 RECT 11.285 1.18 12.3 1.24 ;
 RECT 27.02 0.38 27.12 0.96 ;
 RECT 27.02 1.06 27.12 1.14 ;
 RECT 26.6 0.935 26.83 0.96 ;
 RECT 26.6 0.96 27.12 1.06 ;
 RECT 26.6 1.06 26.83 1.145 ;
 RECT 27.02 1.14 27.29 1.24 ;
 RECT 27.19 1.24 27.29 1.84 ;
 RECT 27.385 0.22 27.615 0.28 ;
 RECT 27.385 0.38 27.615 0.43 ;
 RECT 27.02 0.28 27.615 0.38 ;
 RECT 11.275 1.575 11.375 2.485 ;
 RECT 11.785 1.575 12.015 1.685 ;
 RECT 11.275 1.475 12.015 1.575 ;
 RECT 29.205 0.195 29.305 2.665 ;
 RECT 28.195 0.095 29.305 0.195 ;
 RECT 24.57 1.245 24.67 2.665 ;
 RECT 28.195 0.195 28.295 0.945 ;
 RECT 24.57 1.2 24.855 1.245 ;
 RECT 24.625 1.035 24.855 1.1 ;
 RECT 24.57 2.665 29.305 2.765 ;
 RECT 24.57 1.1 24.9 1.2 ;
 RECT 15.5 0.795 15.665 0.925 ;
 RECT 14.82 0.885 15.05 0.925 ;
 RECT 14.82 1.025 15.05 1.095 ;
 RECT 14.82 0.925 15.665 1.025 ;
 RECT 15.5 0.585 15.73 0.795 ;
 RECT 2.535 1.55 2.775 1.78 ;
 RECT 2.675 1.78 2.775 2.695 ;
 RECT 1.065 1.435 1.635 1.71 ;
 RECT 1.065 0.515 1.165 1.435 ;
 RECT 1.065 1.71 1.165 2.645 ;
 RECT 1.535 0.515 1.635 1.435 ;
 RECT 1.535 1.71 1.635 2.695 ;
 RECT 2.255 1.37 2.355 1.605 ;
 RECT 2.485 0.515 2.585 1.14 ;
 RECT 2.205 1.705 2.305 2.695 ;
 RECT 2.205 1.605 2.355 1.705 ;
 RECT 2.255 1.14 2.585 1.37 ;
 RECT 1.87 0.515 1.97 1.105 ;
 RECT 1.83 1.105 2.075 1.345 ;
 RECT 4.42 0.52 4.52 2.465 ;
 RECT 4.18 0.27 4.52 0.52 ;
 RECT 7.05 1.33 7.19 1.475 ;
 RECT 7.05 1.71 7.15 2.475 ;
 RECT 7.09 0.65 7.19 1.33 ;
 RECT 7.05 1.475 7.28 1.71 ;
 RECT 6.6 0.705 6.7 1.165 ;
 RECT 6.16 1.27 6.26 1.445 ;
 RECT 6.6 0.47 6.885 0.705 ;
 RECT 6.16 1.17 6.7 1.265 ;
 RECT 6.16 1.265 6.535 1.27 ;
 RECT 6.39 1.165 6.7 1.17 ;
 RECT 6.015 1.445 6.26 1.69 ;
 RECT 7.49 0.715 7.59 1.61 ;
 RECT 7.525 1.71 7.625 2.48 ;
 RECT 7.49 1.61 7.625 1.71 ;
 RECT 7.37 0.485 7.61 0.715 ;
 RECT 13.095 0.655 13.195 1.24 ;
 RECT 12.965 1.24 13.195 1.475 ;
 RECT 4.895 0.49 4.995 1.495 ;
 RECT 4.7 1.495 4.995 1.745 ;
 RECT 4.895 1.745 4.995 2.37 ;
 RECT 8.74 0.74 8.84 1.51 ;
 RECT 8.95 1.61 9.05 2.435 ;
 RECT 8.785 2.435 9.05 2.645 ;
 RECT 8.675 0.53 8.905 0.74 ;
 RECT 8.74 1.51 9.05 1.61 ;
 RECT 2.975 0.135 3.075 0.22 ;
 RECT 2.815 0.22 3.075 0.43 ;
 RECT 2.975 0.43 3.075 2.695 ;
 RECT 3.445 0.295 3.545 1.115 ;
 RECT 3.28 1.115 3.545 1.325 ;
 RECT 3.445 1.325 3.545 2.74 ;
 RECT 19.52 0.77 19.62 2.155 ;
 RECT 19.52 0.55 19.62 0.56 ;
 RECT 19.52 0.56 19.775 0.77 ;
 RECT 20.885 0.39 20.985 1.4 ;
 RECT 20.155 0.43 20.255 1.245 ;
 RECT 21.375 0.51 21.475 1.4 ;
 RECT 21.375 1.5 21.475 2.26 ;
 RECT 20.885 1.5 20.985 2.235 ;
 RECT 20.09 0.22 20.32 0.29 ;
 RECT 20.09 0.39 20.32 0.43 ;
 RECT 20.09 0.29 20.985 0.39 ;
 RECT 20.885 1.4 21.475 1.5 ;
 RECT 20.105 1.245 20.335 1.455 ;
 RECT 8.31 2.445 8.57 2.655 ;
 RECT 8.47 1.79 8.57 2.445 ;
 RECT 18.58 1.445 18.68 2.035 ;
 RECT 18.565 2.035 18.795 2.245 ;
 RECT 19.05 0.55 19.15 2.69 ;
 RECT 9.98 1.58 10.08 1.79 ;
 RECT 9.72 1.01 9.82 1.48 ;
 RECT 9.98 2 10.08 2.69 ;
 RECT 9.98 1.79 10.215 2 ;
 RECT 9.72 1.48 10.08 1.58 ;
 RECT 9.98 2.69 19.15 2.79 ;
 RECT 9.42 0.98 9.52 1.615 ;
 RECT 9.28 1.615 9.52 1.825 ;
 RECT 9.42 1.825 9.52 2.675 ;
 RECT 22.4 1.33 23.08 1.43 ;
 RECT 22.4 1.43 22.65 1.46 ;
 RECT 22.4 1.25 22.65 1.33 ;
 RECT 22.98 0.375 23.08 1.33 ;
 RECT 22.4 0.385 22.5 1.25 ;
 RECT 22.4 1.46 22.5 2.69 ;
 RECT 22.98 1.43 23.08 2.695 ;
 RECT 23.585 0.22 23.815 0.275 ;
 RECT 23.585 0.375 23.815 0.43 ;
 RECT 22.98 0.275 23.815 0.375 ;
 RECT 17.55 0.73 17.65 1.39 ;
 RECT 17.415 1.39 17.65 1.6 ;
 RECT 17.55 1.6 17.65 2.39 ;
 RECT 5.735 0.285 5.835 1.52 ;
 RECT 5.235 1.52 5.835 1.62 ;
 RECT 5.735 0.185 14.625 0.195 ;
 RECT 7.79 0.095 14.625 0.185 ;
 RECT 5.735 0.195 7.89 0.285 ;
 RECT 14.525 0.195 14.625 1.29 ;
 RECT 15.42 1.39 15.615 1.405 ;
 RECT 6.555 1.565 6.655 2.675 ;
 RECT 5.67 1.62 5.77 2.675 ;
 RECT 5.235 1.44 5.48 1.52 ;
 RECT 5.235 1.62 5.48 1.69 ;
 RECT 7.79 0.285 7.89 1.24 ;
 RECT 14.525 1.29 15.615 1.39 ;
 RECT 5.67 2.675 6.655 2.775 ;
 RECT 15.42 1.405 15.65 1.615 ;
 RECT 25.805 1.245 25.905 2.02 ;
 RECT 25.675 1.035 25.905 1.245 ;
 RECT 15.915 0.105 18.74 0.205 ;
 RECT 15.915 0.205 16.015 1.91 ;
 RECT 18.64 0.205 18.74 1.265 ;
 RECT 15.095 1.71 15.195 1.91 ;
 RECT 14.01 1.61 15.195 1.71 ;
 RECT 14.01 0.475 14.11 1.61 ;
 RECT 14.56 1.71 14.66 2.425 ;
 RECT 10.675 0.475 10.775 0.895 ;
 RECT 15.095 1.91 16.015 2.01 ;
 RECT 10.675 0.375 14.11 0.475 ;
 RECT 10.55 0.895 10.78 1.105 ;
 RECT 16.225 0.455 18.155 0.535 ;
 RECT 17.925 0.535 18.155 0.6 ;
 RECT 17.925 0.39 18.155 0.435 ;
 RECT 16.305 0.435 18.155 0.455 ;
 LAYER CO ;
 RECT 28.61 2.31 28.74 2.44 ;
 RECT 13.845 2.34 13.975 2.47 ;
 RECT 24.415 0.635 24.545 0.765 ;
 RECT 12.275 1.28 12.405 1.41 ;
 RECT 27.435 0.26 27.565 0.39 ;
 RECT 11.835 1.515 11.965 1.645 ;
 RECT 24.675 1.075 24.805 1.205 ;
 RECT 14.87 0.925 15 1.055 ;
 RECT 1.29 1.51 1.42 1.64 ;
 RECT 0.815 0.735 0.945 0.865 ;
 RECT 3.195 2.31 3.325 2.44 ;
 RECT 1.285 2.015 1.415 2.145 ;
 RECT 1.89 1.155 2.02 1.285 ;
 RECT 3.195 2.05 3.325 2.18 ;
 RECT 2.59 1.6 2.72 1.73 ;
 RECT 3.665 2.01 3.795 2.14 ;
 RECT 3.665 0.735 3.795 0.865 ;
 RECT 2.425 2.075 2.555 2.205 ;
 RECT 1.285 2.275 1.415 2.405 ;
 RECT 3.195 0.545 3.325 0.675 ;
 RECT 3.665 1.75 3.795 1.88 ;
 RECT 0.815 2.015 0.945 2.145 ;
 RECT 2.23 0.735 2.36 0.865 ;
 RECT 2.41 1.19 2.54 1.32 ;
 RECT 7.1 1.525 7.23 1.655 ;
 RECT 12.65 2.225 12.78 2.355 ;
 RECT 21.63 0.975 21.76 1.105 ;
 RECT 22.62 2.64 22.75 2.77 ;
 RECT 4.17 2.115 4.3 2.245 ;
 RECT 21.115 0.36 21.245 0.49 ;
 RECT 23.205 0.63 23.335 0.76 ;
 RECT 27.27 0.595 27.4 0.725 ;
 RECT 6.705 0.525 6.835 0.655 ;
 RECT 7.75 1.825 7.88 1.955 ;
 RECT 27.78 1.49 27.91 1.62 ;
 RECT 6.35 0.88 6.48 1.01 ;
 RECT 14.78 1.87 14.91 2 ;
 RECT 8.22 2.11 8.35 2.24 ;
 RECT 8.035 0.32 8.165 0.45 ;
 RECT 25.55 0.135 25.68 0.265 ;
 RECT 5.295 1.495 5.425 1.625 ;
 RECT 5.245 0.745 5.375 0.875 ;
 RECT 5.115 1.995 5.245 2.125 ;
 RECT 11.95 1.995 12.08 2.125 ;
 RECT 0.315 0.59 0.445 0.72 ;
 RECT 11.505 2.07 11.635 2.2 ;
 RECT 14.275 0.595 14.405 0.725 ;
 RECT 6.07 1.49 6.2 1.62 ;
 RECT 13.015 1.28 13.145 1.41 ;
 RECT 22.145 1.725 22.275 1.855 ;
 RECT 0.315 2.085 0.445 2.215 ;
 RECT 9.71 2.235 9.84 2.365 ;
 RECT 5.225 0.145 5.355 0.275 ;
 RECT 14.275 1.9 14.405 2.03 ;
 RECT 0.315 2.345 0.445 2.475 ;
 RECT 5.38 2.345 5.51 2.475 ;
 RECT 26.33 0.435 26.46 0.565 ;
 RECT 20.625 1.705 20.755 1.835 ;
 RECT 9.98 1.23 10.11 1.36 ;
 RECT 18.8 1.705 18.93 1.835 ;
 RECT 9.17 2.265 9.3 2.395 ;
 RECT 6.82 0.88 6.95 1.01 ;
 RECT 16.83 1.835 16.96 1.965 ;
 RECT 16.7 0.765 16.83 0.895 ;
 RECT 4.64 0.74 4.77 0.87 ;
 RECT 27.945 0.12 28.075 0.25 ;
 RECT 7.425 0.53 7.555 0.66 ;
 RECT 22.145 0.62 22.275 0.75 ;
 RECT 15.675 2.38 15.805 2.51 ;
 RECT 11.95 0.885 12.08 1.015 ;
 RECT 25.08 1.425 25.21 1.555 ;
 RECT 0.315 0.33 0.445 0.46 ;
 RECT 19.865 0.92 19.995 1.05 ;
 RECT 25.55 1.475 25.68 1.605 ;
 RECT 13.75 0.875 13.88 1.005 ;
 RECT 5.955 0.79 6.085 0.92 ;
 RECT 17.77 1.835 17.9 1.965 ;
 RECT 6.8 2.07 6.93 2.2 ;
 RECT 29.505 1.475 29.635 1.605 ;
 RECT 21.63 1.705 21.76 1.835 ;
 RECT 23.205 1.71 23.335 1.84 ;
 RECT 20.625 0.975 20.755 1.105 ;
 RECT 4.17 0.74 4.3 0.87 ;
 RECT 5.89 1.825 6.02 1.955 ;
 RECT 13.75 1.945 13.88 2.075 ;
 RECT 4.64 2.05 4.77 2.18 ;
 RECT 24.83 0.505 24.96 0.635 ;
 RECT 11.025 2.015 11.155 2.145 ;
 RECT 26.765 0.12 26.895 0.25 ;
 RECT 26.33 1.485 26.46 1.615 ;
 RECT 28.725 1.465 28.855 1.595 ;
 RECT 19.27 1.705 19.4 1.835 ;
 RECT 28.725 0.595 28.855 0.725 ;
 RECT 19.745 1.705 19.875 1.835 ;
 RECT 21.03 2.64 21.16 2.77 ;
 RECT 27.41 1.405 27.54 1.535 ;
 RECT 11.03 0.905 11.16 1.035 ;
 RECT 4.24 0.325 4.37 0.455 ;
 RECT 9.17 0.315 9.3 0.445 ;
 RECT 11.505 0.905 11.635 1.035 ;
 RECT 14.78 0.595 14.91 0.725 ;
 RECT 12.84 0.595 12.97 0.725 ;
 RECT 26.935 1.445 27.065 1.575 ;
 RECT 0.315 1.825 0.445 1.955 ;
 RECT 17.805 1.035 17.935 1.165 ;
 RECT 18.39 0.91 18.52 1.04 ;
 RECT 10.2 2.3 10.33 2.43 ;
 RECT 22.705 0.62 22.835 0.75 ;
 RECT 8.69 2.135 8.82 2.265 ;
 RECT 6.305 2.105 6.435 2.235 ;
 RECT 7.27 2.11 7.4 2.24 ;
 RECT 8.725 0.57 8.855 0.7 ;
 RECT 8.835 2.475 8.965 2.605 ;
 RECT 2.865 0.26 2.995 0.39 ;
 RECT 3.33 1.155 3.46 1.285 ;
 RECT 22.47 1.29 22.6 1.42 ;
 RECT 20.155 1.285 20.285 1.415 ;
 RECT 17.975 0.43 18.105 0.56 ;
 RECT 19.595 0.6 19.725 0.73 ;
 RECT 20.14 0.26 20.27 0.39 ;
 RECT 8.36 2.485 8.49 2.615 ;
 RECT 18.615 2.075 18.745 2.205 ;
 RECT 10.035 1.83 10.165 1.96 ;
 RECT 9.33 1.655 9.46 1.785 ;
 RECT 23.635 0.26 23.765 0.39 ;
 RECT 28.575 1.03 28.705 1.16 ;
 RECT 16.275 0.495 16.405 0.625 ;
 RECT 17.465 1.43 17.595 1.56 ;
 RECT 15.55 0.625 15.68 0.755 ;
 RECT 15.47 1.445 15.6 1.575 ;
 RECT 25.725 1.075 25.855 1.205 ;
 RECT 10.6 0.935 10.73 1.065 ;
 RECT 26.65 0.975 26.78 1.105 ;
 RECT 17.13 0.665 17.26 0.795 ;
 RECT 26.17 1.035 26.3 1.165 ;
 RECT 4.76 1.55 4.89 1.68 ;
 RECT 1.285 0.735 1.415 0.865 ;
 LAYER M1 ;
 RECT 3.28 1.115 3.51 1.15 ;
 RECT 3.28 1.29 3.51 1.325 ;
 RECT 27.265 0.73 27.405 1.04 ;
 RECT 27.405 1.18 27.545 1.605 ;
 RECT 27.2 0.59 27.475 0.73 ;
 RECT 28.525 0.99 28.755 1.04 ;
 RECT 27.265 1.04 28.755 1.18 ;
 RECT 28.525 1.18 28.755 1.2 ;
 RECT 27.385 0.29 27.755 0.43 ;
 RECT 27.615 0.43 27.755 0.71 ;
 RECT 27.385 0.22 27.615 0.29 ;
 RECT 29.035 0.85 29.175 1.385 ;
 RECT 28.72 1.525 28.86 1.73 ;
 RECT 27.615 0.71 29.175 0.85 ;
 RECT 28.72 0.51 28.86 0.71 ;
 RECT 28.72 1.385 29.175 1.525 ;
 RECT 24.625 1.225 24.855 1.245 ;
 RECT 24.625 1.195 25.215 1.225 ;
 RECT 24.765 1.015 25.075 1.035 ;
 RECT 24.625 1.035 25.075 1.055 ;
 RECT 24.9 0.64 25.04 1.015 ;
 RECT 25.075 1.225 25.215 1.75 ;
 RECT 24.78 0.5 25.04 0.64 ;
 RECT 25.675 1.035 25.905 1.055 ;
 RECT 25.675 1.195 25.905 1.245 ;
 RECT 24.625 1.055 25.905 1.195 ;
 RECT 26.645 1.145 26.785 1.345 ;
 RECT 26.325 1.485 26.465 1.76 ;
 RECT 26.645 0.73 26.785 0.935 ;
 RECT 26.325 0.355 26.465 0.59 ;
 RECT 26.325 1.345 26.785 1.485 ;
 RECT 26.6 0.935 26.83 1.145 ;
 RECT 26.325 0.59 26.785 0.73 ;
 RECT 23.585 0.36 23.815 0.43 ;
 RECT 25.18 0.36 25.32 0.565 ;
 RECT 23.585 0.22 25.32 0.36 ;
 RECT 25.92 0.705 26.06 0.75 ;
 RECT 26.045 0.995 26.35 1.205 ;
 RECT 26.045 0.89 26.185 0.995 ;
 RECT 25.92 0.75 26.185 0.89 ;
 RECT 25.18 0.565 26.06 0.705 ;
 RECT 18.82 0.775 18.96 1.405 ;
 RECT 19.545 0.56 19.775 0.635 ;
 RECT 17.8 1.405 18.96 1.545 ;
 RECT 17.8 1.545 17.94 1.83 ;
 RECT 17.8 1.17 17.94 1.405 ;
 RECT 16.755 1.83 18.005 1.97 ;
 RECT 17.73 1.03 18.01 1.17 ;
 RECT 21.74 0.36 21.88 0.635 ;
 RECT 18.82 0.635 21.88 0.775 ;
 RECT 22.42 0.36 22.56 1.25 ;
 RECT 22.42 1.25 22.65 1.46 ;
 RECT 21.74 0.22 22.56 0.36 ;
 RECT 17.925 0.28 20.32 0.42 ;
 RECT 17.925 0.42 18.155 0.6 ;
 RECT 20.09 0.22 20.32 0.28 ;
 RECT 20.09 0.42 20.32 0.43 ;
 RECT 11.5 1.04 11.64 2.34 ;
 RECT 11.5 0.895 11.64 0.9 ;
 RECT 11.43 0.9 11.705 1.04 ;
 RECT 12.295 2.055 12.435 2.34 ;
 RECT 11.5 2.34 12.435 2.48 ;
 RECT 12.295 1.915 14.41 2.055 ;
 RECT 13.745 0.765 13.885 1.915 ;
 RECT 13.745 2.055 13.885 2.145 ;
 RECT 14.27 0.525 14.41 1.915 ;
 RECT 14.27 2.055 14.41 2.11 ;
 RECT 14.775 0.525 14.915 0.885 ;
 RECT 14.775 1.095 14.915 2.065 ;
 RECT 14.775 0.885 15.05 1.095 ;
 RECT 15.5 0.585 16.455 0.63 ;
 RECT 16.225 0.63 16.455 0.665 ;
 RECT 16.225 0.455 16.455 0.49 ;
 RECT 15.525 0.49 16.455 0.585 ;
 RECT 15.5 0.63 15.73 0.795 ;
 RECT 17.08 0.57 17.31 0.95 ;
 RECT 5.95 1.67 6.09 1.82 ;
 RECT 5.95 1.96 6.09 2.51 ;
 RECT 8.31 2.445 8.54 2.51 ;
 RECT 8.31 2.65 8.54 2.655 ;
 RECT 5.95 0.5 6.09 1.44 ;
 RECT 5.95 1.44 6.205 1.67 ;
 RECT 5.82 1.82 6.09 1.96 ;
 RECT 5.95 2.51 8.54 2.65 ;
 RECT 3.945 0.875 4.085 1.195 ;
 RECT 3.945 1.335 4.085 2.11 ;
 RECT 3.945 2.25 4.085 2.255 ;
 RECT 3.945 0.735 4.37 0.875 ;
 RECT 3.945 2.11 4.37 2.25 ;
 RECT 3.945 1.195 5.055 1.335 ;
 RECT 4.915 0.6 5.055 1.195 ;
 RECT 6.345 0.36 6.485 2.035 ;
 RECT 5.66 0.36 5.8 0.46 ;
 RECT 5.66 0.22 6.485 0.36 ;
 RECT 6.3 2.17 6.44 2.305 ;
 RECT 4.915 0.46 5.8 0.6 ;
 RECT 6.3 2.035 6.485 2.17 ;
 RECT 7.095 0.895 10.78 1.035 ;
 RECT 10.55 1.035 10.78 1.105 ;
 RECT 7.095 0.66 7.235 0.895 ;
 RECT 6.635 0.52 7.235 0.66 ;
 RECT 7.375 0.73 8.905 0.74 ;
 RECT 8.675 0.53 8.905 0.59 ;
 RECT 7.375 0.485 7.69 0.6 ;
 RECT 17.07 1.23 17.21 1.42 ;
 RECT 15.22 1.09 17.21 1.23 ;
 RECT 15.22 0.385 15.36 1.09 ;
 RECT 13.21 0.385 13.35 0.87 ;
 RECT 13.21 0.255 15.36 0.385 ;
 RECT 13.21 0.245 15.355 0.255 ;
 RECT 12.485 0.87 13.35 1.01 ;
 RECT 12.485 0.73 12.625 0.87 ;
 RECT 7.375 0.6 12.625 0.73 ;
 RECT 8.545 0.59 12.625 0.6 ;
 RECT 17.415 1.39 17.645 1.42 ;
 RECT 17.07 1.42 17.645 1.56 ;
 RECT 17.415 1.56 17.645 1.6 ;
 RECT 4.13 0.22 4.495 0.32 ;
 RECT 3.66 0.32 4.495 0.46 ;
 RECT 4.13 0.46 4.495 0.525 ;
 RECT 3.66 0.46 3.8 2.21 ;
 RECT 0.81 0.68 0.95 1.155 ;
 RECT 0.81 1.295 0.95 2.23 ;
 RECT 1.595 0.36 1.735 1.155 ;
 RECT 0.81 1.155 1.735 1.295 ;
 RECT 2.815 0.36 3.045 0.43 ;
 RECT 1.595 0.22 3.045 0.36 ;
 RECT 19.63 1.7 19.925 1.84 ;
 RECT 19.63 1.84 19.77 2.075 ;
 RECT 18.935 1.84 19.075 2.075 ;
 RECT 18.74 1.7 19.075 1.84 ;
 RECT 18.935 2.075 19.77 2.215 ;
 RECT 19.825 1.055 19.965 1.245 ;
 RECT 19.265 1.385 19.405 1.625 ;
 RECT 20.105 1.385 20.335 1.455 ;
 RECT 19.265 1.245 20.335 1.385 ;
 RECT 19.795 0.915 20.095 1.055 ;
 RECT 19.235 1.625 19.49 1.92 ;
 RECT 20.335 2.205 20.475 2.39 ;
 RECT 16.19 1.895 16.33 2.39 ;
 RECT 16.19 2.39 20.475 2.53 ;
 RECT 15.065 1.755 16.33 1.895 ;
 RECT 15.065 1.895 15.205 2.34 ;
 RECT 13.795 2.3 14.025 2.34 ;
 RECT 13.795 2.48 14.025 2.51 ;
 RECT 13.795 2.34 15.205 2.48 ;
 RECT 20.335 2.065 24.36 2.205 ;
 RECT 24.22 2.205 24.36 2.52 ;
 RECT 28.56 2.48 28.7 2.52 ;
 RECT 24.22 2.52 28.7 2.66 ;
 RECT 28.56 2.27 28.79 2.48 ;
 RECT 16.47 1.56 16.61 2.11 ;
 RECT 16.47 2.11 18.795 2.245 ;
 RECT 16.47 2.245 18.79 2.25 ;
 RECT 18.565 2.035 18.795 2.11 ;
 RECT 15.42 1.405 15.65 1.42 ;
 RECT 15.42 1.56 15.65 1.615 ;
 RECT 15.42 1.42 16.61 1.56 ;
 RECT 11.785 1.475 12.085 1.635 ;
 RECT 11.945 1.02 12.085 1.475 ;
 RECT 11.945 1.775 12.085 2.18 ;
 RECT 11.875 0.88 12.15 1.02 ;
 RECT 11.785 1.635 13.145 1.685 ;
 RECT 13.005 1.415 13.145 1.635 ;
 RECT 11.945 1.685 13.145 1.775 ;
 RECT 12.96 1.275 13.215 1.415 ;
 RECT 7.2 2.105 8.42 2.245 ;
 RECT 9.705 1.365 9.845 2.435 ;
 RECT 7.76 1.365 7.9 1.5 ;
 RECT 6.93 1.64 7.435 1.675 ;
 RECT 6.93 1.5 7.9 1.64 ;
 RECT 11.02 1.04 11.16 1.25 ;
 RECT 11.02 1.39 11.16 2.215 ;
 RECT 11.02 0.885 11.16 0.9 ;
 RECT 7.76 1.25 11.16 1.365 ;
 RECT 7.76 1.225 10.41 1.25 ;
 RECT 10.27 1.365 11.16 1.39 ;
 RECT 10.955 0.9 11.23 1.04 ;
 RECT 5.155 1.475 5.5 1.63 ;
 RECT 5.155 1.63 5.295 1.99 ;
 RECT 5.195 0.88 5.335 1.475 ;
 RECT 5.045 1.99 5.295 2.13 ;
 RECT 5.195 0.74 5.515 0.88 ;
 RECT 6.64 1.82 8.22 1.96 ;
 RECT 8.08 1.79 8.22 1.82 ;
 RECT 6.725 1.96 7.005 2.215 ;
 RECT 6.815 0.805 6.955 1.22 ;
 RECT 6.64 1.22 6.955 1.36 ;
 RECT 6.64 1.36 6.78 1.82 ;
 RECT 9.28 1.615 9.51 1.65 ;
 RECT 9.28 1.79 9.51 1.825 ;
 RECT 8.08 1.65 9.515 1.79 ;
 RECT 2.88 0.87 3.02 1.15 ;
 RECT 2.88 1.29 3.02 2.07 ;
 RECT 2.175 0.73 3.02 0.87 ;
 RECT 2.37 2.07 3.02 2.21 ;
 RECT 2.88 1.15 3.51 1.29 ;
 END
END RSDFFNSRASX1

MACRO RSDFFNSRASX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 32.64 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 25.92 0.59 26.29 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 31.15 1.435 31.49 1.8 ;
 RECT 29.47 1.99 31.335 2.13 ;
 RECT 27.24 2.22 29.61 2.36 ;
 RECT 29.47 1.435 29.61 1.99 ;
 RECT 31.195 1.8 31.335 1.99 ;
 RECT 27.24 1.39 27.38 2.22 ;
 RECT 28.625 1.37 28.765 2.22 ;
 RECT 29.47 2.13 29.61 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 5.145 0.08 5.425 0.295 ;
 RECT 29.59 0.08 29.83 0.26 ;
 RECT 9.075 0.31 9.365 0.45 ;
 RECT 12.76 0.59 13.03 0.73 ;
 RECT 16.685 0.275 17.71 0.415 ;
 RECT 21.22 0.29 21.485 0.45 ;
 RECT 17.57 0.75 18.515 0.89 ;
 RECT 0 -0.08 32.64 0.08 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.625 0.08 4.765 0.97 ;
 RECT 3.18 0.08 3.32 0.74 ;
 RECT 1.27 0.08 1.41 0.93 ;
 RECT 7.97 0.08 8.205 0.46 ;
 RECT 16.685 0.415 16.825 0.945 ;
 RECT 22.855 0.08 22.995 0.92 ;
 RECT 27.24 0.08 27.38 0.36 ;
 RECT 28.455 0.08 28.595 0.35 ;
 RECT 18.375 0.89 18.515 1.11 ;
 RECT 17.57 0.415 17.71 0.75 ;
 RECT 9.155 0.08 9.295 0.31 ;
 RECT 12.825 0.08 12.965 0.59 ;
 RECT 16.685 0.08 16.825 0.275 ;
 RECT 21.275 0.08 21.415 0.29 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 12.57 2.215 12.845 2.355 ;
 RECT 0 2.8 32.64 2.96 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.27 1.965 1.41 2.8 ;
 RECT 3.18 1.99 3.32 2.8 ;
 RECT 4.625 1.98 4.765 2.8 ;
 RECT 5.3 2.34 5.55 2.8 ;
 RECT 8.675 2.45 8.985 2.66 ;
 RECT 8.675 2.07 8.815 2.45 ;
 RECT 9.155 2.13 9.295 2.8 ;
 RECT 12.635 2.195 12.775 2.215 ;
 RECT 10.185 2.355 10.325 2.8 ;
 RECT 15.595 2.335 15.865 2.8 ;
 RECT 21.265 2.58 21.405 2.8 ;
 RECT 22.77 2.56 22.91 2.8 ;
 RECT 23.825 2.57 23.965 2.8 ;
 RECT 8.675 2.66 8.815 2.8 ;
 RECT 12.635 2.355 12.775 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.675 1.475 5.005 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.215 1.16 12.605 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.975 1.725 10.415 2.04 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.435 1.615 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.78 1.59 2.725 1.75 ;
 RECT 1.875 1.09 2.015 1.44 ;
 RECT 1.78 1.44 2.025 1.59 ;
 RECT 2.575 1.75 2.715 1.805 ;
 RECT 2.575 1.53 2.715 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.24 1.115 2.66 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.58 1.27 20.925 1.545 ;
 RECT 20.715 0.93 21.04 1.07 ;
 RECT 21.7 0.93 22.025 1.07 ;
 RECT 20.785 1.71 21.93 1.85 ;
 RECT 20.785 1.85 20.925 1.895 ;
 RECT 20.785 1.545 20.925 1.71 ;
 RECT 20.785 1.07 20.925 1.27 ;
 RECT 20.785 0.915 20.925 0.93 ;
 RECT 21.79 0.925 21.93 0.93 ;
 RECT 21.79 1.85 21.93 1.895 ;
 RECT 21.79 1.07 21.93 1.71 ;
 END
 ANTENNADIFFAREA 0.805 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.195 1.17 22.435 1.41 ;
 RECT 22.295 1.775 24.5 1.915 ;
 RECT 22.295 0.645 22.435 1.17 ;
 RECT 23.355 1.915 23.495 1.92 ;
 RECT 23.355 0.66 23.495 1.775 ;
 RECT 22.295 1.915 22.435 1.925 ;
 RECT 22.295 1.41 22.435 1.775 ;
 END
 ANTENNADIFFAREA 1.186 ;
 END Q

 OBS
 LAYER PO ;
 RECT 17.07 0.835 17.17 2.39 ;
 RECT 27.805 0.215 27.905 0.995 ;
 RECT 27.805 0.995 28.045 1.205 ;
 RECT 27.805 1.205 27.905 2 ;
 RECT 30.2 0.375 30.3 0.99 ;
 RECT 30.2 0.99 30.45 1.2 ;
 RECT 30.2 1.2 30.3 2.27 ;
 RECT 30.2 2.27 30.485 2.48 ;
 RECT 13.48 0.655 13.58 2.305 ;
 RECT 13.785 2.3 14.015 2.305 ;
 RECT 13.785 2.405 14.015 2.51 ;
 RECT 13.48 2.305 14.015 2.405 ;
 RECT 27.025 0.21 27.125 0.755 ;
 RECT 27.025 0.855 27.125 2.2 ;
 RECT 29.89 1.125 29.99 2.2 ;
 RECT 26.06 0.755 27.595 0.84 ;
 RECT 26.06 0.84 27.59 0.855 ;
 RECT 27.495 0.215 27.595 0.755 ;
 RECT 26.06 0.595 26.29 0.755 ;
 RECT 27.025 2.2 29.99 2.3 ;
 RECT 12.19 1.28 12.445 1.45 ;
 RECT 12.19 1.45 12.29 1.655 ;
 RECT 12.19 0.655 12.29 1.18 ;
 RECT 12.19 1.655 13.15 1.755 ;
 RECT 13.05 1.755 13.15 2.355 ;
 RECT 11.275 0.66 11.375 1.18 ;
 RECT 12.19 1.755 12.29 2.51 ;
 RECT 11.275 1.24 12.445 1.28 ;
 RECT 11.275 1.18 12.29 1.24 ;
 RECT 28.715 0.38 28.815 0.96 ;
 RECT 28.715 1.06 28.815 1.14 ;
 RECT 28.295 0.935 28.525 0.96 ;
 RECT 28.295 0.96 28.815 1.06 ;
 RECT 28.295 1.06 28.525 1.145 ;
 RECT 28.715 1.14 28.985 1.24 ;
 RECT 28.885 1.24 28.985 1.84 ;
 RECT 29.08 0.22 29.31 0.28 ;
 RECT 29.08 0.38 29.31 0.43 ;
 RECT 28.715 0.28 29.31 0.38 ;
 RECT 11.265 1.575 11.365 2.485 ;
 RECT 11.775 1.575 12.005 1.685 ;
 RECT 11.265 1.475 12.005 1.575 ;
 RECT 30.9 0.195 31 2.665 ;
 RECT 29.89 0.095 31 0.195 ;
 RECT 26.265 1.245 26.365 2.665 ;
 RECT 29.89 0.195 29.99 0.945 ;
 RECT 26.265 1.2 26.55 1.245 ;
 RECT 26.32 1.035 26.55 1.1 ;
 RECT 26.265 2.665 31 2.765 ;
 RECT 26.265 1.1 26.595 1.2 ;
 RECT 15.49 0.795 15.655 0.925 ;
 RECT 14.81 0.885 15.04 0.925 ;
 RECT 14.81 1.025 15.04 1.095 ;
 RECT 14.81 0.925 15.655 1.025 ;
 RECT 15.49 0.585 15.72 0.795 ;
 RECT 2.525 1.55 2.765 1.78 ;
 RECT 2.665 1.78 2.765 2.695 ;
 RECT 1.055 1.435 1.625 1.71 ;
 RECT 1.055 0.515 1.155 1.435 ;
 RECT 1.055 1.71 1.155 2.645 ;
 RECT 1.525 0.515 1.625 1.435 ;
 RECT 1.525 1.71 1.625 2.695 ;
 RECT 2.245 1.37 2.345 1.605 ;
 RECT 2.475 0.515 2.575 1.14 ;
 RECT 2.195 1.705 2.295 2.695 ;
 RECT 2.195 1.605 2.345 1.705 ;
 RECT 2.245 1.14 2.575 1.37 ;
 RECT 1.86 0.515 1.96 1.105 ;
 RECT 1.82 1.105 2.065 1.345 ;
 RECT 4.41 0.52 4.51 2.465 ;
 RECT 4.17 0.27 4.51 0.52 ;
 RECT 7.04 1.33 7.18 1.475 ;
 RECT 7.04 1.71 7.14 2.475 ;
 RECT 7.08 0.65 7.18 1.33 ;
 RECT 7.04 1.475 7.27 1.71 ;
 RECT 6.59 0.705 6.69 1.165 ;
 RECT 6.15 1.27 6.25 1.445 ;
 RECT 6.59 0.47 6.875 0.705 ;
 RECT 6.15 1.17 6.69 1.265 ;
 RECT 6.15 1.265 6.525 1.27 ;
 RECT 6.38 1.165 6.69 1.17 ;
 RECT 6.005 1.445 6.25 1.69 ;
 RECT 7.48 0.715 7.58 1.61 ;
 RECT 7.515 1.71 7.615 2.48 ;
 RECT 7.48 1.61 7.615 1.71 ;
 RECT 7.36 0.485 7.6 0.715 ;
 RECT 13.085 0.655 13.185 1.24 ;
 RECT 12.955 1.24 13.185 1.475 ;
 RECT 4.885 0.49 4.985 1.495 ;
 RECT 4.69 1.495 4.985 1.745 ;
 RECT 4.885 1.745 4.985 2.37 ;
 RECT 8.705 0.59 9.03 0.74 ;
 RECT 8.93 0.74 9.03 2.45 ;
 RECT 8.755 2.45 9.03 2.66 ;
 RECT 8.705 0.53 8.935 0.59 ;
 RECT 2.8 0.245 3.065 0.455 ;
 RECT 2.965 0.455 3.065 2.695 ;
 RECT 3.435 0.295 3.535 1.115 ;
 RECT 3.245 1.115 3.535 1.325 ;
 RECT 3.435 1.325 3.535 2.765 ;
 RECT 19.51 0.77 19.61 2.155 ;
 RECT 19.51 0.55 19.61 0.56 ;
 RECT 19.51 0.56 19.765 0.77 ;
 RECT 21.05 0.375 21.15 1.41 ;
 RECT 20.145 0.43 20.245 1.245 ;
 RECT 21.54 0.445 21.64 1.41 ;
 RECT 21.54 1.51 21.64 2.645 ;
 RECT 21.05 1.51 21.15 2.57 ;
 RECT 20.145 0.22 20.375 0.275 ;
 RECT 20.145 0.375 20.375 0.43 ;
 RECT 20.145 0.275 21.15 0.375 ;
 RECT 21.05 1.41 21.64 1.51 ;
 RECT 20.095 1.245 20.325 1.455 ;
 RECT 8.3 2.445 8.56 2.655 ;
 RECT 8.46 1.79 8.56 2.445 ;
 RECT 18.57 1.445 18.67 2.035 ;
 RECT 18.555 2.035 18.785 2.245 ;
 RECT 19.04 0.55 19.14 2.69 ;
 RECT 9.97 1.58 10.07 1.735 ;
 RECT 9.71 1.01 9.81 1.48 ;
 RECT 9.97 1.945 10.07 2.69 ;
 RECT 9.97 1.735 10.205 1.945 ;
 RECT 9.71 1.48 10.07 1.58 ;
 RECT 9.97 2.69 19.14 2.79 ;
 RECT 9.41 0.98 9.51 1.615 ;
 RECT 9.27 1.615 9.51 1.825 ;
 RECT 9.41 1.825 9.51 2.605 ;
 RECT 22.555 1.295 24.18 1.395 ;
 RECT 22.555 1.26 22.805 1.295 ;
 RECT 22.555 0.375 22.655 1.26 ;
 RECT 23.135 0.375 23.235 1.295 ;
 RECT 24.08 1.395 24.18 2.685 ;
 RECT 23.61 1.395 23.71 2.69 ;
 RECT 22.555 1.47 22.655 2.69 ;
 RECT 22.555 1.395 22.805 1.47 ;
 RECT 23.135 1.395 23.235 2.715 ;
 RECT 25.28 0.22 25.51 0.275 ;
 RECT 25.28 0.375 25.51 0.43 ;
 RECT 23.135 0.275 25.51 0.375 ;
 RECT 17.54 0.73 17.64 1.39 ;
 RECT 17.405 1.39 17.64 1.6 ;
 RECT 17.54 1.6 17.64 2.39 ;
 RECT 5.725 0.285 5.825 1.52 ;
 RECT 5.225 1.52 5.825 1.62 ;
 RECT 5.725 0.185 14.615 0.195 ;
 RECT 7.78 0.095 14.615 0.185 ;
 RECT 5.725 0.195 7.88 0.285 ;
 RECT 14.515 0.195 14.615 1.29 ;
 RECT 15.41 1.39 15.605 1.405 ;
 RECT 6.545 1.565 6.645 2.675 ;
 RECT 5.66 1.62 5.76 2.675 ;
 RECT 5.225 1.44 5.47 1.52 ;
 RECT 5.225 1.62 5.47 1.69 ;
 RECT 7.78 0.285 7.88 1.24 ;
 RECT 14.515 1.29 15.605 1.39 ;
 RECT 5.66 2.675 6.645 2.775 ;
 RECT 15.41 1.405 15.64 1.615 ;
 RECT 27.5 1.245 27.6 2.02 ;
 RECT 27.37 1.035 27.6 1.245 ;
 RECT 15.905 0.105 18.73 0.205 ;
 RECT 15.905 0.205 16.005 1.91 ;
 RECT 18.63 0.205 18.73 1.265 ;
 RECT 15.085 1.71 15.185 1.91 ;
 RECT 14 1.61 15.185 1.71 ;
 RECT 14 0.475 14.1 1.61 ;
 RECT 14.55 1.71 14.65 2.425 ;
 RECT 10.665 0.475 10.765 0.895 ;
 RECT 15.085 1.91 16.005 2.01 ;
 RECT 10.665 0.375 14.1 0.475 ;
 RECT 10.54 0.895 10.77 1.105 ;
 RECT 16.215 0.455 18.145 0.535 ;
 RECT 17.915 0.535 18.145 0.6 ;
 RECT 17.915 0.39 18.145 0.435 ;
 RECT 16.295 0.435 18.145 0.455 ;
 RECT 16.215 0.535 16.445 0.665 ;
 RECT 17.07 0.535 17.3 0.835 ;
 LAYER CO ;
 RECT 26.11 0.635 26.24 0.765 ;
 RECT 12.265 1.28 12.395 1.41 ;
 RECT 29.13 0.26 29.26 0.39 ;
 RECT 11.825 1.515 11.955 1.645 ;
 RECT 26.37 1.075 26.5 1.205 ;
 RECT 14.86 0.925 14.99 1.055 ;
 RECT 0.805 0.735 0.935 0.865 ;
 RECT 3.185 2.31 3.315 2.44 ;
 RECT 1.275 2.015 1.405 2.145 ;
 RECT 1.88 1.155 2.01 1.285 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 2.58 1.6 2.71 1.73 ;
 RECT 3.655 2.01 3.785 2.14 ;
 RECT 3.655 0.735 3.785 0.865 ;
 RECT 2.415 2.075 2.545 2.205 ;
 RECT 1.275 2.275 1.405 2.405 ;
 RECT 3.185 0.545 3.315 0.675 ;
 RECT 3.655 1.75 3.785 1.88 ;
 RECT 0.805 2.015 0.935 2.145 ;
 RECT 2.22 0.735 2.35 0.865 ;
 RECT 2.4 1.19 2.53 1.32 ;
 RECT 28.965 0.595 29.095 0.725 ;
 RECT 6.695 0.525 6.825 0.655 ;
 RECT 7.74 1.825 7.87 1.955 ;
 RECT 29.475 1.49 29.605 1.62 ;
 RECT 6.34 0.88 6.47 1.01 ;
 RECT 14.77 1.87 14.9 2 ;
 RECT 8.21 2.11 8.34 2.24 ;
 RECT 8.025 0.32 8.155 0.45 ;
 RECT 27.245 0.135 27.375 0.265 ;
 RECT 5.285 1.495 5.415 1.625 ;
 RECT 5.235 0.745 5.365 0.875 ;
 RECT 5.105 1.995 5.235 2.125 ;
 RECT 11.94 1.995 12.07 2.125 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 11.495 2.07 11.625 2.2 ;
 RECT 14.265 0.595 14.395 0.725 ;
 RECT 6.06 1.49 6.19 1.62 ;
 RECT 13.005 1.28 13.135 1.41 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 23.83 2.64 23.96 2.77 ;
 RECT 23.36 1.72 23.49 1.85 ;
 RECT 23.36 0.73 23.49 0.86 ;
 RECT 20.79 0.935 20.92 1.065 ;
 RECT 21.28 0.315 21.41 0.445 ;
 RECT 22.3 1.735 22.43 1.865 ;
 RECT 22.775 2.635 22.905 2.765 ;
 RECT 21.795 1.715 21.925 1.845 ;
 RECT 21.27 2.635 21.4 2.765 ;
 RECT 24.3 1.78 24.43 1.91 ;
 RECT 22.3 0.72 22.43 0.85 ;
 RECT 9.7 2.165 9.83 2.295 ;
 RECT 5.215 0.145 5.345 0.275 ;
 RECT 14.265 1.9 14.395 2.03 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 5.37 2.345 5.5 2.475 ;
 RECT 28.025 0.435 28.155 0.565 ;
 RECT 9.97 1.23 10.1 1.36 ;
 RECT 18.79 1.705 18.92 1.835 ;
 RECT 9.16 2.195 9.29 2.325 ;
 RECT 6.81 0.88 6.94 1.01 ;
 RECT 16.82 1.835 16.95 1.965 ;
 RECT 16.69 0.765 16.82 0.895 ;
 RECT 4.63 0.74 4.76 0.87 ;
 RECT 29.64 0.12 29.77 0.25 ;
 RECT 7.415 0.53 7.545 0.66 ;
 RECT 15.665 2.38 15.795 2.51 ;
 RECT 11.94 0.885 12.07 1.015 ;
 RECT 26.775 1.425 26.905 1.555 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 19.855 0.92 19.985 1.05 ;
 RECT 27.245 1.475 27.375 1.605 ;
 RECT 13.74 0.875 13.87 1.005 ;
 RECT 5.945 0.79 6.075 0.92 ;
 RECT 17.76 1.835 17.89 1.965 ;
 RECT 6.79 2.07 6.92 2.2 ;
 RECT 31.2 1.475 31.33 1.605 ;
 RECT 4.16 0.74 4.29 0.87 ;
 RECT 5.88 1.825 6.01 1.955 ;
 RECT 13.74 1.945 13.87 2.075 ;
 RECT 4.63 2.05 4.76 2.18 ;
 RECT 26.525 0.505 26.655 0.635 ;
 RECT 11.015 2.015 11.145 2.145 ;
 RECT 28.46 0.12 28.59 0.25 ;
 RECT 28.025 1.485 28.155 1.615 ;
 RECT 30.42 1.465 30.55 1.595 ;
 RECT 19.26 1.705 19.39 1.835 ;
 RECT 30.42 0.595 30.55 0.725 ;
 RECT 7.09 1.525 7.22 1.655 ;
 RECT 12.64 2.225 12.77 2.355 ;
 RECT 4.16 2.115 4.29 2.245 ;
 RECT 19.735 1.705 19.865 1.835 ;
 RECT 29.105 1.405 29.235 1.535 ;
 RECT 11.02 0.905 11.15 1.035 ;
 RECT 4.23 0.325 4.36 0.455 ;
 RECT 9.16 0.315 9.29 0.445 ;
 RECT 11.495 0.905 11.625 1.035 ;
 RECT 14.77 0.595 14.9 0.725 ;
 RECT 12.83 0.595 12.96 0.725 ;
 RECT 28.63 1.445 28.76 1.575 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 17.795 1.035 17.925 1.165 ;
 RECT 18.38 0.91 18.51 1.04 ;
 RECT 10.19 2.43 10.32 2.56 ;
 RECT 8.68 2.135 8.81 2.265 ;
 RECT 6.295 2.105 6.425 2.235 ;
 RECT 7.26 2.11 7.39 2.24 ;
 RECT 8.805 2.49 8.935 2.62 ;
 RECT 8.755 0.57 8.885 0.7 ;
 RECT 2.85 0.285 2.98 0.415 ;
 RECT 3.295 1.155 3.425 1.285 ;
 RECT 22.625 1.3 22.755 1.43 ;
 RECT 20.145 1.285 20.275 1.415 ;
 RECT 17.965 0.43 18.095 0.56 ;
 RECT 19.585 0.6 19.715 0.73 ;
 RECT 20.195 0.26 20.325 0.39 ;
 RECT 8.35 2.485 8.48 2.615 ;
 RECT 18.605 2.075 18.735 2.205 ;
 RECT 10.025 1.775 10.155 1.905 ;
 RECT 9.32 1.655 9.45 1.785 ;
 RECT 25.33 0.26 25.46 0.39 ;
 RECT 30.27 1.03 30.4 1.16 ;
 RECT 16.265 0.495 16.395 0.625 ;
 RECT 17.455 1.43 17.585 1.56 ;
 RECT 15.54 0.625 15.67 0.755 ;
 RECT 15.46 1.445 15.59 1.575 ;
 RECT 27.42 1.075 27.55 1.205 ;
 RECT 10.59 0.935 10.72 1.065 ;
 RECT 28.345 0.975 28.475 1.105 ;
 RECT 17.12 0.665 17.25 0.795 ;
 RECT 27.865 1.035 27.995 1.165 ;
 RECT 30.305 2.31 30.435 2.44 ;
 RECT 13.835 2.34 13.965 2.47 ;
 RECT 4.75 1.55 4.88 1.68 ;
 RECT 20.79 1.715 20.92 1.845 ;
 RECT 22.86 0.72 22.99 0.85 ;
 RECT 21.795 0.935 21.925 1.065 ;
 RECT 1.275 0.735 1.405 0.865 ;
 RECT 1.28 1.51 1.41 1.64 ;
 LAYER M1 ;
 RECT 28.02 1.485 28.16 1.76 ;
 RECT 28.34 0.73 28.48 0.935 ;
 RECT 28.02 0.355 28.16 0.59 ;
 RECT 28.02 1.345 28.48 1.485 ;
 RECT 28.295 0.935 28.525 1.145 ;
 RECT 28.02 0.59 28.48 0.73 ;
 RECT 25.28 0.36 25.51 0.43 ;
 RECT 26.875 0.36 27.015 0.565 ;
 RECT 25.28 0.22 27.015 0.36 ;
 RECT 27.615 0.705 27.755 0.75 ;
 RECT 27.74 0.995 28.045 1.205 ;
 RECT 27.74 0.89 27.88 0.995 ;
 RECT 27.615 0.75 27.88 0.89 ;
 RECT 26.875 0.565 27.755 0.705 ;
 RECT 14.765 0.525 14.905 0.885 ;
 RECT 14.765 1.095 14.905 2.065 ;
 RECT 14.765 0.885 15.04 1.095 ;
 RECT 18.81 0.775 18.95 1.405 ;
 RECT 19.535 0.56 19.765 0.635 ;
 RECT 17.79 1.405 18.95 1.545 ;
 RECT 17.79 1.545 17.93 1.83 ;
 RECT 16.745 1.83 17.995 1.97 ;
 RECT 17.79 1.17 17.93 1.405 ;
 RECT 17.72 1.03 18 1.17 ;
 RECT 21.685 0.38 21.825 0.635 ;
 RECT 18.81 0.635 21.825 0.775 ;
 RECT 22.575 0.38 22.715 1.26 ;
 RECT 21.685 0.24 22.715 0.38 ;
 RECT 22.575 1.26 22.805 1.47 ;
 RECT 20.145 0.22 20.375 0.28 ;
 RECT 20.145 0.42 20.375 0.43 ;
 RECT 17.915 0.28 20.375 0.42 ;
 RECT 17.915 0.42 18.145 0.6 ;
 RECT 15.49 0.585 16.445 0.63 ;
 RECT 16.215 0.63 16.445 0.665 ;
 RECT 16.215 0.455 16.445 0.49 ;
 RECT 15.515 0.49 16.445 0.585 ;
 RECT 15.49 0.63 15.72 0.795 ;
 RECT 17.07 0.57 17.3 0.95 ;
 RECT 11.49 1.04 11.63 2.34 ;
 RECT 11.49 0.895 11.63 0.9 ;
 RECT 11.42 0.9 11.695 1.04 ;
 RECT 12.285 2.055 12.425 2.34 ;
 RECT 11.49 2.34 12.425 2.48 ;
 RECT 13.42 1.66 13.56 1.915 ;
 RECT 12.285 1.915 13.56 2.055 ;
 RECT 14.26 0.525 14.4 1.52 ;
 RECT 14.26 1.66 14.4 2.11 ;
 RECT 13.735 0.765 13.875 1.52 ;
 RECT 13.735 1.66 13.875 2.145 ;
 RECT 13.42 1.52 14.4 1.66 ;
 RECT 5.94 1.67 6.08 1.82 ;
 RECT 5.94 1.96 6.08 2.51 ;
 RECT 8.3 2.445 8.53 2.51 ;
 RECT 8.3 2.65 8.53 2.655 ;
 RECT 5.94 0.5 6.08 1.44 ;
 RECT 5.94 1.44 6.195 1.67 ;
 RECT 5.81 1.82 6.08 1.96 ;
 RECT 5.94 2.51 8.53 2.65 ;
 RECT 7.085 0.895 10.77 1.035 ;
 RECT 10.54 1.035 10.77 1.105 ;
 RECT 7.085 0.66 7.225 0.895 ;
 RECT 6.625 0.52 7.225 0.66 ;
 RECT 5.185 0.88 5.325 1.475 ;
 RECT 5.145 1.63 5.285 1.99 ;
 RECT 5.145 1.475 5.49 1.63 ;
 RECT 5.035 1.99 5.285 2.13 ;
 RECT 5.185 0.74 5.505 0.88 ;
 RECT 7.365 0.71 11.46 0.745 ;
 RECT 8.705 0.53 8.935 0.605 ;
 RECT 7.365 0.485 7.68 0.605 ;
 RECT 17.06 1.23 17.2 1.42 ;
 RECT 15.21 1.09 17.2 1.23 ;
 RECT 15.21 0.385 15.35 1.09 ;
 RECT 13.2 0.385 13.34 0.875 ;
 RECT 13.2 0.255 15.35 0.385 ;
 RECT 13.2 0.245 15.345 0.255 ;
 RECT 12.48 0.875 13.34 1.015 ;
 RECT 12.48 0.71 12.62 0.875 ;
 RECT 7.365 0.605 12.62 0.71 ;
 RECT 11.21 0.57 12.62 0.605 ;
 RECT 17.405 1.39 17.635 1.42 ;
 RECT 17.06 1.42 17.635 1.56 ;
 RECT 17.405 1.56 17.635 1.6 ;
 RECT 2.87 0.87 3.01 1.15 ;
 RECT 2.87 1.29 3.01 2.07 ;
 RECT 2.36 2.07 3.01 2.21 ;
 RECT 2.165 0.73 3.01 0.87 ;
 RECT 3.245 1.115 3.475 1.15 ;
 RECT 3.245 1.29 3.475 1.325 ;
 RECT 2.87 1.15 3.475 1.29 ;
 RECT 3.935 1.335 4.075 2.11 ;
 RECT 3.935 2.25 4.075 2.255 ;
 RECT 3.935 0.875 4.075 1.195 ;
 RECT 3.935 2.11 4.36 2.25 ;
 RECT 3.935 0.735 4.36 0.875 ;
 RECT 3.935 1.195 5.045 1.335 ;
 RECT 4.905 0.6 5.045 1.195 ;
 RECT 6.335 0.36 6.475 2.035 ;
 RECT 5.65 0.22 6.475 0.36 ;
 RECT 5.65 0.36 5.79 0.46 ;
 RECT 6.29 2.17 6.43 2.305 ;
 RECT 6.29 2.035 6.475 2.17 ;
 RECT 4.905 0.46 5.79 0.6 ;
 RECT 3.65 0.46 3.79 2.21 ;
 RECT 4.12 0.22 4.485 0.32 ;
 RECT 4.12 0.46 4.485 0.525 ;
 RECT 3.65 0.32 4.485 0.46 ;
 RECT 0.8 0.68 0.94 1.155 ;
 RECT 0.8 1.295 0.94 2.23 ;
 RECT 1.585 0.385 1.725 1.155 ;
 RECT 0.8 1.155 1.725 1.295 ;
 RECT 2.8 0.385 3.03 0.455 ;
 RECT 1.585 0.245 3.03 0.385 ;
 RECT 16.18 1.895 16.32 2.39 ;
 RECT 20.325 2.205 20.465 2.39 ;
 RECT 16.18 2.39 20.465 2.53 ;
 RECT 15.055 1.755 16.32 1.895 ;
 RECT 15.055 1.895 15.195 2.34 ;
 RECT 13.785 2.3 14.015 2.34 ;
 RECT 13.785 2.48 14.015 2.51 ;
 RECT 13.785 2.34 15.195 2.48 ;
 RECT 20.325 2.065 26.055 2.205 ;
 RECT 25.915 2.205 26.055 2.52 ;
 RECT 30.255 2.48 30.395 2.52 ;
 RECT 25.915 2.52 30.395 2.66 ;
 RECT 30.255 2.27 30.485 2.48 ;
 RECT 19.815 1.055 19.955 1.245 ;
 RECT 19.255 1.385 19.395 1.625 ;
 RECT 20.095 1.385 20.325 1.455 ;
 RECT 19.255 1.245 20.325 1.385 ;
 RECT 19.785 0.915 20.085 1.055 ;
 RECT 19.225 1.625 19.48 1.92 ;
 RECT 19.62 1.7 19.915 1.84 ;
 RECT 19.62 1.84 19.76 2.075 ;
 RECT 18.925 1.84 19.065 2.075 ;
 RECT 18.73 1.7 19.065 1.84 ;
 RECT 18.925 2.075 19.76 2.215 ;
 RECT 16.46 1.56 16.6 2.11 ;
 RECT 16.46 2.11 18.785 2.245 ;
 RECT 16.46 2.245 18.78 2.25 ;
 RECT 18.555 2.035 18.785 2.11 ;
 RECT 15.41 1.405 15.64 1.42 ;
 RECT 15.41 1.56 15.64 1.615 ;
 RECT 15.41 1.42 16.6 1.56 ;
 RECT 11.935 1.02 12.075 1.475 ;
 RECT 11.775 1.475 12.075 1.635 ;
 RECT 11.935 1.775 12.075 2.18 ;
 RECT 11.86 0.88 12.135 1.02 ;
 RECT 11.935 1.685 13.14 1.775 ;
 RECT 13 1.415 13.14 1.635 ;
 RECT 11.775 1.635 13.14 1.685 ;
 RECT 12.95 1.275 13.205 1.415 ;
 RECT 7.19 2.105 8.41 2.245 ;
 RECT 9.695 1.365 9.835 2.36 ;
 RECT 7.75 1.365 7.89 1.5 ;
 RECT 6.92 1.64 7.425 1.675 ;
 RECT 6.92 1.5 7.89 1.64 ;
 RECT 11.01 1.04 11.15 1.25 ;
 RECT 11.01 1.39 11.15 2.215 ;
 RECT 11.01 0.885 11.15 0.9 ;
 RECT 7.75 1.25 11.15 1.365 ;
 RECT 7.75 1.225 10.4 1.25 ;
 RECT 10.26 1.365 11.15 1.39 ;
 RECT 10.945 0.9 11.22 1.04 ;
 RECT 6.63 1.82 8.21 1.96 ;
 RECT 8.07 1.79 8.21 1.82 ;
 RECT 6.63 1.22 6.945 1.36 ;
 RECT 6.805 0.805 6.945 1.22 ;
 RECT 6.715 1.96 6.995 2.215 ;
 RECT 6.63 1.36 6.77 1.82 ;
 RECT 9.27 1.615 9.5 1.65 ;
 RECT 9.27 1.79 9.5 1.825 ;
 RECT 8.07 1.65 9.505 1.79 ;
 RECT 28.96 0.73 29.1 1.04 ;
 RECT 29.1 1.18 29.24 1.605 ;
 RECT 28.895 0.59 29.17 0.73 ;
 RECT 30.22 0.99 30.45 1.04 ;
 RECT 28.96 1.04 30.45 1.18 ;
 RECT 30.22 1.18 30.45 1.2 ;
 RECT 29.08 0.29 29.45 0.43 ;
 RECT 29.31 0.43 29.45 0.71 ;
 RECT 29.08 0.22 29.31 0.29 ;
 RECT 30.73 0.85 30.87 1.385 ;
 RECT 30.415 1.525 30.555 1.73 ;
 RECT 29.31 0.71 30.87 0.85 ;
 RECT 30.415 0.51 30.555 0.71 ;
 RECT 30.415 1.385 30.87 1.525 ;
 RECT 26.32 1.225 26.55 1.245 ;
 RECT 26.32 1.195 26.91 1.225 ;
 RECT 26.46 1.015 26.77 1.035 ;
 RECT 26.32 1.035 26.77 1.055 ;
 RECT 26.595 0.64 26.735 1.015 ;
 RECT 26.77 1.225 26.91 1.75 ;
 RECT 26.475 0.5 26.735 0.64 ;
 RECT 27.37 1.035 27.6 1.055 ;
 RECT 27.37 1.195 27.6 1.245 ;
 RECT 26.32 1.055 27.6 1.195 ;
 RECT 28.34 1.145 28.48 1.345 ;
 END
END RSDFFNSRASX2

MACRO RSDFFNSRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.52 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.08 1.16 18.445 1.4 ;
 RECT 18.305 0.695 18.445 1.16 ;
 RECT 19.365 1.905 19.505 1.91 ;
 RECT 18.305 1.765 19.505 1.905 ;
 RECT 19.365 0.71 19.505 1.765 ;
 RECT 18.305 1.4 18.445 1.765 ;
 END
 ANTENNADIFFAREA 0.729 ;
 END Q

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.79 1.475 5.12 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.35 1.16 10.68 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 16.78 1.7 17.925 1.75 ;
 RECT 16.565 1.75 17.925 1.84 ;
 RECT 16.565 1.84 16.92 1.99 ;
 RECT 17.785 0.915 17.925 1.7 ;
 RECT 16.78 0.905 16.92 1.7 ;
 RECT 17.785 1.84 17.925 1.92 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 27.52 2.96 ;
 RECT 1.36 2.005 1.5 2.8 ;
 RECT 5.415 2.34 5.665 2.8 ;
 RECT 10.77 2.375 10.91 2.8 ;
 RECT 4.74 1.98 4.88 2.8 ;
 RECT 3.27 2.03 3.41 2.8 ;
 RECT 15.205 2.57 15.345 2.8 ;
 RECT 14.36 2.57 14.5 2.8 ;
 RECT 8.67 2.07 8.81 2.8 ;
 RECT 0.385 1.74 0.525 2.8 ;
 RECT 18.78 2.57 18.92 2.8 ;
 RECT 17.265 2.57 17.405 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 27.52 0.08 ;
 RECT 17.215 0.28 17.48 0.44 ;
 RECT 3.27 0.08 3.41 0.78 ;
 RECT 8.085 0.08 8.32 0.595 ;
 RECT 4.74 0.08 4.88 1.055 ;
 RECT 24.345 0.08 24.585 0.31 ;
 RECT 21.995 0.08 22.135 0.31 ;
 RECT 15.21 0.08 15.35 0.525 ;
 RECT 1.36 0.08 1.5 0.97 ;
 RECT 5.485 0.08 5.625 0.39 ;
 RECT 18.865 0.08 19.005 0.965 ;
 RECT 23.21 0.08 23.35 0.325 ;
 RECT 0.35 0.08 0.49 0.775 ;
 RECT 10.96 0.08 11.1 0.815 ;
 RECT 14.135 0.08 14.275 1.155 ;
 RECT 17.27 0.08 17.41 0.28 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.33 1.155 2.75 1.415 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.18 1.475 1.705 1.75 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.965 1.13 2.105 1.48 ;
 RECT 1.87 1.63 2.815 1.79 ;
 RECT 1.87 1.48 2.115 1.63 ;
 RECT 2.665 1.79 2.805 1.845 ;
 RECT 2.665 1.57 2.805 1.63 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 25.905 1.41 26.245 1.775 ;
 RECT 24.225 1.965 26.09 2.105 ;
 RECT 21.995 2.195 24.365 2.335 ;
 RECT 24.225 1.41 24.365 1.965 ;
 RECT 25.95 1.775 26.09 1.965 ;
 RECT 21.995 1.365 22.135 2.195 ;
 RECT 23.38 1.345 23.52 2.195 ;
 RECT 24.225 2.105 24.365 2.195 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.565 0.57 21.045 0.78 ;
 RECT 20.565 0.78 20.935 0.865 ;
 RECT 20.565 0.565 20.935 0.57 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 OBS
 LAYER PO ;
 RECT 16.425 0.84 16.525 1.3 ;
 RECT 15.895 1.46 15.995 2.56 ;
 RECT 15.735 1.4 15.995 1.46 ;
 RECT 15.735 1.3 16.525 1.4 ;
 RECT 16.41 0.63 16.64 0.84 ;
 RECT 22.12 1.01 22.355 1.22 ;
 RECT 22.255 1.22 22.355 1.995 ;
 RECT 23.47 0.355 23.57 0.985 ;
 RECT 23.47 0.255 24.205 0.355 ;
 RECT 23.975 0.355 24.205 0.465 ;
 RECT 23.64 1.215 23.74 1.815 ;
 RECT 23.08 1.115 23.74 1.215 ;
 RECT 23.08 0.985 23.57 1.115 ;
 RECT 18.55 1.285 19.245 1.385 ;
 RECT 18.55 1.385 18.76 1.435 ;
 RECT 19.145 0.38 19.245 1.285 ;
 RECT 18.55 1.2 18.76 1.285 ;
 RECT 18.565 0.47 18.665 1.2 ;
 RECT 18.565 1.435 18.665 2.645 ;
 RECT 19.145 1.385 19.245 2.645 ;
 RECT 19.815 0.205 20.045 0.28 ;
 RECT 19.815 0.38 20.045 0.435 ;
 RECT 19.145 0.28 20.045 0.38 ;
 RECT 11.615 2.69 13.265 2.695 ;
 RECT 13.09 2.54 13.265 2.69 ;
 RECT 12.405 2.695 13.265 2.79 ;
 RECT 11.615 0.655 11.715 2.595 ;
 RECT 11.615 2.595 12.505 2.69 ;
 RECT 13.09 2.33 13.32 2.54 ;
 RECT 4.285 0.27 4.625 0.52 ;
 RECT 4.525 0.52 4.625 2.465 ;
 RECT 11.22 0.655 11.32 1.24 ;
 RECT 11.09 1.24 11.32 1.475 ;
 RECT 8.76 1.61 9.025 1.82 ;
 RECT 8.925 1.82 9.025 2.49 ;
 RECT 8.555 0.66 8.655 1.51 ;
 RECT 8.555 1.51 9.025 1.61 ;
 RECT 21.02 1.175 21.305 1.305 ;
 RECT 21.02 1.305 21.12 2.64 ;
 RECT 24.645 0.19 24.745 0.94 ;
 RECT 24.645 0.09 25.755 0.19 ;
 RECT 25.655 0.19 25.755 2.64 ;
 RECT 21.02 1.075 21.35 1.175 ;
 RECT 21.02 2.64 25.755 2.74 ;
 RECT 17.045 0.39 17.145 1.4 ;
 RECT 16.04 0.225 16.27 0.29 ;
 RECT 16.04 0.39 16.27 0.435 ;
 RECT 16.04 0.29 17.145 0.39 ;
 RECT 17.045 1.5 17.145 2.26 ;
 RECT 17.535 0.505 17.635 1.4 ;
 RECT 17.535 1.5 17.635 2.26 ;
 RECT 17.045 1.4 17.635 1.5 ;
 RECT 5 0.57 5.1 1.495 ;
 RECT 4.805 1.495 5.1 1.745 ;
 RECT 5 1.745 5.1 2.37 ;
 RECT 7.195 1.475 7.505 1.71 ;
 RECT 7.195 0.65 7.295 1.475 ;
 RECT 7.195 1.71 7.295 2.475 ;
 RECT 5.775 1.62 5.875 2.375 ;
 RECT 5.84 0.185 12.75 0.19 ;
 RECT 12.65 0.19 12.75 1.29 ;
 RECT 5.84 0.19 7.995 0.285 ;
 RECT 5.84 0.285 5.94 1.52 ;
 RECT 6.66 1.565 6.76 2.375 ;
 RECT 13.44 1.285 13.67 1.29 ;
 RECT 13.44 1.39 13.67 1.615 ;
 RECT 12.65 1.29 13.67 1.39 ;
 RECT 5.34 1.44 5.585 1.52 ;
 RECT 5.34 1.62 5.585 1.69 ;
 RECT 5.34 1.52 5.94 1.62 ;
 RECT 7.895 0.09 12.75 0.185 ;
 RECT 7.895 0.285 7.995 1.24 ;
 RECT 5.775 2.375 6.76 2.475 ;
 RECT 2.755 1.82 2.855 2.735 ;
 RECT 2.615 1.59 2.855 1.82 ;
 RECT 1.95 0.555 2.05 1.145 ;
 RECT 1.91 1.145 2.155 1.385 ;
 RECT 3.525 0.335 3.625 1.155 ;
 RECT 3.525 1.365 3.625 2.745 ;
 RECT 3.335 1.155 3.625 1.365 ;
 RECT 1.145 1.475 1.715 1.75 ;
 RECT 1.145 0.555 1.245 1.475 ;
 RECT 1.145 1.75 1.245 2.685 ;
 RECT 1.615 0.555 1.715 1.475 ;
 RECT 1.615 1.75 1.715 2.735 ;
 RECT 2.335 1.41 2.435 1.645 ;
 RECT 2.565 0.555 2.665 1.18 ;
 RECT 2.285 1.745 2.385 2.735 ;
 RECT 2.285 1.645 2.435 1.745 ;
 RECT 2.335 1.18 2.665 1.41 ;
 RECT 3.055 0.405 3.155 2.735 ;
 RECT 2.85 0.175 3.155 0.405 ;
 RECT 8.455 1.79 8.555 2.465 ;
 RECT 8.24 2.465 8.555 2.71 ;
 RECT 6.705 0.705 6.805 1.17 ;
 RECT 6.705 0.47 6.99 0.705 ;
 RECT 6.12 1.17 6.805 1.27 ;
 RECT 6.12 1.27 6.365 1.46 ;
 RECT 13.85 0.19 13.95 1.795 ;
 RECT 13.85 0.09 15.565 0.19 ;
 RECT 8.945 0.47 9.13 0.5 ;
 RECT 13.155 1.71 13.255 1.795 ;
 RECT 15.465 0.19 15.565 1.18 ;
 RECT 13.155 1.795 13.95 1.895 ;
 RECT 12.135 0.47 12.235 1.61 ;
 RECT 12.685 1.71 12.785 2.445 ;
 RECT 8.9 0.5 9.13 0.71 ;
 RECT 8.945 0.37 12.235 0.47 ;
 RECT 12.135 1.61 13.255 1.71 ;
 RECT 15.46 1.635 15.56 1.66 ;
 RECT 15.46 1.87 15.56 2.565 ;
 RECT 15.46 1.66 15.715 1.87 ;
 RECT 14.615 0.64 14.715 1.26 ;
 RECT 14.41 1.26 14.715 1.47 ;
 RECT 14.615 1.47 14.715 2.21 ;
 RECT 10.325 1.45 10.425 1.655 ;
 RECT 10.325 1.755 10.425 2.57 ;
 RECT 10.325 1.655 11.285 1.755 ;
 RECT 11.185 1.755 11.285 2.355 ;
 RECT 10.325 0.655 10.425 1.13 ;
 RECT 10.325 1.23 10.425 1.24 ;
 RECT 9.41 0.66 9.51 1.13 ;
 RECT 10.325 1.24 10.58 1.45 ;
 RECT 9.41 1.13 10.425 1.23 ;
 RECT 24.955 0.37 25.055 1.01 ;
 RECT 24.955 1.01 25.205 1.22 ;
 RECT 24.955 1.22 25.055 2.245 ;
 RECT 24.955 2.245 25.24 2.455 ;
 RECT 9.4 1.575 9.5 2.485 ;
 RECT 9.91 1.41 10.14 1.475 ;
 RECT 9.4 1.475 10.14 1.575 ;
 RECT 9.91 1.575 10.14 1.62 ;
 RECT 22.56 0.19 22.66 0.97 ;
 RECT 22.56 0.97 22.8 1.18 ;
 RECT 22.56 1.18 22.66 1.975 ;
 RECT 21.78 0.87 21.88 2.175 ;
 RECT 20.815 0.77 22.35 0.78 ;
 RECT 21.78 0.73 22.35 0.77 ;
 RECT 21.78 2.175 24.58 2.275 ;
 RECT 24.48 1.125 24.58 2.175 ;
 RECT 20.82 0.78 22.35 0.83 ;
 RECT 20.82 0.83 21.88 0.87 ;
 RECT 22.25 0.19 22.35 0.73 ;
 RECT 21.78 0.185 21.88 0.73 ;
 RECT 20.815 0.57 21.045 0.77 ;
 RECT 15.735 1.25 15.995 1.3 ;
 RECT 15.895 0.61 15.995 1.25 ;
 LAYER CO ;
 RECT 24.025 0.295 24.155 0.425 ;
 RECT 22.62 1.01 22.75 1.14 ;
 RECT 16.46 0.67 16.59 0.8 ;
 RECT 22.17 1.05 22.3 1.18 ;
 RECT 11.875 0.875 12.005 1.005 ;
 RECT 7.325 1.525 7.455 1.655 ;
 RECT 4.345 0.325 4.475 0.455 ;
 RECT 24.395 0.115 24.525 0.245 ;
 RECT 23.215 0.11 23.345 0.24 ;
 RECT 21.53 1.4 21.66 1.53 ;
 RECT 23.695 0.59 23.825 0.72 ;
 RECT 3.745 2.05 3.875 2.18 ;
 RECT 1.37 1.55 1.5 1.68 ;
 RECT 3.275 2.09 3.405 2.22 ;
 RECT 2.49 1.23 2.62 1.36 ;
 RECT 1.365 2.315 1.495 2.445 ;
 RECT 2.67 1.64 2.8 1.77 ;
 RECT 24.23 1.465 24.36 1.595 ;
 RECT 23.385 1.42 23.515 1.55 ;
 RECT 25.175 1.44 25.305 1.57 ;
 RECT 22 1.45 22.13 1.58 ;
 RECT 12.905 1.87 13.035 2 ;
 RECT 4.865 1.55 4.995 1.68 ;
 RECT 6.925 0.88 7.055 1.01 ;
 RECT 12.4 0.595 12.53 0.725 ;
 RECT 10.075 1.885 10.205 2.015 ;
 RECT 5.995 1.825 6.125 1.955 ;
 RECT 12.4 1.9 12.53 2.03 ;
 RECT 8.205 2.125 8.335 2.255 ;
 RECT 4.275 2.115 4.405 2.245 ;
 RECT 25.175 0.59 25.305 0.72 ;
 RECT 22.78 1.46 22.91 1.59 ;
 RECT 22.78 0.41 22.91 0.54 ;
 RECT 23.86 1.38 23.99 1.51 ;
 RECT 21.28 0.505 21.41 0.635 ;
 RECT 25.955 1.45 26.085 1.58 ;
 RECT 22 0.11 22.13 0.24 ;
 RECT 6.905 2.07 7.035 2.2 ;
 RECT 15.21 2.64 15.34 2.77 ;
 RECT 0.39 2.085 0.52 2.215 ;
 RECT 10.775 2.445 10.905 2.575 ;
 RECT 4.275 0.79 4.405 0.92 ;
 RECT 14.365 2.64 14.495 2.77 ;
 RECT 17.79 0.975 17.92 1.105 ;
 RECT 0.39 1.825 0.52 1.955 ;
 RECT 14.835 1.705 14.965 1.835 ;
 RECT 6.81 0.525 6.94 0.655 ;
 RECT 6.455 0.88 6.585 1.01 ;
 RECT 18.31 0.77 18.44 0.9 ;
 RECT 8.28 2.515 8.41 2.645 ;
 RECT 8.135 0.455 8.265 0.585 ;
 RECT 6.06 0.905 6.19 1.035 ;
 RECT 16.115 0.83 16.245 0.96 ;
 RECT 19.37 0.78 19.5 0.91 ;
 RECT 14.14 0.955 14.27 1.085 ;
 RECT 4.745 2.05 4.875 2.18 ;
 RECT 10.965 0.62 11.095 0.75 ;
 RECT 6.41 2.105 6.54 2.235 ;
 RECT 9.63 2.07 9.76 2.2 ;
 RECT 8.675 2.135 8.805 2.265 ;
 RECT 8.815 1.63 8.945 1.76 ;
 RECT 18.31 1.725 18.44 1.855 ;
 RECT 5.35 0.88 5.48 1.01 ;
 RECT 9.63 0.88 9.76 1.01 ;
 RECT 14.835 0.96 14.965 1.09 ;
 RECT 0.39 2.345 0.52 2.475 ;
 RECT 4.745 0.79 4.875 0.92 ;
 RECT 9.145 0.93 9.275 1.06 ;
 RECT 1.365 0.775 1.495 0.905 ;
 RECT 3.275 2.35 3.405 2.48 ;
 RECT 2.505 2.115 2.635 2.245 ;
 RECT 1.365 2.055 1.495 2.185 ;
 RECT 0.895 2.055 1.025 2.185 ;
 RECT 3.745 1.79 3.875 1.92 ;
 RECT 1.97 1.195 2.1 1.325 ;
 RECT 3.385 1.195 3.515 1.325 ;
 RECT 2.9 0.225 3.03 0.355 ;
 RECT 0.895 0.775 1.025 0.905 ;
 RECT 3.745 0.775 3.875 0.905 ;
 RECT 3.275 0.585 3.405 0.715 ;
 RECT 2.31 0.775 2.44 0.905 ;
 RECT 16.785 0.975 16.915 1.105 ;
 RECT 5.49 0.21 5.62 0.34 ;
 RECT 17.27 2.64 17.4 2.77 ;
 RECT 9.145 2.015 9.275 2.145 ;
 RECT 7.415 2.125 7.545 2.255 ;
 RECT 5.485 2.345 5.615 2.475 ;
 RECT 18.59 1.25 18.72 1.38 ;
 RECT 0.355 0.33 0.485 0.46 ;
 RECT 15.535 1.7 15.665 1.83 ;
 RECT 23.13 1.025 23.26 1.155 ;
 RECT 6.175 1.265 6.305 1.395 ;
 RECT 25.025 1.05 25.155 1.18 ;
 RECT 14.46 1.3 14.59 1.43 ;
 RECT 21.125 1.135 21.255 1.265 ;
 RECT 13.49 1.445 13.62 1.575 ;
 RECT 13.14 2.37 13.27 2.5 ;
 RECT 20.865 0.61 20.995 0.74 ;
 RECT 8.95 0.54 9.08 0.67 ;
 RECT 9.96 1.45 10.09 1.58 ;
 RECT 0.355 0.59 0.485 0.72 ;
 RECT 11.875 1.945 12.005 2.075 ;
 RECT 10.075 0.88 10.205 1.01 ;
 RECT 5.4 1.495 5.53 1.625 ;
 RECT 18.785 2.64 18.915 2.77 ;
 RECT 11.14 1.28 11.27 1.41 ;
 RECT 16.785 1.72 16.915 1.85 ;
 RECT 5.22 1.995 5.35 2.125 ;
 RECT 19.37 1.71 19.5 1.84 ;
 RECT 15.215 0.33 15.345 0.46 ;
 RECT 17.79 1.72 17.92 1.85 ;
 RECT 12.905 0.595 13.035 0.725 ;
 RECT 16.115 1.78 16.245 1.91 ;
 RECT 17.275 0.305 17.405 0.435 ;
 RECT 18.87 0.77 19 0.9 ;
 RECT 15.785 1.29 15.915 1.42 ;
 RECT 10.4 1.28 10.53 1.41 ;
 RECT 25.06 2.285 25.19 2.415 ;
 RECT 19.865 0.265 19.995 0.395 ;
 RECT 16.09 0.265 16.22 0.395 ;
 LAYER M1 ;
 RECT 23.08 0.985 23.31 1.195 ;
 RECT 22.775 0.565 23.235 0.705 ;
 RECT 6.74 0.52 7.34 0.66 ;
 RECT 7.2 0.66 7.34 1.015 ;
 RECT 8.745 0.505 9.13 0.71 ;
 RECT 8.9 0.5 9.13 0.505 ;
 RECT 7.2 1.015 8.885 1.155 ;
 RECT 8.745 0.71 8.885 1.015 ;
 RECT 6.055 1.435 6.195 1.82 ;
 RECT 6.055 1.96 6.195 2.51 ;
 RECT 6.055 0.5 6.195 1.225 ;
 RECT 6.055 1.225 6.355 1.435 ;
 RECT 5.925 1.82 6.195 1.96 ;
 RECT 6.055 2.51 8.53 2.65 ;
 RECT 13.09 2.42 13.32 2.54 ;
 RECT 13.09 2.28 20.695 2.42 ;
 RECT 20.555 2.42 20.695 2.505 ;
 RECT 25.01 2.455 25.15 2.505 ;
 RECT 20.555 2.505 25.15 2.645 ;
 RECT 25.01 2.245 25.24 2.455 ;
 RECT 3.74 0.57 3.88 2.25 ;
 RECT 4.235 0.22 4.6 0.43 ;
 RECT 3.74 0.43 4.6 0.57 ;
 RECT 4.235 0.57 4.6 0.615 ;
 RECT 14.415 0.805 14.555 1.26 ;
 RECT 14.41 1.26 14.64 1.295 ;
 RECT 14.41 1.435 14.64 1.47 ;
 RECT 13.82 1.295 14.64 1.435 ;
 RECT 13.82 1.105 13.96 1.295 ;
 RECT 12.9 0.525 13.04 0.965 ;
 RECT 12.9 1.105 13.04 2.065 ;
 RECT 12.9 0.965 13.96 1.105 ;
 RECT 16.11 0.435 16.25 0.665 ;
 RECT 16.11 0.805 16.25 1.98 ;
 RECT 14.415 0.665 16.25 0.805 ;
 RECT 16.11 0.22 16.25 0.225 ;
 RECT 16.04 0.225 16.27 0.435 ;
 RECT 24.065 0.465 24.205 0.685 ;
 RECT 23.975 0.255 24.205 0.465 ;
 RECT 24.065 0.685 25.625 0.825 ;
 RECT 25.485 0.825 25.625 1.36 ;
 RECT 25.17 1.5 25.31 1.705 ;
 RECT 25.17 0.485 25.31 0.685 ;
 RECT 25.17 1.36 25.625 1.5 ;
 RECT 19.815 0.36 20.045 0.435 ;
 RECT 21.63 0.36 21.77 0.54 ;
 RECT 19.815 0.225 21.77 0.36 ;
 RECT 19.85 0.22 21.77 0.225 ;
 RECT 22.495 0.535 22.635 0.54 ;
 RECT 22.495 0.68 22.635 0.97 ;
 RECT 21.63 0.54 22.635 0.68 ;
 RECT 22.495 0.97 22.8 1.18 ;
 RECT 14.83 1.37 15.965 1.46 ;
 RECT 14.83 1.095 14.97 1.37 ;
 RECT 14.83 1.46 15.96 1.51 ;
 RECT 14.83 1.51 14.97 1.7 ;
 RECT 15.735 1.25 15.965 1.37 ;
 RECT 14.765 1.7 15.04 1.84 ;
 RECT 14.76 0.955 15.03 1.095 ;
 RECT 16.41 0.72 16.64 0.84 ;
 RECT 17.68 0.37 17.82 0.58 ;
 RECT 16.41 0.63 17.82 0.72 ;
 RECT 16.42 0.58 17.82 0.63 ;
 RECT 18.585 0.37 18.725 1.46 ;
 RECT 17.68 0.23 18.725 0.37 ;
 RECT 21.525 1.2 21.665 1.725 ;
 RECT 21.075 1.17 21.665 1.2 ;
 RECT 21.35 0.64 21.49 0.99 ;
 RECT 21.075 1.2 21.305 1.305 ;
 RECT 21.215 0.99 21.525 1.03 ;
 RECT 21.23 0.5 21.49 0.64 ;
 RECT 22.12 1.01 22.35 1.03 ;
 RECT 21.07 1.03 22.35 1.17 ;
 RECT 22.12 1.17 22.35 1.22 ;
 RECT 9.625 0.82 9.765 2.225 ;
 RECT 10.475 2.165 10.615 2.225 ;
 RECT 9.625 2.225 10.615 2.365 ;
 RECT 12.395 0.525 12.535 2.025 ;
 RECT 11.87 0.765 12.01 2.025 ;
 RECT 10.475 2.025 12.535 2.165 ;
 RECT 23.69 0.48 23.83 1.08 ;
 RECT 23.855 1.22 23.995 1.58 ;
 RECT 24.975 1.01 25.205 1.08 ;
 RECT 23.69 1.08 25.205 1.22 ;
 RECT 5.26 1.63 5.4 1.99 ;
 RECT 5.26 1.475 5.605 1.63 ;
 RECT 5.345 0.81 5.485 1.475 ;
 RECT 5.15 1.99 5.4 2.13 ;
 RECT 4.05 0.925 4.19 1.195 ;
 RECT 4.05 1.335 4.19 2.11 ;
 RECT 4.05 0.785 4.475 0.925 ;
 RECT 4.05 2.11 4.475 2.25 ;
 RECT 4.05 1.195 5.16 1.335 ;
 RECT 5.02 0.67 5.16 1.195 ;
 RECT 5.765 0.22 6.59 0.36 ;
 RECT 6.45 0.36 6.59 0.9 ;
 RECT 6.525 1.08 6.665 1.945 ;
 RECT 5.02 0.53 5.905 0.67 ;
 RECT 5.765 0.36 5.905 0.53 ;
 RECT 6.45 0.9 6.665 1.08 ;
 RECT 6.405 1.945 6.665 2.17 ;
 RECT 6.405 2.17 6.545 2.305 ;
 RECT 10.07 0.81 10.21 1.41 ;
 RECT 9.91 1.41 10.21 1.62 ;
 RECT 10.07 1.62 10.21 1.735 ;
 RECT 10.07 1.875 10.21 2.085 ;
 RECT 11.12 1.49 11.26 1.735 ;
 RECT 10.07 1.735 11.26 1.875 ;
 RECT 11.045 1.235 11.39 1.49 ;
 RECT 0.89 0.72 1.03 1.195 ;
 RECT 0.89 1.335 1.03 2.27 ;
 RECT 1.675 0.36 1.815 1.195 ;
 RECT 0.89 1.195 1.815 1.335 ;
 RECT 1.675 0.22 3.1 0.36 ;
 RECT 8.185 1.79 8.325 1.82 ;
 RECT 6.92 0.805 7.06 1.82 ;
 RECT 6.83 1.96 7.11 2.215 ;
 RECT 6.83 1.82 8.325 1.96 ;
 RECT 8.76 1.58 9 1.65 ;
 RECT 8.185 1.65 9 1.79 ;
 RECT 8.76 1.79 9 1.835 ;
 RECT 15.485 1.87 15.67 1.985 ;
 RECT 13.435 1.43 13.67 1.615 ;
 RECT 13.435 1.615 13.575 1.985 ;
 RECT 13.44 1.405 13.67 1.43 ;
 RECT 13.435 1.985 15.67 2.125 ;
 RECT 15.485 1.66 15.715 1.87 ;
 RECT 7.255 1.52 8.005 1.66 ;
 RECT 7.865 1.44 8.005 1.52 ;
 RECT 9.14 0.865 9.28 1.3 ;
 RECT 9.14 1.44 9.28 2.215 ;
 RECT 7.865 1.3 9.28 1.44 ;
 RECT 7.305 2.12 8.405 2.26 ;
 RECT 2.96 0.91 3.1 1.19 ;
 RECT 2.96 1.33 3.1 2.11 ;
 RECT 2.255 0.77 3.1 0.91 ;
 RECT 2.45 2.11 3.1 2.25 ;
 RECT 3.38 1.145 3.52 1.19 ;
 RECT 3.38 1.33 3.52 1.375 ;
 RECT 2.96 1.19 3.52 1.33 ;
 RECT 23.08 1.195 23.22 1.32 ;
 RECT 22.775 1.46 22.915 1.735 ;
 RECT 23.095 0.705 23.235 0.985 ;
 RECT 22.775 0.33 22.915 0.565 ;
 RECT 22.775 1.32 23.22 1.46 ;
 END
END RSDFFNSRX1

MACRO RSDFFNSRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.84 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.08 1.16 18.435 1.4 ;
 RECT 18.205 0.695 18.345 1.16 ;
 RECT 18.205 1.765 20.42 1.905 ;
 RECT 18.205 1.4 18.345 1.765 ;
 RECT 20.28 0.71 20.42 1.765 ;
 RECT 19.335 0.71 19.475 1.765 ;
 END
 ANTENNADIFFAREA 1.112 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 27.84 2.96 ;
 RECT 1.36 2.005 1.5 2.8 ;
 RECT 5.415 2.34 5.665 2.8 ;
 RECT 14.645 2.57 14.785 2.8 ;
 RECT 10.77 2.375 10.91 2.8 ;
 RECT 4.74 1.98 4.88 2.8 ;
 RECT 18.68 2.57 18.82 2.8 ;
 RECT 3.27 2.03 3.41 2.8 ;
 RECT 0.385 1.74 0.525 2.8 ;
 RECT 16.38 2.57 16.52 2.8 ;
 RECT 19.665 2.57 19.805 2.8 ;
 RECT 13.8 2.57 13.94 2.8 ;
 RECT 8.67 2.07 8.81 2.8 ;
 RECT 17.33 2.57 17.47 2.8 ;
 END
 END VDD

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.18 1.475 1.705 1.75 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.79 1.475 5.12 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.82 0.57 21.3 0.78 ;
 RECT 20.82 0.565 21.19 0.57 ;
 RECT 20.82 0.78 21.19 0.865 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 27.84 0.08 ;
 RECT 16.88 0.28 17.145 0.44 ;
 RECT 3.27 0.08 3.41 0.78 ;
 RECT 8.085 0.08 8.32 0.595 ;
 RECT 4.74 0.08 4.88 1.055 ;
 RECT 24.6 0.08 24.84 0.31 ;
 RECT 22.25 0.08 22.39 0.31 ;
 RECT 13.575 0.08 13.715 1.155 ;
 RECT 5.485 0.08 5.625 0.39 ;
 RECT 0.35 0.08 0.49 0.775 ;
 RECT 18.865 0.08 19.005 0.965 ;
 RECT 10.96 0.08 11.1 0.815 ;
 RECT 23.465 0.08 23.605 0.325 ;
 RECT 19.81 0.08 19.95 0.965 ;
 RECT 14.65 0.08 14.79 0.525 ;
 RECT 1.36 0.08 1.5 0.97 ;
 RECT 16.935 0.08 17.075 0.28 ;
 END
 END VSS

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.965 1.13 2.105 1.48 ;
 RECT 1.87 1.63 2.815 1.79 ;
 RECT 1.87 1.48 2.115 1.63 ;
 RECT 2.665 1.79 2.805 1.845 ;
 RECT 2.665 1.57 2.805 1.63 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.16 1.41 26.5 1.775 ;
 RECT 24.48 1.965 26.345 2.105 ;
 RECT 22.25 2.195 24.62 2.335 ;
 RECT 26.205 1.775 26.345 1.965 ;
 RECT 24.48 1.41 24.62 1.965 ;
 RECT 22.25 1.365 22.39 2.195 ;
 RECT 23.635 1.345 23.775 2.195 ;
 RECT 24.48 2.105 24.62 2.195 ;
 END
 END VDDG

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.35 1.16 10.68 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.33 1.155 2.75 1.415 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 16.245 1.205 16.6 1.445 ;
 RECT 15.85 1.705 18.005 1.845 ;
 RECT 16.455 0.88 16.595 1.205 ;
 RECT 17.465 0.89 17.605 1.705 ;
 RECT 16.455 1.445 16.595 1.705 ;
 END
 ANTENNADIFFAREA 0.794 ;
 END QN

 OBS
 LAYER PO ;
 RECT 4.525 0.52 4.625 2.465 ;
 RECT 4.285 0.27 4.625 0.52 ;
 RECT 11.22 0.655 11.32 1.24 ;
 RECT 11.09 1.24 11.32 1.475 ;
 RECT 16.71 0.39 16.81 1.4 ;
 RECT 17.19 0.37 17.29 1.4 ;
 RECT 17.585 1.5 17.685 2.275 ;
 RECT 16.17 1.4 17.685 1.5 ;
 RECT 16.17 1.5 16.27 2.275 ;
 RECT 17.12 1.5 17.22 2.275 ;
 RECT 16.645 1.5 16.745 2.275 ;
 RECT 15.84 0.29 16.81 0.39 ;
 RECT 15.84 0.22 16.07 0.29 ;
 RECT 15.84 0.39 16.07 0.43 ;
 RECT 8.76 1.61 9.025 1.82 ;
 RECT 8.925 1.82 9.025 2.49 ;
 RECT 8.555 0.66 8.655 1.51 ;
 RECT 8.555 1.51 9.025 1.61 ;
 RECT 3.055 0.405 3.155 2.735 ;
 RECT 2.85 0.175 3.155 0.405 ;
 RECT 11.615 2.69 13.265 2.695 ;
 RECT 13.09 2.54 13.265 2.69 ;
 RECT 12.405 2.695 13.265 2.79 ;
 RECT 11.615 0.655 11.715 2.595 ;
 RECT 11.615 2.595 12.505 2.69 ;
 RECT 13.09 2.33 13.32 2.54 ;
 RECT 21.275 1.175 21.56 1.305 ;
 RECT 21.275 1.305 21.375 2.64 ;
 RECT 24.9 0.19 25 0.94 ;
 RECT 24.9 0.09 26.01 0.19 ;
 RECT 25.91 0.19 26.01 2.64 ;
 RECT 21.275 1.075 21.605 1.175 ;
 RECT 21.275 2.64 26.01 2.74 ;
 RECT 1.95 0.555 2.05 1.145 ;
 RECT 1.91 1.145 2.155 1.385 ;
 RECT 22.035 0.87 22.135 2.175 ;
 RECT 21.07 0.77 22.605 0.78 ;
 RECT 22.035 0.73 22.605 0.77 ;
 RECT 24.735 1.125 24.835 2.175 ;
 RECT 21.075 0.78 22.605 0.83 ;
 RECT 21.075 0.83 22.135 0.87 ;
 RECT 22.505 0.19 22.605 0.73 ;
 RECT 22.035 0.185 22.135 0.73 ;
 RECT 21.07 0.57 21.3 0.77 ;
 RECT 22.035 2.175 24.835 2.275 ;
 RECT 14.055 0.64 14.155 1.26 ;
 RECT 13.85 1.26 14.155 1.47 ;
 RECT 14.055 1.47 14.155 2.21 ;
 RECT 18.46 1.2 18.76 1.285 ;
 RECT 18.46 0.525 18.56 1.2 ;
 RECT 18.46 1.285 20.17 1.385 ;
 RECT 20.065 0.36 20.165 1.285 ;
 RECT 18.46 1.435 18.56 2.645 ;
 RECT 18.46 1.385 18.76 1.435 ;
 RECT 18.95 1.385 19.05 2.645 ;
 RECT 19.59 0.525 19.69 1.285 ;
 RECT 19.92 1.385 20.02 2.645 ;
 RECT 19.445 1.385 19.545 2.645 ;
 RECT 19.12 0.52 19.22 1.285 ;
 RECT 20.36 0.19 20.59 0.26 ;
 RECT 20.36 0.36 20.59 0.435 ;
 RECT 20.065 0.26 20.59 0.36 ;
 RECT 23.725 0.355 23.825 0.985 ;
 RECT 23.895 1.215 23.995 1.815 ;
 RECT 23.335 1.115 23.995 1.215 ;
 RECT 23.335 0.985 23.825 1.115 ;
 RECT 24.23 0.355 24.46 0.465 ;
 RECT 23.725 0.255 24.46 0.355 ;
 RECT 3.525 0.335 3.625 1.155 ;
 RECT 3.525 1.365 3.625 2.745 ;
 RECT 3.335 1.155 3.625 1.365 ;
 RECT 2.755 1.82 2.855 2.735 ;
 RECT 2.615 1.59 2.855 1.82 ;
 RECT 8.455 1.79 8.555 2.465 ;
 RECT 8.24 2.465 8.555 2.71 ;
 RECT 7.195 1.475 7.505 1.71 ;
 RECT 7.195 0.65 7.295 1.475 ;
 RECT 7.195 1.71 7.295 2.475 ;
 RECT 12.65 0.19 12.75 1.29 ;
 RECT 12.65 1.29 13.555 1.39 ;
 RECT 5.84 0.285 5.94 1.52 ;
 RECT 5.34 1.52 5.94 1.62 ;
 RECT 6.66 1.565 6.76 2.375 ;
 RECT 13.325 1.39 13.555 1.82 ;
 RECT 5.775 1.62 5.875 2.375 ;
 RECT 5.34 1.44 5.585 1.52 ;
 RECT 5.34 1.62 5.585 1.69 ;
 RECT 5.84 0.185 12.75 0.19 ;
 RECT 7.895 0.09 12.75 0.185 ;
 RECT 5.84 0.19 7.995 0.285 ;
 RECT 7.895 0.285 7.995 1.24 ;
 RECT 5.775 2.375 6.76 2.475 ;
 RECT 1.145 1.475 1.715 1.75 ;
 RECT 1.145 0.555 1.245 1.475 ;
 RECT 1.145 1.75 1.245 2.685 ;
 RECT 1.615 0.555 1.715 1.475 ;
 RECT 1.615 1.75 1.715 2.735 ;
 RECT 2.565 0.555 2.665 1.18 ;
 RECT 2.335 1.41 2.435 1.645 ;
 RECT 2.335 1.18 2.665 1.41 ;
 RECT 2.285 1.645 2.435 1.745 ;
 RECT 2.285 1.745 2.385 2.735 ;
 RECT 13.19 0.09 15.005 0.19 ;
 RECT 14.905 0.19 15.005 1.18 ;
 RECT 13.19 0.19 13.42 0.45 ;
 RECT 8.945 0.47 9.13 0.5 ;
 RECT 12.685 1.71 12.785 2.445 ;
 RECT 12 0.47 12.235 0.59 ;
 RECT 12.135 0.59 12.235 1.61 ;
 RECT 8.9 0.5 9.13 0.71 ;
 RECT 12.135 1.61 12.785 1.71 ;
 RECT 8.945 0.37 12.235 0.47 ;
 RECT 14.9 1.635 15 1.66 ;
 RECT 14.9 1.66 15.155 1.87 ;
 RECT 14.9 1.87 15 2.565 ;
 RECT 25.21 2.245 25.495 2.455 ;
 RECT 25.21 1.22 25.31 2.245 ;
 RECT 25.21 0.37 25.31 1.01 ;
 RECT 25.21 1.01 25.46 1.22 ;
 RECT 22.375 1.01 22.61 1.22 ;
 RECT 22.51 1.22 22.61 1.995 ;
 RECT 9.4 1.575 9.5 2.485 ;
 RECT 9.91 1.41 10.14 1.475 ;
 RECT 9.91 1.575 10.14 1.62 ;
 RECT 9.4 1.475 10.14 1.575 ;
 RECT 10.325 1.45 10.425 1.655 ;
 RECT 10.325 1.755 10.425 2.57 ;
 RECT 10.325 1.655 11.285 1.755 ;
 RECT 11.185 1.755 11.285 2.355 ;
 RECT 10.325 0.655 10.425 1.13 ;
 RECT 10.325 1.23 10.425 1.24 ;
 RECT 9.41 0.66 9.51 1.13 ;
 RECT 10.325 1.24 10.58 1.45 ;
 RECT 9.41 1.13 10.425 1.23 ;
 RECT 15.335 1.195 15.435 1.25 ;
 RECT 15.18 1.25 15.435 1.46 ;
 RECT 15.335 1.46 15.435 2.56 ;
 RECT 15.865 0.84 15.965 1.095 ;
 RECT 15.335 0.61 15.435 1.095 ;
 RECT 15.335 1.095 15.965 1.195 ;
 RECT 15.85 0.63 16.08 0.84 ;
 RECT 22.815 0.19 22.915 0.97 ;
 RECT 22.815 0.97 23.055 1.18 ;
 RECT 22.815 1.18 22.915 1.975 ;
 RECT 5 0.57 5.1 1.495 ;
 RECT 4.805 1.495 5.1 1.745 ;
 RECT 5 1.745 5.1 2.37 ;
 RECT 6.705 0.705 6.805 1.17 ;
 RECT 6.12 1.17 6.805 1.27 ;
 RECT 6.12 1.27 6.365 1.46 ;
 RECT 6.705 0.47 6.99 0.705 ;
 LAYER CO ;
 RECT 11.875 0.875 12.005 1.005 ;
 RECT 25.43 1.44 25.56 1.57 ;
 RECT 17.805 1.71 17.935 1.84 ;
 RECT 5.22 1.995 5.35 2.125 ;
 RECT 12.4 0.595 12.53 0.725 ;
 RECT 6.06 0.905 6.19 1.035 ;
 RECT 19.185 1.77 19.315 1.9 ;
 RECT 12.4 1.9 12.53 2.03 ;
 RECT 7.325 1.525 7.455 1.655 ;
 RECT 6.81 0.525 6.94 0.655 ;
 RECT 4.865 1.55 4.995 1.68 ;
 RECT 23.64 1.42 23.77 1.55 ;
 RECT 10.075 1.885 10.205 2.015 ;
 RECT 18.87 0.77 19 0.9 ;
 RECT 18.685 2.64 18.815 2.77 ;
 RECT 6.925 0.88 7.055 1.01 ;
 RECT 3.745 0.775 3.875 0.905 ;
 RECT 14.275 0.96 14.405 1.09 ;
 RECT 7.415 2.125 7.545 2.255 ;
 RECT 21.535 0.505 21.665 0.635 ;
 RECT 8.205 2.125 8.335 2.255 ;
 RECT 3.275 2.35 3.405 2.48 ;
 RECT 0.355 0.59 0.485 0.72 ;
 RECT 4.275 2.115 4.405 2.245 ;
 RECT 14.655 0.33 14.785 0.46 ;
 RECT 0.895 2.055 1.025 2.185 ;
 RECT 10.075 0.88 10.205 1.01 ;
 RECT 1.365 2.055 1.495 2.185 ;
 RECT 11.875 1.945 12.005 2.075 ;
 RECT 15.555 1.78 15.685 1.91 ;
 RECT 1.365 0.775 1.495 0.905 ;
 RECT 11.14 1.28 11.27 1.41 ;
 RECT 16.46 0.95 16.59 1.08 ;
 RECT 12.905 0.595 13.035 0.725 ;
 RECT 1.97 1.195 2.1 1.325 ;
 RECT 22.255 1.45 22.385 1.58 ;
 RECT 3.275 0.585 3.405 0.715 ;
 RECT 6.905 2.07 7.035 2.2 ;
 RECT 15.555 0.83 15.685 0.96 ;
 RECT 2.505 2.115 2.635 2.245 ;
 RECT 19.34 0.79 19.47 0.92 ;
 RECT 9.145 2.015 9.275 2.145 ;
 RECT 26.21 1.45 26.34 1.58 ;
 RECT 3.385 1.195 3.515 1.325 ;
 RECT 5.485 2.345 5.615 2.475 ;
 RECT 13.805 2.64 13.935 2.77 ;
 RECT 10.775 2.445 10.905 2.575 ;
 RECT 3.745 2.05 3.875 2.18 ;
 RECT 21.12 0.61 21.25 0.74 ;
 RECT 8.95 0.54 9.08 0.67 ;
 RECT 13.9 1.3 14.03 1.43 ;
 RECT 20.41 0.265 20.54 0.395 ;
 RECT 24.28 0.295 24.41 0.425 ;
 RECT 22.255 0.11 22.385 0.24 ;
 RECT 23.035 0.41 23.165 0.54 ;
 RECT 18.59 1.25 18.72 1.38 ;
 RECT 25.43 0.59 25.56 0.72 ;
 RECT 9.63 2.07 9.76 2.2 ;
 RECT 0.895 0.775 1.025 0.905 ;
 RECT 1.365 2.315 1.495 2.445 ;
 RECT 8.675 2.135 8.805 2.265 ;
 RECT 17.335 2.64 17.465 2.77 ;
 RECT 4.345 0.325 4.475 0.455 ;
 RECT 23.035 1.46 23.165 1.59 ;
 RECT 24.115 1.38 24.245 1.51 ;
 RECT 24.485 1.465 24.615 1.595 ;
 RECT 2.31 0.775 2.44 0.905 ;
 RECT 4.745 0.79 4.875 0.92 ;
 RECT 14.275 1.705 14.405 1.835 ;
 RECT 8.135 0.455 8.265 0.585 ;
 RECT 17.47 0.96 17.6 1.09 ;
 RECT 8.28 2.515 8.41 2.645 ;
 RECT 6.455 0.88 6.585 1.01 ;
 RECT 5.4 1.495 5.53 1.625 ;
 RECT 5.995 1.825 6.125 1.955 ;
 RECT 4.275 0.79 4.405 0.92 ;
 RECT 13.58 0.955 13.71 1.085 ;
 RECT 16.87 1.71 17 1.84 ;
 RECT 2.9 0.225 3.03 0.355 ;
 RECT 5.35 0.88 5.48 1.01 ;
 RECT 0.355 0.33 0.485 0.46 ;
 RECT 18.21 0.77 18.34 0.9 ;
 RECT 5.49 0.21 5.62 0.34 ;
 RECT 3.745 1.79 3.875 1.92 ;
 RECT 9.145 0.93 9.275 1.06 ;
 RECT 6.41 2.105 6.54 2.235 ;
 RECT 13.24 0.28 13.37 0.41 ;
 RECT 12.05 0.42 12.18 0.55 ;
 RECT 15.89 0.26 16.02 0.39 ;
 RECT 25.315 2.285 25.445 2.415 ;
 RECT 15.23 1.29 15.36 1.42 ;
 RECT 23.385 1.025 23.515 1.155 ;
 RECT 14.975 1.7 15.105 1.83 ;
 RECT 25.28 1.05 25.41 1.18 ;
 RECT 22.425 1.05 22.555 1.18 ;
 RECT 13.375 1.65 13.505 1.78 ;
 RECT 21.38 1.135 21.51 1.265 ;
 RECT 9.96 1.45 10.09 1.58 ;
 RECT 6.175 1.265 6.305 1.395 ;
 RECT 10.4 1.28 10.53 1.41 ;
 RECT 15.9 0.67 16.03 0.8 ;
 RECT 22.875 1.01 23.005 1.14 ;
 RECT 13.14 2.37 13.27 2.5 ;
 RECT 20.285 0.78 20.415 0.91 ;
 RECT 19.815 0.78 19.945 0.91 ;
 RECT 20.145 1.77 20.275 1.9 ;
 RECT 19.67 2.64 19.8 2.77 ;
 RECT 15.92 1.71 16.05 1.84 ;
 RECT 16.385 2.64 16.515 2.77 ;
 RECT 1.37 1.55 1.5 1.68 ;
 RECT 23.47 0.11 23.6 0.24 ;
 RECT 2.67 1.64 2.8 1.77 ;
 RECT 0.39 1.825 0.52 1.955 ;
 RECT 14.65 2.64 14.78 2.77 ;
 RECT 8.815 1.63 8.945 1.76 ;
 RECT 0.39 2.345 0.52 2.475 ;
 RECT 0.39 2.085 0.52 2.215 ;
 RECT 4.745 2.05 4.875 2.18 ;
 RECT 24.65 0.115 24.78 0.245 ;
 RECT 12.905 1.87 13.035 2 ;
 RECT 18.21 1.725 18.34 1.855 ;
 RECT 16.94 0.305 17.07 0.435 ;
 RECT 9.63 0.88 9.76 1.01 ;
 RECT 10.965 0.62 11.095 0.75 ;
 RECT 21.785 1.4 21.915 1.53 ;
 RECT 2.49 1.23 2.62 1.36 ;
 RECT 23.95 0.59 24.08 0.72 ;
 RECT 3.275 2.09 3.405 2.22 ;
 LAYER M1 ;
 RECT 14.27 1.395 14.41 1.7 ;
 RECT 15.18 1.25 15.41 1.255 ;
 RECT 15.18 1.395 15.41 1.46 ;
 RECT 14.205 1.7 14.48 1.84 ;
 RECT 14.2 0.955 14.47 1.095 ;
 RECT 23.335 1.195 23.475 1.32 ;
 RECT 23.03 1.46 23.17 1.735 ;
 RECT 23.35 0.705 23.49 0.985 ;
 RECT 23.03 0.33 23.17 0.565 ;
 RECT 23.03 1.32 23.475 1.46 ;
 RECT 23.03 0.565 23.49 0.705 ;
 RECT 23.335 0.985 23.565 1.195 ;
 RECT 10.07 1.62 10.21 1.735 ;
 RECT 10.07 1.875 10.21 2.085 ;
 RECT 10.07 0.81 10.21 1.41 ;
 RECT 9.91 1.41 10.21 1.62 ;
 RECT 10.07 1.735 11.27 1.875 ;
 RECT 11.13 1.415 11.27 1.735 ;
 RECT 11.09 1.275 11.34 1.415 ;
 RECT 6.055 1.435 6.195 1.82 ;
 RECT 6.055 1.96 6.195 2.51 ;
 RECT 6.055 0.5 6.195 1.225 ;
 RECT 6.055 1.225 6.355 1.435 ;
 RECT 5.925 1.82 6.195 1.96 ;
 RECT 6.055 2.51 8.53 2.65 ;
 RECT 15.85 0.72 16.08 0.84 ;
 RECT 17.345 0.37 17.485 0.58 ;
 RECT 15.85 0.58 17.485 0.72 ;
 RECT 18.585 0.37 18.725 1.46 ;
 RECT 17.345 0.23 18.725 0.37 ;
 RECT 13.09 2.42 13.32 2.54 ;
 RECT 20.81 2.42 20.95 2.505 ;
 RECT 13.09 2.28 20.95 2.42 ;
 RECT 25.265 2.455 25.405 2.505 ;
 RECT 25.265 2.245 25.495 2.455 ;
 RECT 20.81 2.505 25.405 2.645 ;
 RECT 21.605 0.64 21.745 0.99 ;
 RECT 21.33 1.17 21.92 1.2 ;
 RECT 21.78 1.2 21.92 1.725 ;
 RECT 21.47 0.99 21.78 1.03 ;
 RECT 21.33 1.2 21.56 1.305 ;
 RECT 21.485 0.5 21.745 0.64 ;
 RECT 22.375 1.01 22.605 1.03 ;
 RECT 21.325 1.03 22.605 1.17 ;
 RECT 22.375 1.17 22.605 1.22 ;
 RECT 9.625 0.82 9.765 2.225 ;
 RECT 10.475 2.165 10.615 2.225 ;
 RECT 9.625 2.225 10.615 2.365 ;
 RECT 12.395 0.525 12.535 2.025 ;
 RECT 11.87 0.765 12.01 2.025 ;
 RECT 10.475 2.025 12.535 2.165 ;
 RECT 23.945 0.48 24.085 1.08 ;
 RECT 24.11 1.22 24.25 1.58 ;
 RECT 25.23 1.01 25.46 1.08 ;
 RECT 23.945 1.08 25.46 1.22 ;
 RECT 0.89 0.72 1.03 1.195 ;
 RECT 0.89 1.335 1.03 2.27 ;
 RECT 1.675 0.36 1.815 1.195 ;
 RECT 0.89 1.195 1.815 1.335 ;
 RECT 1.675 0.22 3.1 0.36 ;
 RECT 6.74 0.52 7.34 0.66 ;
 RECT 7.2 0.66 7.34 1.015 ;
 RECT 8.745 0.505 9.13 0.71 ;
 RECT 8.9 0.5 9.13 0.505 ;
 RECT 7.2 1.015 8.885 1.155 ;
 RECT 8.745 0.71 8.885 1.015 ;
 RECT 20.36 0.36 20.59 0.435 ;
 RECT 21.885 0.36 22.025 0.54 ;
 RECT 20.35 0.22 22.025 0.36 ;
 RECT 22.75 0.97 23.055 1.18 ;
 RECT 22.75 0.68 22.89 0.97 ;
 RECT 21.885 0.54 22.89 0.68 ;
 RECT 22.75 0.535 22.89 0.54 ;
 RECT 24.32 0.465 24.46 0.685 ;
 RECT 24.23 0.255 24.46 0.465 ;
 RECT 25.74 0.825 25.88 1.36 ;
 RECT 24.32 0.685 25.88 0.825 ;
 RECT 25.425 1.5 25.565 1.705 ;
 RECT 25.425 0.485 25.565 0.685 ;
 RECT 25.425 1.36 25.88 1.5 ;
 RECT 13.855 0.805 13.995 1.26 ;
 RECT 13.85 1.26 14.08 1.3 ;
 RECT 13.85 1.44 14.08 1.47 ;
 RECT 12.9 1.3 14.08 1.44 ;
 RECT 12.9 0.525 13.04 1.3 ;
 RECT 12.9 1.44 13.04 2.065 ;
 RECT 13.855 0.665 15.69 0.805 ;
 RECT 15.55 0.43 15.69 0.665 ;
 RECT 15.55 0.805 15.69 1.98 ;
 RECT 15.55 0.22 16.07 0.43 ;
 RECT 4.05 0.925 4.19 1.195 ;
 RECT 4.05 1.335 4.19 2.11 ;
 RECT 4.05 0.785 4.475 0.925 ;
 RECT 4.05 2.11 4.475 2.25 ;
 RECT 4.05 1.195 5.16 1.335 ;
 RECT 5.02 0.67 5.16 1.195 ;
 RECT 5.765 0.22 6.59 0.36 ;
 RECT 6.45 0.36 6.59 0.9 ;
 RECT 6.525 1.08 6.665 1.945 ;
 RECT 5.02 0.53 5.905 0.67 ;
 RECT 5.765 0.36 5.905 0.53 ;
 RECT 6.45 0.9 6.665 1.08 ;
 RECT 6.405 1.945 6.665 2.17 ;
 RECT 6.405 2.17 6.545 2.305 ;
 RECT 14.925 1.87 15.11 1.985 ;
 RECT 13.355 1.82 13.495 1.985 ;
 RECT 13.355 1.985 15.11 2.125 ;
 RECT 14.925 1.66 15.155 1.87 ;
 RECT 13.325 1.61 13.555 1.82 ;
 RECT 3.74 0.57 3.88 2.25 ;
 RECT 4.235 0.22 4.6 0.43 ;
 RECT 4.235 0.57 4.6 0.615 ;
 RECT 3.74 0.43 4.6 0.57 ;
 RECT 5.26 1.63 5.4 1.99 ;
 RECT 5.345 0.81 5.485 1.475 ;
 RECT 5.26 1.475 5.605 1.63 ;
 RECT 5.15 1.99 5.4 2.13 ;
 RECT 8.185 1.79 8.325 1.82 ;
 RECT 6.92 0.805 7.06 1.82 ;
 RECT 6.83 1.96 7.11 2.215 ;
 RECT 6.83 1.82 8.325 1.96 ;
 RECT 8.76 1.58 9 1.65 ;
 RECT 8.185 1.65 9 1.79 ;
 RECT 8.76 1.79 9 1.835 ;
 RECT 13.19 0.38 13.42 0.45 ;
 RECT 12 0.24 13.435 0.38 ;
 RECT 12 0.38 12.23 0.59 ;
 RECT 2.96 0.91 3.1 1.19 ;
 RECT 2.96 1.33 3.1 2.11 ;
 RECT 2.255 0.77 3.1 0.91 ;
 RECT 2.45 2.11 3.1 2.25 ;
 RECT 2.96 1.19 3.52 1.33 ;
 RECT 3.38 1.145 3.52 1.19 ;
 RECT 3.38 1.33 3.52 1.375 ;
 RECT 7.865 1.44 8.005 1.52 ;
 RECT 7.255 1.52 8.005 1.66 ;
 RECT 9.14 0.865 9.28 1.3 ;
 RECT 7.865 1.3 9.28 1.44 ;
 RECT 9.14 1.44 9.28 2.215 ;
 RECT 7.305 2.12 8.405 2.26 ;
 RECT 14.27 1.095 14.41 1.255 ;
 RECT 14.27 1.255 15.41 1.395 ;
 END
END RSDFFNSRX2

MACRO RSDFFSRARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 28.48 BY 2.88 ;
 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.78 0.735 8.855 0.875 ;
 RECT 11.59 0.245 13.96 0.385 ;
 RECT 7.78 0.445 8.11 0.735 ;
 RECT 8.715 0.36 8.855 0.735 ;
 RECT 10.615 0.99 11.73 1.13 ;
 RECT 13.82 1.05 15.57 1.19 ;
 RECT 15.43 0.74 15.57 1.05 ;
 RECT 15.465 0.53 15.695 0.555 ;
 RECT 15.43 0.555 15.695 0.74 ;
 RECT 10.615 0.36 10.755 0.99 ;
 RECT 8.715 0.22 10.755 0.36 ;
 RECT 11.59 0.385 11.73 0.99 ;
 RECT 13.82 0.385 13.96 1.05 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 28.48 0.08 ;
 RECT 25.28 0.08 25.52 0.26 ;
 RECT 18.565 0.335 18.87 0.475 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.995 0.08 5.135 1.055 ;
 RECT 3.32 0.08 3.46 0.85 ;
 RECT 5.74 0.08 5.88 0.39 ;
 RECT 8.34 0.08 8.575 0.595 ;
 RECT 11.215 0.08 11.355 0.815 ;
 RECT 14.775 0.08 14.915 0.5 ;
 RECT 16.58 0.08 16.72 0.525 ;
 RECT 22.93 0.08 23.07 0.36 ;
 RECT 20.345 0.08 20.485 0.82 ;
 RECT 24.145 0.08 24.285 0.35 ;
 RECT 1.345 0.08 1.595 0.255 ;
 RECT 18.65 0.08 18.79 0.335 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 28.48 2.96 ;
 RECT 1.41 2.005 1.55 2.8 ;
 RECT 0.295 1.74 0.435 2.8 ;
 RECT 5.67 2.34 5.92 2.8 ;
 RECT 3.32 2.03 3.46 2.8 ;
 RECT 4.995 1.98 5.135 2.8 ;
 RECT 8.925 2.07 9.065 2.8 ;
 RECT 11.025 2.375 11.165 2.8 ;
 RECT 15.25 2.57 15.39 2.8 ;
 RECT 16.575 2.57 16.715 2.8 ;
 RECT 18.67 2.57 18.81 2.8 ;
 RECT 20.26 2.57 20.4 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5 1.475 5.375 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.08 1.15 19.32 1.4 ;
 RECT 19.12 0.915 19.26 1.15 ;
 RECT 18.18 1.765 19.26 1.905 ;
 RECT 19.12 1.4 19.26 1.765 ;
 RECT 18.18 0.905 18.32 1.765 ;
 END
 ANTENNADIFFAREA 0.532 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.72 1.765 20.985 1.905 ;
 RECT 19.72 1.905 19.98 2.12 ;
 RECT 19.785 0.55 19.925 1.765 ;
 RECT 20.845 1.905 20.985 1.93 ;
 RECT 20.845 1.64 20.985 1.765 ;
 END
 ANTENNADIFFAREA 0.499 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.335 2.12 11.67 2.46 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.04 0.41 1.41 0.62 ;
 RECT 1.155 0.62 1.41 0.76 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.985 1.215 2.165 1.425 ;
 RECT 1.795 1.63 2.865 1.79 ;
 RECT 1.795 1.425 2.165 1.63 ;
 RECT 2.715 1.79 2.855 1.845 ;
 RECT 2.715 1.57 2.855 1.63 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.44 1.16 2.715 1.42 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.84 1.435 27.18 1.8 ;
 RECT 25.16 1.99 27.025 2.13 ;
 RECT 22.93 2.22 25.3 2.36 ;
 RECT 25.16 1.435 25.3 1.99 ;
 RECT 26.885 1.8 27.025 1.99 ;
 RECT 22.93 1.39 23.07 2.22 ;
 RECT 24.315 1.37 24.455 2.22 ;
 RECT 25.16 2.13 25.3 2.22 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 21.61 0.59 21.98 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 OBS
 LAYER PO ;
 RECT 23.985 0.935 24.215 0.96 ;
 RECT 23.985 0.96 24.505 1.06 ;
 RECT 23.985 1.06 24.215 1.145 ;
 RECT 24.77 0.22 25 0.28 ;
 RECT 24.77 0.38 25 0.43 ;
 RECT 24.405 0.28 25 0.38 ;
 RECT 26.59 0.195 26.69 2.665 ;
 RECT 25.58 0.095 26.69 0.195 ;
 RECT 21.955 1.245 22.055 2.665 ;
 RECT 21.955 1.2 22.24 1.245 ;
 RECT 25.58 0.195 25.68 0.945 ;
 RECT 22.01 1.035 22.24 1.1 ;
 RECT 21.955 2.665 26.69 2.765 ;
 RECT 21.955 1.1 22.285 1.2 ;
 RECT 23.495 0.215 23.595 0.995 ;
 RECT 23.495 0.995 23.735 1.205 ;
 RECT 23.495 1.205 23.595 2 ;
 RECT 25.89 0.375 25.99 0.99 ;
 RECT 25.89 0.99 26.14 1.2 ;
 RECT 25.89 1.2 25.99 2.27 ;
 RECT 25.89 2.27 26.175 2.48 ;
 RECT 22.715 0.21 22.815 0.755 ;
 RECT 22.715 0.855 22.815 2.2 ;
 RECT 25.58 1.125 25.68 2.2 ;
 RECT 21.75 0.755 23.285 0.84 ;
 RECT 21.75 0.84 23.28 0.855 ;
 RECT 23.185 0.215 23.285 0.755 ;
 RECT 21.75 0.595 21.98 0.755 ;
 RECT 22.715 2.2 25.68 2.3 ;
 RECT 10.58 0.66 10.68 1.13 ;
 RECT 10.58 1.23 10.68 1.655 ;
 RECT 9.665 0.66 9.765 1.13 ;
 RECT 10.58 1.655 11.54 1.755 ;
 RECT 11.44 1.755 11.54 2.25 ;
 RECT 10.58 1.755 10.68 2.57 ;
 RECT 9.665 1.13 10.68 1.23 ;
 RECT 11.44 2.25 11.67 2.46 ;
 RECT 14.115 0.685 14.345 0.875 ;
 RECT 13.445 0.82 13.675 0.875 ;
 RECT 13.445 0.975 13.675 1.03 ;
 RECT 13.445 0.875 14.35 0.975 ;
 RECT 16.83 1.635 16.93 1.66 ;
 RECT 16.83 1.66 17.085 1.87 ;
 RECT 16.83 1.87 16.93 2.565 ;
 RECT 17.49 0.19 17.59 0.22 ;
 RECT 18.435 0.19 18.535 1.435 ;
 RECT 18.435 1.535 18.535 2.26 ;
 RECT 18.905 0.5 19.005 1.435 ;
 RECT 18.905 1.535 19.005 2.26 ;
 RECT 17.49 0.09 18.535 0.19 ;
 RECT 18.43 1.435 19.005 1.535 ;
 RECT 17.36 0.22 17.59 0.43 ;
 RECT 17.105 1.25 17.365 1.3 ;
 RECT 17.265 0.61 17.365 1.25 ;
 RECT 17.105 1.4 17.365 1.46 ;
 RECT 17.265 1.46 17.365 2.56 ;
 RECT 17.795 0.68 17.895 1.3 ;
 RECT 17.105 1.3 17.895 1.4 ;
 RECT 17.78 0.47 18.01 0.68 ;
 RECT 15.505 0.51 15.605 0.53 ;
 RECT 15.505 0.74 15.605 2.21 ;
 RECT 15.465 0.53 15.695 0.74 ;
 RECT 15.035 0.54 15.285 0.695 ;
 RECT 15.035 0.695 15.135 2.21 ;
 RECT 15.055 0.485 15.285 0.54 ;
 RECT 11.87 2.69 13.78 2.695 ;
 RECT 13.68 2.54 13.78 2.69 ;
 RECT 12.66 2.695 13.78 2.79 ;
 RECT 11.87 0.66 11.97 2.595 ;
 RECT 11.87 2.595 12.76 2.69 ;
 RECT 13.68 2.33 13.91 2.54 ;
 RECT 6.415 0.185 13.005 0.19 ;
 RECT 12.905 1.355 14 1.39 ;
 RECT 12.905 0.19 13.005 1.29 ;
 RECT 12.905 1.29 13.995 1.355 ;
 RECT 6.415 0.285 6.515 0.51 ;
 RECT 6.415 0.19 8.25 0.285 ;
 RECT 8.15 0.285 8.25 1.24 ;
 RECT 8.15 0.09 13.005 0.185 ;
 RECT 13.77 1.39 14 1.565 ;
 RECT 6.375 0.51 6.62 0.755 ;
 RECT 13.475 1.71 13.575 1.76 ;
 RECT 9.2 0.48 9.385 0.5 ;
 RECT 16.835 0.19 16.935 1.18 ;
 RECT 14.535 0.19 14.635 1.76 ;
 RECT 13.475 1.76 14.635 1.86 ;
 RECT 12.39 0.48 12.49 1.61 ;
 RECT 12.94 1.71 13.04 2.445 ;
 RECT 14.535 0.09 16.935 0.19 ;
 RECT 12.39 1.61 13.575 1.71 ;
 RECT 9.2 0.38 12.49 0.48 ;
 RECT 9.155 0.5 9.385 0.71 ;
 RECT 9.655 1.575 9.755 2.485 ;
 RECT 10.165 1.41 10.395 1.475 ;
 RECT 10.165 1.575 10.395 1.62 ;
 RECT 9.655 1.475 10.395 1.575 ;
 RECT 2 0.555 2.1 1.215 ;
 RECT 1.96 1.215 2.205 1.455 ;
 RECT 7.41 1.33 7.55 1.475 ;
 RECT 7.41 1.71 7.51 2.475 ;
 RECT 7.45 0.65 7.55 1.33 ;
 RECT 7.41 1.475 7.64 1.71 ;
 RECT 3.105 0.58 3.205 2.79 ;
 RECT 2.9 0.35 3.205 0.58 ;
 RECT 2.665 1.59 2.905 1.82 ;
 RECT 2.805 1.82 2.905 2.79 ;
 RECT 3.575 0.35 3.675 1.2 ;
 RECT 3.575 1.41 3.675 2.79 ;
 RECT 3.395 1.2 3.675 1.41 ;
 RECT 2.385 1.41 2.485 1.645 ;
 RECT 2.61 0.555 2.71 1.18 ;
 RECT 2.335 1.745 2.435 2.79 ;
 RECT 2.335 1.645 2.485 1.745 ;
 RECT 2.385 1.18 2.71 1.41 ;
 RECT 7.85 0.695 7.95 1.61 ;
 RECT 7.885 1.71 7.985 2.48 ;
 RECT 7.85 1.61 7.985 1.71 ;
 RECT 7.73 0.465 7.97 0.695 ;
 RECT 9.015 1.61 9.28 1.82 ;
 RECT 9.18 1.82 9.28 2.49 ;
 RECT 8.81 0.66 8.91 1.51 ;
 RECT 8.81 1.51 9.28 1.61 ;
 RECT 6.915 1.595 7.015 2.48 ;
 RECT 6.375 1.445 6.62 1.495 ;
 RECT 6.375 1.595 6.62 1.69 ;
 RECT 6.375 1.495 7.015 1.595 ;
 RECT 11.475 0.66 11.575 1.24 ;
 RECT 11.345 1.24 11.575 1.475 ;
 RECT 5.255 0.655 5.355 1.495 ;
 RECT 5.06 1.495 5.355 1.745 ;
 RECT 5.255 1.745 5.355 2.37 ;
 RECT 4.78 0.52 4.88 2.465 ;
 RECT 4.54 0.27 4.88 0.52 ;
 RECT 5.595 1.52 6.195 1.62 ;
 RECT 6.96 0.47 7.245 0.705 ;
 RECT 6.96 0.705 7.06 1.165 ;
 RECT 6.095 0.585 6.195 1.165 ;
 RECT 6.095 1.265 6.195 1.52 ;
 RECT 6.03 1.62 6.13 2.69 ;
 RECT 8.71 1.79 8.81 2.69 ;
 RECT 5.595 1.44 5.84 1.52 ;
 RECT 5.595 1.62 5.84 1.69 ;
 RECT 6.095 1.165 7.06 1.265 ;
 RECT 6.03 2.69 8.81 2.79 ;
 RECT 1.195 0.62 1.295 1.195 ;
 RECT 1.195 1.195 1.765 1.295 ;
 RECT 1.195 1.295 1.295 2.745 ;
 RECT 1.665 0.555 1.765 1.195 ;
 RECT 1.665 1.295 1.765 2.79 ;
 RECT 1.04 0.41 1.295 0.62 ;
 RECT 23.19 1.245 23.29 2.02 ;
 RECT 23.06 1.035 23.29 1.245 ;
 RECT 20.045 0.19 20.145 1.2 ;
 RECT 20.045 1.435 20.145 2.555 ;
 RECT 20.625 1.43 20.725 2.565 ;
 RECT 20.03 1.2 20.24 1.33 ;
 RECT 20.03 1.43 20.24 1.435 ;
 RECT 20.03 1.33 20.725 1.43 ;
 RECT 21.17 0.19 21.27 0.22 ;
 RECT 20.045 0.09 21.27 0.19 ;
 RECT 21.17 0.22 21.4 0.43 ;
 RECT 24.405 1.06 24.505 1.14 ;
 RECT 24.405 0.38 24.505 0.96 ;
 RECT 24.405 1.14 24.675 1.24 ;
 RECT 24.575 1.24 24.675 1.84 ;
 LAYER CO ;
 RECT 2.36 0.79 2.49 0.92 ;
 RECT 0.81 0.79 0.94 0.92 ;
 RECT 20.85 1.71 20.98 1.84 ;
 RECT 20.265 2.64 20.395 2.77 ;
 RECT 19.79 1.725 19.92 1.855 ;
 RECT 6.25 1.825 6.38 1.955 ;
 RECT 11.395 1.28 11.525 1.41 ;
 RECT 9.4 2.015 9.53 2.145 ;
 RECT 0.3 2.085 0.43 2.215 ;
 RECT 10.33 0.88 10.46 1.01 ;
 RECT 12.13 1.945 12.26 2.075 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 11.22 0.62 11.35 0.75 ;
 RECT 0.3 2.345 0.43 2.475 ;
 RECT 7.785 0.515 7.915 0.645 ;
 RECT 7.16 2.07 7.29 2.2 ;
 RECT 5 0.875 5.13 1.005 ;
 RECT 8.39 0.455 8.52 0.585 ;
 RECT 6.43 1.49 6.56 1.62 ;
 RECT 6.43 0.555 6.56 0.685 ;
 RECT 7.18 0.88 7.31 1.01 ;
 RECT 4.6 0.325 4.73 0.455 ;
 RECT 4.53 0.875 4.66 1.005 ;
 RECT 8.93 2.135 9.06 2.265 ;
 RECT 5.74 2.345 5.87 2.475 ;
 RECT 9.885 2.07 10.015 2.2 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 4.53 2.115 4.66 2.245 ;
 RECT 7.63 2.125 7.76 2.255 ;
 RECT 6.315 0.905 6.445 1.035 ;
 RECT 6.665 2.105 6.795 2.235 ;
 RECT 5.605 0.875 5.735 1.005 ;
 RECT 5 2.05 5.13 2.18 ;
 RECT 8.11 1.825 8.24 1.955 ;
 RECT 5.12 1.55 5.25 1.68 ;
 RECT 1.09 0.45 1.22 0.58 ;
 RECT 23.11 1.075 23.24 1.205 ;
 RECT 25.96 1.03 26.09 1.16 ;
 RECT 21.22 0.26 21.35 0.39 ;
 RECT 24.035 0.975 24.165 1.105 ;
 RECT 24.82 0.26 24.95 0.39 ;
 RECT 22.06 1.075 22.19 1.205 ;
 RECT 23.555 1.035 23.685 1.165 ;
 RECT 25.995 2.31 26.125 2.44 ;
 RECT 21.8 0.635 21.93 0.765 ;
 RECT 11.49 2.29 11.62 2.42 ;
 RECT 14.165 0.725 14.295 0.855 ;
 RECT 13.495 0.86 13.625 0.99 ;
 RECT 17.83 0.51 17.96 0.64 ;
 RECT 16.905 1.7 17.035 1.83 ;
 RECT 17.41 0.26 17.54 0.39 ;
 RECT 17.155 1.29 17.285 1.42 ;
 RECT 15.515 0.57 15.645 0.7 ;
 RECT 15.105 0.525 15.235 0.655 ;
 RECT 13.73 2.37 13.86 2.5 ;
 RECT 13.82 1.395 13.95 1.525 ;
 RECT 9.205 0.54 9.335 0.67 ;
 RECT 10.215 1.45 10.345 1.58 ;
 RECT 20.07 1.25 20.2 1.38 ;
 RECT 20.35 0.62 20.48 0.75 ;
 RECT 2.02 1.265 2.15 1.395 ;
 RECT 3.795 0.79 3.925 0.92 ;
 RECT 1.415 0.12 1.545 0.25 ;
 RECT 1.415 2.055 1.545 2.185 ;
 RECT 1.415 2.315 1.545 2.445 ;
 RECT 3.795 2.05 3.925 2.18 ;
 RECT 3.325 2.35 3.455 2.48 ;
 RECT 2.53 1.23 2.66 1.36 ;
 RECT 17.485 0.83 17.615 0.96 ;
 RECT 16.585 0.33 16.715 0.46 ;
 RECT 17.485 1.78 17.615 1.91 ;
 RECT 16.58 2.64 16.71 2.77 ;
 RECT 14.78 0.3 14.91 0.43 ;
 RECT 15.725 0.975 15.855 1.105 ;
 RECT 15.725 1.705 15.855 1.835 ;
 RECT 15.255 2.64 15.385 2.77 ;
 RECT 14.785 1.7 14.915 1.83 ;
 RECT 11.03 2.445 11.16 2.575 ;
 RECT 24.795 1.405 24.925 1.535 ;
 RECT 22.215 0.505 22.345 0.635 ;
 RECT 23.715 1.485 23.845 1.615 ;
 RECT 24.15 0.12 24.28 0.25 ;
 RECT 25.165 1.49 25.295 1.62 ;
 RECT 22.935 1.475 23.065 1.605 ;
 RECT 24.32 1.445 24.45 1.575 ;
 RECT 25.33 0.12 25.46 0.25 ;
 RECT 26.11 1.465 26.24 1.595 ;
 RECT 22.935 0.135 23.065 0.265 ;
 RECT 26.89 1.475 27.02 1.605 ;
 RECT 23.715 0.435 23.845 0.565 ;
 RECT 26.11 0.595 26.24 0.725 ;
 RECT 22.465 1.425 22.595 1.555 ;
 RECT 24.655 0.595 24.785 0.725 ;
 RECT 5.745 0.21 5.875 0.34 ;
 RECT 0.3 1.825 0.43 1.955 ;
 RECT 8.46 2.125 8.59 2.255 ;
 RECT 5.475 1.995 5.605 2.125 ;
 RECT 7.46 1.525 7.59 1.655 ;
 RECT 6.71 0.88 6.84 1.01 ;
 RECT 9.4 0.93 9.53 1.06 ;
 RECT 7.065 0.525 7.195 0.655 ;
 RECT 10.33 1.995 10.46 2.125 ;
 RECT 9.885 0.88 10.015 1.01 ;
 RECT 5.655 1.495 5.785 1.625 ;
 RECT 12.13 0.88 12.26 1.01 ;
 RECT 9.07 1.63 9.2 1.76 ;
 RECT 18.655 0.34 18.785 0.47 ;
 RECT 18.675 2.64 18.805 2.77 ;
 RECT 19.125 1.705 19.255 1.835 ;
 RECT 19.125 0.975 19.255 1.105 ;
 RECT 18.185 0.975 18.315 1.105 ;
 RECT 13.16 0.595 13.29 0.725 ;
 RECT 13.16 1.87 13.29 2 ;
 RECT 12.655 0.595 12.785 0.725 ;
 RECT 12.655 1.9 12.785 2.03 ;
 RECT 18.185 1.705 18.315 1.835 ;
 RECT 19.79 0.625 19.92 0.755 ;
 RECT 3.795 1.79 3.925 1.92 ;
 RECT 3.325 0.6 3.455 0.73 ;
 RECT 3.445 1.24 3.575 1.37 ;
 RECT 2.555 2.115 2.685 2.245 ;
 RECT 3.325 2.09 3.455 2.22 ;
 RECT 2.72 1.64 2.85 1.77 ;
 RECT 0.945 2.055 1.075 2.185 ;
 RECT 2.95 0.4 3.08 0.53 ;
 LAYER M1 ;
 RECT 10.325 1.62 10.465 2.18 ;
 RECT 11.075 1.275 11.595 1.415 ;
 RECT 3.01 0.925 3.15 1.245 ;
 RECT 3.01 1.385 3.15 2.11 ;
 RECT 2.285 0.785 3.15 0.925 ;
 RECT 2.5 2.11 3.15 2.25 ;
 RECT 3.01 1.245 3.58 1.385 ;
 RECT 3.44 1.19 3.58 1.245 ;
 RECT 3.44 1.385 3.58 1.42 ;
 RECT 5.515 1.63 5.655 1.99 ;
 RECT 5.515 1.475 5.86 1.63 ;
 RECT 5.6 0.825 5.74 1.475 ;
 RECT 5.405 1.99 5.655 2.13 ;
 RECT 24.65 0.73 24.79 1.04 ;
 RECT 24.79 1.18 24.93 1.605 ;
 RECT 24.585 0.59 24.86 0.73 ;
 RECT 25.91 0.99 26.14 1.04 ;
 RECT 24.65 1.04 26.14 1.18 ;
 RECT 25.91 1.18 26.14 1.2 ;
 RECT 24.77 0.29 25.14 0.43 ;
 RECT 25 0.43 25.14 0.71 ;
 RECT 24.77 0.22 25 0.29 ;
 RECT 26.42 0.85 26.56 1.385 ;
 RECT 26.105 1.525 26.245 1.73 ;
 RECT 25 0.71 26.56 0.85 ;
 RECT 26.105 0.51 26.245 0.71 ;
 RECT 26.105 1.385 26.56 1.525 ;
 RECT 22.01 1.225 22.24 1.245 ;
 RECT 22.01 1.195 22.6 1.225 ;
 RECT 22.15 1.015 22.46 1.035 ;
 RECT 22.01 1.035 22.46 1.055 ;
 RECT 22.285 0.64 22.425 1.015 ;
 RECT 22.46 1.225 22.6 1.75 ;
 RECT 22.165 0.5 22.425 0.64 ;
 RECT 23.06 1.035 23.29 1.055 ;
 RECT 23.06 1.195 23.29 1.245 ;
 RECT 22.01 1.055 23.29 1.195 ;
 RECT 24.03 1.145 24.17 1.345 ;
 RECT 23.71 1.485 23.85 1.76 ;
 RECT 24.03 0.73 24.17 0.935 ;
 RECT 23.71 0.355 23.85 0.59 ;
 RECT 23.71 1.345 24.17 1.485 ;
 RECT 23.985 0.935 24.215 1.145 ;
 RECT 23.71 0.59 24.17 0.73 ;
 RECT 21.17 0.36 21.4 0.43 ;
 RECT 22.565 0.36 22.705 0.565 ;
 RECT 21.17 0.22 22.705 0.36 ;
 RECT 23.305 0.705 23.445 0.75 ;
 RECT 23.43 0.995 23.735 1.205 ;
 RECT 23.43 0.89 23.57 0.995 ;
 RECT 23.305 0.75 23.57 0.89 ;
 RECT 22.565 0.565 23.445 0.705 ;
 RECT 17.78 0.475 18.385 0.625 ;
 RECT 17.78 0.47 18.01 0.475 ;
 RECT 17.78 0.635 18.01 0.68 ;
 RECT 19.165 0.37 19.305 0.625 ;
 RECT 17.78 0.625 19.305 0.635 ;
 RECT 18.245 0.635 19.305 0.765 ;
 RECT 19.165 0.765 19.305 0.77 ;
 RECT 20.065 0.37 20.205 1.46 ;
 RECT 19.165 0.23 20.205 0.37 ;
 RECT 13.445 0.82 13.675 0.855 ;
 RECT 13.445 0.995 13.675 1.03 ;
 RECT 13.155 0.525 13.295 0.855 ;
 RECT 13.155 0.995 13.295 2.065 ;
 RECT 13.155 0.855 13.675 0.995 ;
 RECT 10.73 1.875 10.87 2.33 ;
 RECT 10.73 2.47 10.87 2.475 ;
 RECT 9.88 2.33 10.87 2.47 ;
 RECT 9.88 0.82 10.02 2.33 ;
 RECT 9.88 2.47 10.02 2.475 ;
 RECT 11.81 1.875 11.95 2.295 ;
 RECT 12.125 0.765 12.265 2.295 ;
 RECT 12.65 0.525 12.79 2.295 ;
 RECT 10.73 1.735 11.95 1.875 ;
 RECT 11.81 2.295 12.79 2.435 ;
 RECT 15.055 0.36 15.285 0.68 ;
 RECT 14.12 0.68 15.285 0.685 ;
 RECT 14.12 0.895 15.285 0.91 ;
 RECT 14.115 0.685 15.285 0.895 ;
 RECT 15.055 0.22 16.435 0.36 ;
 RECT 16.295 0.36 16.435 0.675 ;
 RECT 16.295 0.675 17.62 0.815 ;
 RECT 17.36 0.23 17.62 0.43 ;
 RECT 17.36 0.22 17.59 0.23 ;
 RECT 17.48 0.43 17.62 0.675 ;
 RECT 17.48 0.815 17.62 1.98 ;
 RECT 6.31 0.5 6.565 0.965 ;
 RECT 6.31 0.965 6.45 1.44 ;
 RECT 6.31 1.44 6.565 1.67 ;
 RECT 6.31 1.67 6.45 1.82 ;
 RECT 6.18 1.82 6.45 1.96 ;
 RECT 6.995 0.52 7.64 0.66 ;
 RECT 7.5 0.66 7.64 1.015 ;
 RECT 9 0.505 9.385 0.71 ;
 RECT 7.5 1.015 9.14 1.155 ;
 RECT 9 0.71 9.14 1.015 ;
 RECT 9.155 0.5 9.385 0.505 ;
 RECT 4.305 1.01 4.445 1.195 ;
 RECT 4.305 1.335 4.445 2.11 ;
 RECT 4.305 2.25 4.445 2.255 ;
 RECT 4.305 0.87 4.73 1.01 ;
 RECT 4.305 2.11 4.73 2.25 ;
 RECT 4.305 1.195 5.415 1.335 ;
 RECT 5.275 0.67 5.415 1.195 ;
 RECT 6.705 0.36 6.845 2.035 ;
 RECT 6.02 0.22 6.845 0.36 ;
 RECT 5.275 0.53 6.16 0.67 ;
 RECT 6.66 2.17 6.8 2.305 ;
 RECT 6.66 2.035 6.845 2.17 ;
 RECT 6.02 0.36 6.16 0.53 ;
 RECT 3.79 0.5 3.93 2.25 ;
 RECT 3.79 0.36 4.855 0.5 ;
 RECT 4.49 0.22 4.855 0.36 ;
 RECT 4.49 0.5 4.855 0.615 ;
 RECT 1.705 0.535 1.845 1.14 ;
 RECT 0.805 1.14 1.845 1.28 ;
 RECT 0.94 1.28 1.08 2.27 ;
 RECT 0.805 0.925 0.945 1.14 ;
 RECT 0.74 0.785 0.99 0.925 ;
 RECT 1.705 0.395 3.15 0.535 ;
 RECT 13.68 2.42 13.91 2.54 ;
 RECT 21.16 2.42 21.3 2.52 ;
 RECT 13.68 2.28 21.3 2.42 ;
 RECT 25.945 2.48 26.085 2.52 ;
 RECT 25.945 2.27 26.175 2.48 ;
 RECT 21.16 2.52 26.085 2.66 ;
 RECT 14.78 1.51 14.92 1.695 ;
 RECT 14.71 1.695 14.99 1.835 ;
 RECT 15.72 0.905 15.86 1.37 ;
 RECT 15.72 1.51 15.86 1.7 ;
 RECT 17.105 1.25 17.335 1.37 ;
 RECT 14.78 1.37 17.335 1.51 ;
 RECT 15.655 1.7 15.93 1.84 ;
 RECT 13.815 1.565 13.955 1.985 ;
 RECT 13.815 1.985 17.085 2.125 ;
 RECT 16.855 1.66 17.085 1.985 ;
 RECT 13.77 1.355 14 1.565 ;
 RECT 8.12 1.44 8.26 1.52 ;
 RECT 7.39 1.52 8.26 1.66 ;
 RECT 9.395 0.865 9.535 1.3 ;
 RECT 8.12 1.3 9.535 1.44 ;
 RECT 9.395 1.44 9.535 2.215 ;
 RECT 7.56 2.12 8.66 2.26 ;
 RECT 7 1.22 7.315 1.36 ;
 RECT 7.175 0.805 7.315 1.22 ;
 RECT 7.085 1.96 7.365 2.215 ;
 RECT 7 1.36 7.14 1.82 ;
 RECT 7 1.82 8.58 1.96 ;
 RECT 8.44 1.79 8.58 1.82 ;
 RECT 9.015 1.58 9.255 1.65 ;
 RECT 8.44 1.65 9.255 1.79 ;
 RECT 9.015 1.79 9.255 1.835 ;
 RECT 11.075 1.415 11.215 1.455 ;
 RECT 10.165 1.455 11.215 1.595 ;
 RECT 10.165 1.41 10.465 1.455 ;
 RECT 10.325 0.81 10.465 1.41 ;
 RECT 10.165 1.595 10.465 1.62 ;
 END
END RSDFFSRARX1

MACRO RSDFFSRARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 30.72 BY 2.88 ;
 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.78 0.735 8.855 0.875 ;
 RECT 11.59 0.245 13.96 0.385 ;
 RECT 7.78 0.445 8.11 0.735 ;
 RECT 8.715 0.36 8.855 0.735 ;
 RECT 10.615 0.99 11.73 1.13 ;
 RECT 13.82 1.05 15.57 1.19 ;
 RECT 15.43 0.74 15.57 1.05 ;
 RECT 15.465 0.53 15.695 0.555 ;
 RECT 15.43 0.555 15.695 0.74 ;
 RECT 10.615 0.36 10.755 0.99 ;
 RECT 8.715 0.22 10.755 0.36 ;
 RECT 11.59 0.385 11.73 0.99 ;
 RECT 13.82 0.385 13.96 1.05 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 30.72 0.08 ;
 RECT 27.39 0.08 27.63 0.26 ;
 RECT 18.8 0.35 19.065 0.49 ;
 RECT 19.74 0.35 20.045 0.49 ;
 RECT 1.41 0.08 1.55 1.045 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.995 0.08 5.135 1.055 ;
 RECT 3.32 0.08 3.46 0.85 ;
 RECT 5.74 0.08 5.88 0.39 ;
 RECT 8.34 0.08 8.575 0.595 ;
 RECT 11.215 0.08 11.355 0.815 ;
 RECT 14.775 0.08 14.915 0.5 ;
 RECT 16.58 0.08 16.72 0.525 ;
 RECT 25.04 0.08 25.18 0.36 ;
 RECT 21.52 0.08 21.66 0.82 ;
 RECT 26.255 0.08 26.395 0.35 ;
 RECT 18.875 0.08 19.015 0.35 ;
 RECT 19.825 0.08 19.965 0.35 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 30.72 2.96 ;
 RECT 1.41 2.005 1.55 2.8 ;
 RECT 0.295 1.74 0.435 2.8 ;
 RECT 5.67 2.34 5.92 2.8 ;
 RECT 3.32 2.03 3.46 2.8 ;
 RECT 4.995 1.98 5.135 2.8 ;
 RECT 11.025 2.375 11.165 2.8 ;
 RECT 8.925 2.07 9.065 2.8 ;
 RECT 15.25 2.57 15.39 2.8 ;
 RECT 18.845 2.57 18.985 2.8 ;
 RECT 16.575 2.57 16.715 2.8 ;
 RECT 19.845 2.57 19.985 2.8 ;
 RECT 21.435 2.57 21.575 2.8 ;
 RECT 22.49 2.57 22.63 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.985 1.475 5.375 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.395 1.765 20.605 1.905 ;
 RECT 20.295 1.905 20.605 2.04 ;
 RECT 20.295 0.915 20.435 1.765 ;
 RECT 18.395 0.915 18.535 1.765 ;
 RECT 19.355 0.915 19.495 1.765 ;
 END
 ANTENNADIFFAREA 0.788 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.96 1.765 23.1 1.905 ;
 RECT 20.68 0.84 21.1 1.085 ;
 RECT 20.96 0.55 21.1 0.84 ;
 RECT 22.96 1.905 23.1 1.97 ;
 RECT 22.96 1.7 23.1 1.765 ;
 RECT 22.02 1.905 22.16 1.91 ;
 RECT 22.02 0.56 22.16 1.765 ;
 RECT 20.96 1.905 21.1 1.925 ;
 RECT 20.96 1.085 21.1 1.765 ;
 END
 ANTENNADIFFAREA 0.942 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.335 2.12 11.67 2.495 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.23 1.475 1.755 1.75 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.015 1.79 2.36 2.04 ;
 RECT 2.715 1.79 2.855 1.845 ;
 RECT 2.715 1.57 2.855 1.63 ;
 RECT 2.015 1.175 2.155 1.63 ;
 RECT 2.015 1.63 2.865 1.79 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.38 1.135 2.74 1.4 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 28.95 1.435 29.29 1.8 ;
 RECT 27.27 1.99 29.135 2.13 ;
 RECT 25.04 2.22 27.41 2.36 ;
 RECT 28.995 1.8 29.135 1.99 ;
 RECT 27.27 1.435 27.41 1.99 ;
 RECT 25.04 1.39 25.18 2.22 ;
 RECT 26.425 1.37 26.565 2.22 ;
 RECT 27.27 2.13 27.41 2.22 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 23.72 0.59 24.09 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 OBS
 LAYER PO ;
 RECT 26.095 1.06 26.325 1.145 ;
 RECT 26.515 1.14 26.785 1.24 ;
 RECT 26.685 1.24 26.785 1.84 ;
 RECT 26.88 0.22 27.11 0.28 ;
 RECT 26.88 0.38 27.11 0.43 ;
 RECT 26.515 0.28 27.11 0.38 ;
 RECT 28.7 0.195 28.8 2.665 ;
 RECT 27.69 0.095 28.8 0.195 ;
 RECT 24.065 1.245 24.165 2.665 ;
 RECT 24.065 1.2 24.35 1.245 ;
 RECT 27.69 0.195 27.79 0.945 ;
 RECT 24.12 1.035 24.35 1.1 ;
 RECT 24.065 2.665 28.8 2.765 ;
 RECT 24.065 1.1 24.395 1.2 ;
 RECT 25.605 0.215 25.705 0.995 ;
 RECT 25.605 0.995 25.845 1.205 ;
 RECT 25.605 1.205 25.705 2 ;
 RECT 28 0.375 28.1 0.99 ;
 RECT 28 0.99 28.25 1.2 ;
 RECT 28 1.2 28.1 2.27 ;
 RECT 28 2.27 28.285 2.48 ;
 RECT 24.825 0.855 24.925 2.2 ;
 RECT 27.69 1.125 27.79 2.2 ;
 RECT 23.86 0.755 25.395 0.84 ;
 RECT 23.86 0.84 25.39 0.855 ;
 RECT 25.295 0.215 25.395 0.755 ;
 RECT 24.825 0.21 24.925 0.755 ;
 RECT 23.86 0.595 24.09 0.755 ;
 RECT 24.825 2.2 27.79 2.3 ;
 RECT 10.58 0.66 10.68 1.13 ;
 RECT 10.58 1.23 10.68 1.655 ;
 RECT 9.665 0.66 9.765 1.13 ;
 RECT 10.58 1.655 11.54 1.755 ;
 RECT 11.44 1.755 11.54 2.285 ;
 RECT 10.58 1.755 10.68 2.57 ;
 RECT 9.665 1.13 10.68 1.23 ;
 RECT 11.44 2.285 11.67 2.495 ;
 RECT 14.115 0.685 14.345 0.875 ;
 RECT 13.445 0.82 13.675 0.875 ;
 RECT 13.445 0.975 13.675 1.03 ;
 RECT 13.445 0.875 14.35 0.975 ;
 RECT 16.83 1.635 16.93 1.66 ;
 RECT 16.83 1.66 17.085 1.87 ;
 RECT 16.83 1.87 16.93 2.565 ;
 RECT 18.66 0.19 18.76 1.435 ;
 RECT 17.49 0.19 17.59 0.22 ;
 RECT 19.14 0.56 19.24 1.435 ;
 RECT 20.08 0.555 20.18 1.435 ;
 RECT 20.08 1.535 20.18 2.21 ;
 RECT 19.61 0.555 19.71 1.435 ;
 RECT 19.61 1.535 19.71 2.205 ;
 RECT 19.14 1.535 19.24 2.205 ;
 RECT 18.66 1.535 18.76 2.215 ;
 RECT 17.49 0.09 18.76 0.19 ;
 RECT 18.66 1.435 20.18 1.535 ;
 RECT 17.36 0.22 17.59 0.43 ;
 RECT 17.105 1.25 17.365 1.3 ;
 RECT 17.265 0.61 17.365 1.25 ;
 RECT 17.105 1.4 17.365 1.46 ;
 RECT 17.265 1.46 17.365 2.56 ;
 RECT 17.795 0.84 17.895 1.3 ;
 RECT 17.105 1.3 17.895 1.4 ;
 RECT 17.78 0.63 18.01 0.84 ;
 RECT 15.505 0.51 15.605 0.53 ;
 RECT 15.505 0.74 15.605 2.21 ;
 RECT 15.465 0.53 15.695 0.74 ;
 RECT 15.035 0.54 15.285 0.695 ;
 RECT 15.035 0.695 15.135 2.21 ;
 RECT 15.055 0.485 15.285 0.54 ;
 RECT 11.87 2.69 13.78 2.695 ;
 RECT 13.68 2.54 13.78 2.69 ;
 RECT 12.66 2.695 13.78 2.79 ;
 RECT 11.87 0.66 11.97 2.595 ;
 RECT 11.87 2.595 12.76 2.69 ;
 RECT 13.68 2.33 13.91 2.54 ;
 RECT 6.415 0.185 13.005 0.19 ;
 RECT 12.905 1.355 14 1.39 ;
 RECT 12.905 0.19 13.005 1.29 ;
 RECT 12.905 1.29 13.995 1.355 ;
 RECT 6.415 0.285 6.515 0.51 ;
 RECT 6.415 0.19 8.25 0.285 ;
 RECT 8.15 0.285 8.25 1.24 ;
 RECT 8.15 0.09 13.005 0.185 ;
 RECT 13.77 1.39 14 1.565 ;
 RECT 6.375 0.51 6.62 0.755 ;
 RECT 13.475 1.71 13.575 1.76 ;
 RECT 9.2 0.48 9.385 0.5 ;
 RECT 16.835 0.19 16.935 1.18 ;
 RECT 14.535 0.19 14.635 1.76 ;
 RECT 13.475 1.76 14.635 1.86 ;
 RECT 12.39 0.48 12.49 1.61 ;
 RECT 12.94 1.71 13.04 2.445 ;
 RECT 14.535 0.09 16.935 0.19 ;
 RECT 12.39 1.61 13.575 1.71 ;
 RECT 9.2 0.38 12.49 0.48 ;
 RECT 9.155 0.5 9.385 0.71 ;
 RECT 9.655 1.575 9.755 2.485 ;
 RECT 10.165 1.41 10.395 1.475 ;
 RECT 10.165 1.575 10.395 1.62 ;
 RECT 9.655 1.475 10.395 1.575 ;
 RECT 1.195 1.475 1.765 1.75 ;
 RECT 1.665 0.555 1.765 1.475 ;
 RECT 1.665 1.75 1.765 2.79 ;
 RECT 1.195 0.555 1.295 1.475 ;
 RECT 1.195 1.75 1.295 2.745 ;
 RECT 2 0.555 2.1 1.225 ;
 RECT 1.96 1.225 2.205 1.465 ;
 RECT 3.105 0.57 3.205 2.79 ;
 RECT 2.9 0.34 3.205 0.57 ;
 RECT 2.665 1.59 2.905 1.82 ;
 RECT 2.805 1.82 2.905 2.79 ;
 RECT 3.575 0.35 3.675 1.2 ;
 RECT 3.575 1.41 3.675 2.79 ;
 RECT 3.395 1.2 3.675 1.41 ;
 RECT 2.385 1.41 2.485 1.645 ;
 RECT 2.61 0.555 2.71 1.18 ;
 RECT 2.335 1.745 2.435 2.79 ;
 RECT 2.335 1.645 2.485 1.745 ;
 RECT 2.385 1.18 2.715 1.41 ;
 RECT 7.85 0.695 7.95 1.61 ;
 RECT 7.885 1.71 7.985 2.48 ;
 RECT 7.85 1.61 7.985 1.71 ;
 RECT 7.73 0.465 7.97 0.695 ;
 RECT 9.015 1.61 9.28 1.82 ;
 RECT 9.18 1.82 9.28 2.49 ;
 RECT 8.81 0.66 8.91 1.51 ;
 RECT 8.81 1.51 9.28 1.61 ;
 RECT 6.915 1.595 7.015 2.48 ;
 RECT 6.375 1.445 6.62 1.495 ;
 RECT 6.375 1.595 6.62 1.69 ;
 RECT 6.375 1.495 7.015 1.595 ;
 RECT 11.475 0.66 11.575 1.24 ;
 RECT 11.345 1.24 11.575 1.475 ;
 RECT 5.255 0.655 5.355 1.495 ;
 RECT 5.06 1.495 5.355 1.745 ;
 RECT 5.255 1.745 5.355 2.37 ;
 RECT 4.78 0.52 4.88 2.465 ;
 RECT 4.54 0.27 4.88 0.52 ;
 RECT 7.41 1.33 7.55 1.475 ;
 RECT 7.41 1.71 7.51 2.475 ;
 RECT 7.45 0.65 7.55 1.33 ;
 RECT 7.41 1.475 7.64 1.71 ;
 RECT 6.095 1.265 6.195 1.52 ;
 RECT 5.595 1.52 6.195 1.62 ;
 RECT 6.03 1.62 6.13 2.69 ;
 RECT 8.71 1.79 8.81 2.69 ;
 RECT 5.595 1.44 5.84 1.52 ;
 RECT 5.595 1.62 5.84 1.69 ;
 RECT 6.96 0.705 7.06 1.165 ;
 RECT 6.095 0.585 6.195 1.165 ;
 RECT 6.96 0.47 7.245 0.705 ;
 RECT 6.03 2.69 8.81 2.79 ;
 RECT 6.095 1.165 7.06 1.265 ;
 RECT 25.3 1.245 25.4 2.02 ;
 RECT 25.17 1.035 25.4 1.245 ;
 RECT 21.22 0.385 21.32 1.2 ;
 RECT 21.8 0.19 21.9 1.33 ;
 RECT 21.205 1.2 21.415 1.33 ;
 RECT 21.205 1.43 21.415 1.435 ;
 RECT 21.205 1.33 22.845 1.43 ;
 RECT 21.22 1.435 21.32 2.555 ;
 RECT 22.745 1.43 22.845 2.555 ;
 RECT 22.275 1.43 22.375 2.555 ;
 RECT 21.8 1.43 21.9 2.565 ;
 RECT 23.28 0.19 23.38 0.22 ;
 RECT 21.8 0.09 23.38 0.19 ;
 RECT 23.28 0.22 23.51 0.43 ;
 RECT 26.515 0.38 26.615 0.96 ;
 RECT 26.515 1.06 26.615 1.14 ;
 RECT 26.095 0.935 26.325 0.96 ;
 RECT 26.095 0.96 26.615 1.06 ;
 LAYER CO ;
 RECT 9.4 2.015 9.53 2.145 ;
 RECT 0.3 2.085 0.43 2.215 ;
 RECT 10.33 0.88 10.46 1.01 ;
 RECT 12.13 1.945 12.26 2.075 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 11.22 0.62 11.35 0.75 ;
 RECT 0.3 2.345 0.43 2.475 ;
 RECT 7.785 0.515 7.915 0.645 ;
 RECT 7.16 2.07 7.29 2.2 ;
 RECT 5 0.875 5.13 1.005 ;
 RECT 8.39 0.455 8.52 0.585 ;
 RECT 6.43 1.49 6.56 1.62 ;
 RECT 6.43 0.555 6.56 0.685 ;
 RECT 7.18 0.88 7.31 1.01 ;
 RECT 4.6 0.325 4.73 0.455 ;
 RECT 4.53 0.875 4.66 1.005 ;
 RECT 8.93 2.135 9.06 2.265 ;
 RECT 5.74 2.345 5.87 2.475 ;
 RECT 9.885 2.07 10.015 2.2 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 4.53 2.115 4.66 2.245 ;
 RECT 7.63 2.125 7.76 2.255 ;
 RECT 6.315 0.905 6.445 1.035 ;
 RECT 6.665 2.105 6.795 2.235 ;
 RECT 5.605 0.875 5.735 1.005 ;
 RECT 5 2.05 5.13 2.18 ;
 RECT 8.11 1.825 8.24 1.955 ;
 RECT 5.12 1.55 5.25 1.68 ;
 RECT 5.745 0.21 5.875 0.34 ;
 RECT 0.3 1.825 0.43 1.955 ;
 RECT 8.46 2.125 8.59 2.255 ;
 RECT 5.475 1.995 5.605 2.125 ;
 RECT 7.46 1.525 7.59 1.655 ;
 RECT 6.71 0.88 6.84 1.01 ;
 RECT 25.22 1.075 25.35 1.205 ;
 RECT 28.07 1.03 28.2 1.16 ;
 RECT 23.33 0.26 23.46 0.39 ;
 RECT 26.145 0.975 26.275 1.105 ;
 RECT 26.93 0.26 27.06 0.39 ;
 RECT 24.17 1.075 24.3 1.205 ;
 RECT 25.665 1.035 25.795 1.165 ;
 RECT 28.105 2.31 28.235 2.44 ;
 RECT 23.91 0.635 24.04 0.765 ;
 RECT 11.49 2.325 11.62 2.455 ;
 RECT 14.165 0.725 14.295 0.855 ;
 RECT 13.495 0.86 13.625 0.99 ;
 RECT 17.83 0.67 17.96 0.8 ;
 RECT 16.905 1.7 17.035 1.83 ;
 RECT 17.41 0.26 17.54 0.39 ;
 RECT 17.155 1.29 17.285 1.42 ;
 RECT 15.515 0.57 15.645 0.7 ;
 RECT 15.105 0.525 15.235 0.655 ;
 RECT 13.73 2.37 13.86 2.5 ;
 RECT 13.82 1.395 13.95 1.525 ;
 RECT 9.205 0.54 9.335 0.67 ;
 RECT 10.215 1.45 10.345 1.58 ;
 RECT 2.02 1.275 2.15 1.405 ;
 RECT 3.795 0.79 3.925 0.92 ;
 RECT 1.42 1.55 1.55 1.68 ;
 RECT 1.415 0.79 1.545 0.92 ;
 RECT 1.415 2.055 1.545 2.185 ;
 RECT 1.415 2.315 1.545 2.445 ;
 RECT 3.795 2.05 3.925 2.18 ;
 RECT 3.325 2.35 3.455 2.48 ;
 RECT 2.54 1.23 2.67 1.36 ;
 RECT 17.485 0.83 17.615 0.96 ;
 RECT 16.585 0.33 16.715 0.46 ;
 RECT 17.485 1.78 17.615 1.91 ;
 RECT 16.58 2.64 16.71 2.77 ;
 RECT 14.78 0.3 14.91 0.43 ;
 RECT 15.725 0.975 15.855 1.105 ;
 RECT 15.725 1.705 15.855 1.835 ;
 RECT 15.255 2.64 15.385 2.77 ;
 RECT 14.785 1.7 14.915 1.83 ;
 RECT 11.03 2.445 11.16 2.575 ;
 RECT 26.905 1.405 27.035 1.535 ;
 RECT 24.325 0.505 24.455 0.635 ;
 RECT 25.825 1.485 25.955 1.615 ;
 RECT 26.26 0.12 26.39 0.25 ;
 RECT 27.275 1.49 27.405 1.62 ;
 RECT 25.045 1.475 25.175 1.605 ;
 RECT 26.43 1.445 26.56 1.575 ;
 RECT 27.44 0.12 27.57 0.25 ;
 RECT 28.22 1.465 28.35 1.595 ;
 RECT 25.045 0.135 25.175 0.265 ;
 RECT 29 1.475 29.13 1.605 ;
 RECT 25.825 0.435 25.955 0.565 ;
 RECT 28.22 0.595 28.35 0.725 ;
 RECT 24.575 1.425 24.705 1.555 ;
 RECT 26.765 0.595 26.895 0.725 ;
 RECT 9.4 0.93 9.53 1.06 ;
 RECT 7.065 0.525 7.195 0.655 ;
 RECT 10.33 1.995 10.46 2.125 ;
 RECT 9.885 0.88 10.015 1.01 ;
 RECT 5.655 1.495 5.785 1.625 ;
 RECT 12.13 0.88 12.26 1.01 ;
 RECT 9.07 1.63 9.2 1.76 ;
 RECT 22.495 2.64 22.625 2.77 ;
 RECT 22.965 1.77 23.095 1.9 ;
 RECT 19.83 0.355 19.96 0.485 ;
 RECT 19.85 2.64 19.98 2.77 ;
 RECT 20.3 1.705 20.43 1.835 ;
 RECT 20.3 0.975 20.43 1.105 ;
 RECT 19.36 0.975 19.49 1.105 ;
 RECT 18.88 0.355 19.01 0.485 ;
 RECT 18.4 0.975 18.53 1.105 ;
 RECT 13.16 0.595 13.29 0.725 ;
 RECT 13.16 1.87 13.29 2 ;
 RECT 12.655 0.595 12.785 0.725 ;
 RECT 12.655 1.9 12.785 2.03 ;
 RECT 19.36 1.705 19.49 1.835 ;
 RECT 20.965 0.625 21.095 0.755 ;
 RECT 3.795 1.79 3.925 1.92 ;
 RECT 3.325 0.6 3.455 0.73 ;
 RECT 3.445 1.24 3.575 1.37 ;
 RECT 2.555 2.115 2.685 2.245 ;
 RECT 3.325 2.09 3.455 2.22 ;
 RECT 2.72 1.64 2.85 1.77 ;
 RECT 0.945 2.055 1.075 2.185 ;
 RECT 2.95 0.39 3.08 0.52 ;
 RECT 2.36 0.79 2.49 0.92 ;
 RECT 0.945 0.79 1.075 0.92 ;
 RECT 22.025 0.63 22.155 0.76 ;
 RECT 22.025 1.71 22.155 1.84 ;
 RECT 21.44 2.64 21.57 2.77 ;
 RECT 18.85 2.64 18.98 2.77 ;
 RECT 18.4 1.705 18.53 1.835 ;
 RECT 20.965 1.725 21.095 1.855 ;
 RECT 21.245 1.25 21.375 1.38 ;
 RECT 21.525 0.62 21.655 0.75 ;
 RECT 6.25 1.825 6.38 1.955 ;
 RECT 11.395 1.28 11.525 1.41 ;
 LAYER M1 ;
 RECT 7.56 2.12 8.66 2.26 ;
 RECT 10.73 1.875 10.87 2.33 ;
 RECT 10.73 2.47 10.87 2.475 ;
 RECT 9.88 2.33 10.87 2.47 ;
 RECT 9.88 0.82 10.02 2.33 ;
 RECT 9.88 2.47 10.02 2.475 ;
 RECT 11.81 1.875 11.95 2.295 ;
 RECT 12.65 0.525 12.79 2.295 ;
 RECT 12.125 0.765 12.265 2.295 ;
 RECT 11.81 2.295 12.79 2.435 ;
 RECT 10.73 1.735 11.95 1.875 ;
 RECT 7 1.22 7.315 1.36 ;
 RECT 7.175 0.805 7.315 1.22 ;
 RECT 7.085 1.96 7.365 2.215 ;
 RECT 7 1.36 7.14 1.82 ;
 RECT 7 1.82 8.58 1.96 ;
 RECT 8.44 1.79 8.58 1.82 ;
 RECT 9.015 1.58 9.255 1.65 ;
 RECT 9.015 1.79 9.255 1.835 ;
 RECT 8.44 1.65 9.255 1.79 ;
 RECT 11.075 1.415 11.215 1.455 ;
 RECT 10.165 1.455 11.215 1.595 ;
 RECT 10.165 1.41 10.465 1.455 ;
 RECT 10.325 0.81 10.465 1.41 ;
 RECT 10.165 1.595 10.465 1.62 ;
 RECT 10.325 1.62 10.465 2.18 ;
 RECT 11.075 1.275 11.595 1.415 ;
 RECT 3.01 0.925 3.15 1.245 ;
 RECT 3.01 1.385 3.15 2.11 ;
 RECT 2.285 0.785 3.15 0.925 ;
 RECT 2.5 2.11 3.15 2.25 ;
 RECT 3.01 1.245 3.58 1.385 ;
 RECT 3.44 1.19 3.58 1.245 ;
 RECT 3.44 1.385 3.58 1.42 ;
 RECT 5.515 1.63 5.655 1.99 ;
 RECT 5.515 1.475 5.86 1.63 ;
 RECT 5.6 0.825 5.74 1.475 ;
 RECT 5.405 1.99 5.655 2.13 ;
 RECT 26.88 0.29 27.25 0.43 ;
 RECT 27.11 0.43 27.25 0.71 ;
 RECT 26.88 0.22 27.11 0.29 ;
 RECT 28.53 0.85 28.67 1.385 ;
 RECT 28.215 1.525 28.355 1.73 ;
 RECT 27.11 0.71 28.67 0.85 ;
 RECT 28.215 0.51 28.355 0.71 ;
 RECT 28.215 1.385 28.67 1.525 ;
 RECT 26.14 1.145 26.28 1.345 ;
 RECT 25.82 1.485 25.96 1.76 ;
 RECT 26.14 0.73 26.28 0.935 ;
 RECT 25.82 0.355 25.96 0.59 ;
 RECT 25.82 1.345 26.28 1.485 ;
 RECT 26.095 0.935 26.325 1.145 ;
 RECT 25.82 0.59 26.28 0.73 ;
 RECT 24.12 1.225 24.35 1.245 ;
 RECT 24.12 1.195 24.71 1.225 ;
 RECT 24.26 1.015 24.57 1.035 ;
 RECT 24.12 1.035 24.57 1.055 ;
 RECT 24.395 0.64 24.535 1.015 ;
 RECT 24.57 1.225 24.71 1.75 ;
 RECT 24.275 0.5 24.535 0.64 ;
 RECT 25.17 1.035 25.4 1.055 ;
 RECT 25.17 1.195 25.4 1.245 ;
 RECT 24.12 1.055 25.4 1.195 ;
 RECT 23.28 0.36 23.51 0.43 ;
 RECT 24.675 0.36 24.815 0.565 ;
 RECT 23.28 0.22 24.815 0.36 ;
 RECT 25.415 0.705 25.555 0.75 ;
 RECT 25.54 0.995 25.845 1.205 ;
 RECT 25.54 0.89 25.68 0.995 ;
 RECT 25.415 0.75 25.68 0.89 ;
 RECT 24.675 0.565 25.555 0.705 ;
 RECT 17.78 0.63 18.01 0.635 ;
 RECT 17.78 0.775 18.01 0.84 ;
 RECT 20.365 0.37 20.505 0.635 ;
 RECT 17.775 0.635 20.505 0.775 ;
 RECT 21.24 0.37 21.38 1.46 ;
 RECT 20.365 0.23 21.38 0.37 ;
 RECT 15.055 0.36 15.285 0.68 ;
 RECT 14.12 0.68 15.285 0.685 ;
 RECT 14.12 0.895 15.285 0.91 ;
 RECT 14.115 0.685 15.285 0.895 ;
 RECT 15.055 0.22 16.435 0.36 ;
 RECT 16.295 0.36 16.435 0.675 ;
 RECT 16.295 0.675 17.62 0.815 ;
 RECT 17.36 0.23 17.62 0.43 ;
 RECT 17.36 0.22 17.59 0.23 ;
 RECT 17.48 0.43 17.62 0.675 ;
 RECT 17.48 0.815 17.62 1.98 ;
 RECT 6.995 0.52 7.64 0.66 ;
 RECT 7.5 0.66 7.64 1.015 ;
 RECT 9 0.505 9.385 0.71 ;
 RECT 7.5 1.015 9.14 1.155 ;
 RECT 9 0.71 9.14 1.015 ;
 RECT 9.155 0.5 9.385 0.505 ;
 RECT 6.31 0.5 6.565 0.965 ;
 RECT 6.31 1.67 6.45 1.82 ;
 RECT 6.31 0.965 6.45 1.44 ;
 RECT 6.31 1.44 6.565 1.67 ;
 RECT 6.18 1.82 6.45 1.96 ;
 RECT 4.305 1.01 4.445 1.195 ;
 RECT 4.305 1.335 4.445 2.11 ;
 RECT 4.305 2.25 4.445 2.255 ;
 RECT 4.305 0.87 4.73 1.01 ;
 RECT 4.305 2.11 4.73 2.25 ;
 RECT 5.275 0.67 5.415 1.195 ;
 RECT 4.305 1.195 5.415 1.335 ;
 RECT 6.705 0.36 6.845 2.035 ;
 RECT 5.275 0.53 6.16 0.67 ;
 RECT 6.02 0.22 6.845 0.36 ;
 RECT 6.66 2.17 6.8 2.305 ;
 RECT 6.66 2.035 6.845 2.17 ;
 RECT 6.02 0.36 6.16 0.53 ;
 RECT 3.79 0.5 3.93 2.25 ;
 RECT 3.79 0.36 4.855 0.5 ;
 RECT 4.49 0.22 4.855 0.36 ;
 RECT 4.49 0.5 4.855 0.615 ;
 RECT 0.94 0.72 1.08 1.195 ;
 RECT 0.94 1.335 1.08 2.27 ;
 RECT 1.725 0.525 1.865 1.195 ;
 RECT 0.94 1.195 1.865 1.335 ;
 RECT 1.725 0.385 3.15 0.525 ;
 RECT 13.68 2.42 13.91 2.54 ;
 RECT 23.28 2.42 23.42 2.52 ;
 RECT 13.68 2.28 23.42 2.42 ;
 RECT 28.055 2.48 28.195 2.52 ;
 RECT 28.055 2.27 28.285 2.48 ;
 RECT 23.28 2.52 28.195 2.66 ;
 RECT 26.9 1.18 27.04 1.605 ;
 RECT 26.76 0.73 26.9 1.04 ;
 RECT 26.695 0.59 26.97 0.73 ;
 RECT 28.02 0.99 28.25 1.04 ;
 RECT 28.02 1.18 28.25 1.2 ;
 RECT 26.76 1.04 28.25 1.18 ;
 RECT 14.78 1.51 14.92 1.695 ;
 RECT 14.71 1.695 14.99 1.835 ;
 RECT 15.72 0.905 15.86 1.37 ;
 RECT 15.72 1.51 15.86 1.7 ;
 RECT 17.105 1.25 17.335 1.37 ;
 RECT 14.78 1.37 17.335 1.51 ;
 RECT 15.655 1.7 15.93 1.84 ;
 RECT 13.155 0.525 13.295 0.855 ;
 RECT 13.155 0.995 13.295 2.065 ;
 RECT 13.445 0.82 13.675 0.855 ;
 RECT 13.445 0.995 13.675 1.03 ;
 RECT 13.155 0.855 13.675 0.995 ;
 RECT 13.815 1.565 13.955 1.985 ;
 RECT 13.815 1.985 17.085 2.125 ;
 RECT 16.855 1.66 17.085 1.985 ;
 RECT 13.77 1.355 14 1.565 ;
 RECT 8.12 1.44 8.26 1.52 ;
 RECT 7.39 1.52 8.26 1.66 ;
 RECT 9.395 0.865 9.535 1.3 ;
 RECT 8.12 1.3 9.535 1.44 ;
 RECT 9.395 1.44 9.535 2.215 ;
 END
END RSDFFSRARX2

MACRO RSDFFSRASRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 31.04 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 24.225 0.59 24.595 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 29.455 1.435 29.795 1.8 ;
 RECT 27.775 1.99 29.64 2.13 ;
 RECT 25.545 2.22 27.915 2.36 ;
 RECT 27.775 1.435 27.915 1.99 ;
 RECT 29.5 1.8 29.64 1.99 ;
 RECT 25.545 1.39 25.685 2.22 ;
 RECT 26.93 1.37 27.07 2.22 ;
 RECT 27.775 2.13 27.915 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 31.04 0.08 ;
 RECT 27.895 0.08 28.135 0.26 ;
 RECT 5.155 0.08 5.435 0.295 ;
 RECT 9.085 0.31 9.375 0.45 ;
 RECT 12.77 0.59 13.045 0.73 ;
 RECT 21.055 0.335 21.32 0.495 ;
 RECT 16.695 0.275 17.72 0.415 ;
 RECT 17.58 0.75 18.525 0.89 ;
 RECT 25.545 0.08 25.685 0.36 ;
 RECT 26.76 0.08 26.9 0.35 ;
 RECT 0.31 0.08 0.45 0.775 ;
 RECT 1.28 0.08 1.42 0.93 ;
 RECT 4.635 0.08 4.775 0.97 ;
 RECT 3.19 0.08 3.33 0.74 ;
 RECT 7.98 0.08 8.215 0.46 ;
 RECT 22.7 0.08 22.84 0.82 ;
 RECT 9.165 0.08 9.305 0.31 ;
 RECT 12.835 0.08 12.975 0.59 ;
 RECT 21.11 0.08 21.25 0.335 ;
 RECT 16.695 0.415 16.835 0.945 ;
 RECT 16.695 0.08 16.835 0.275 ;
 RECT 18.385 0.89 18.525 1.11 ;
 RECT 17.58 0.415 17.72 0.75 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.51 1.205 20.865 1.445 ;
 RECT 20.62 0.915 20.76 1.205 ;
 RECT 21.625 1.84 21.765 1.885 ;
 RECT 21.625 0.915 21.765 1.7 ;
 RECT 20.62 1.84 20.76 1.885 ;
 RECT 20.62 1.7 21.765 1.84 ;
 RECT 20.62 1.445 20.76 1.7 ;
 END
 ANTENNADIFFAREA 0.58 ;
 END QN

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.685 1.475 5.015 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.02 1.095 22.28 1.335 ;
 RECT 22.14 0.51 22.28 1.095 ;
 RECT 23.2 1.905 23.34 1.91 ;
 RECT 22.14 1.765 23.34 1.905 ;
 RECT 23.2 0.56 23.34 1.765 ;
 RECT 22.14 1.905 22.28 1.915 ;
 RECT 22.14 1.335 22.28 1.765 ;
 END
 ANTENNADIFFAREA 0.533 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.225 1.16 12.62 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.375 0.505 7.78 0.605 ;
 RECT 7.375 0.675 11.67 0.745 ;
 RECT 11.53 0.535 12.435 0.605 ;
 RECT 7.375 0.605 12.435 0.675 ;
 RECT 13.21 1.01 13.35 1.015 ;
 RECT 12.295 0.87 13.35 1.01 ;
 RECT 13.21 0.245 15.355 0.255 ;
 RECT 13.21 0.255 15.36 0.385 ;
 RECT 15.22 1.09 17.21 1.23 ;
 RECT 17.415 1.56 17.645 1.6 ;
 RECT 17.07 1.42 17.645 1.56 ;
 RECT 17.415 1.39 17.645 1.42 ;
 RECT 12.295 0.675 12.435 0.87 ;
 RECT 13.21 0.385 13.35 0.87 ;
 RECT 15.22 0.385 15.36 1.09 ;
 RECT 17.07 1.23 17.21 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.985 1.745 10.425 2.07 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.1 1.435 1.625 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.79 1.59 2.735 1.75 ;
 RECT 1.885 1.09 2.025 1.44 ;
 RECT 1.79 1.44 2.035 1.59 ;
 RECT 2.585 1.75 2.725 1.805 ;
 RECT 2.585 1.53 2.725 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.25 1.115 2.67 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 31.04 2.96 ;
 RECT 20.965 2.6 21.23 2.8 ;
 RECT 22.555 2.6 22.82 2.8 ;
 RECT 12.58 2.215 12.855 2.355 ;
 RECT 1.28 1.965 1.42 2.8 ;
 RECT 0.31 1.74 0.45 2.8 ;
 RECT 5.31 2.34 5.56 2.8 ;
 RECT 3.19 1.99 3.33 2.8 ;
 RECT 4.635 1.98 4.775 2.8 ;
 RECT 9.165 2.17 9.305 2.8 ;
 RECT 10.195 2.21 10.335 2.8 ;
 RECT 15.605 2.335 15.875 2.8 ;
 RECT 12.645 2.355 12.785 2.8 ;
 RECT 12.645 2.195 12.785 2.215 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 25.805 1.245 25.905 2.02 ;
 RECT 25.675 1.035 25.905 1.245 ;
 RECT 15.915 0.105 18.74 0.205 ;
 RECT 15.915 0.205 16.015 1.91 ;
 RECT 18.64 0.205 18.74 1.265 ;
 RECT 15.095 1.71 15.195 1.91 ;
 RECT 14.01 1.61 15.195 1.71 ;
 RECT 14.01 0.475 14.11 1.61 ;
 RECT 14.56 1.71 14.66 2.425 ;
 RECT 10.675 0.475 10.775 0.895 ;
 RECT 15.095 1.91 16.015 2.01 ;
 RECT 10.675 0.375 14.11 0.475 ;
 RECT 10.55 0.895 10.78 1.105 ;
 RECT 16.225 0.455 18.155 0.535 ;
 RECT 17.925 0.535 18.155 0.6 ;
 RECT 17.925 0.39 18.155 0.435 ;
 RECT 16.305 0.435 18.155 0.455 ;
 RECT 16.225 0.535 16.455 0.665 ;
 RECT 17.08 0.535 17.31 0.835 ;
 RECT 17.08 0.835 17.18 2.39 ;
 RECT 26.11 0.215 26.21 0.995 ;
 RECT 26.11 0.995 26.35 1.205 ;
 RECT 26.11 1.205 26.21 2 ;
 RECT 28.505 0.375 28.605 0.99 ;
 RECT 28.505 0.99 28.755 1.2 ;
 RECT 28.505 1.2 28.605 2.27 ;
 RECT 28.505 2.27 28.79 2.48 ;
 RECT 13.49 0.655 13.59 2.305 ;
 RECT 13.795 2.3 14.025 2.305 ;
 RECT 13.795 2.405 14.025 2.51 ;
 RECT 13.49 2.305 14.025 2.405 ;
 RECT 25.33 0.21 25.43 0.755 ;
 RECT 25.33 0.855 25.43 2.2 ;
 RECT 28.195 1.125 28.295 2.2 ;
 RECT 24.365 0.755 25.9 0.84 ;
 RECT 24.365 0.84 25.895 0.855 ;
 RECT 25.8 0.215 25.9 0.755 ;
 RECT 24.365 0.595 24.595 0.755 ;
 RECT 25.33 2.2 28.295 2.3 ;
 RECT 12.2 1.28 12.455 1.45 ;
 RECT 12.2 1.45 12.3 1.655 ;
 RECT 12.2 0.655 12.3 1.18 ;
 RECT 12.2 1.655 13.16 1.755 ;
 RECT 13.06 1.755 13.16 2.355 ;
 RECT 11.285 0.66 11.385 1.18 ;
 RECT 12.2 1.755 12.3 2.51 ;
 RECT 11.285 1.24 12.455 1.28 ;
 RECT 11.285 1.18 12.3 1.24 ;
 RECT 27.02 0.38 27.12 0.96 ;
 RECT 27.02 1.06 27.12 1.14 ;
 RECT 26.6 0.935 26.83 0.96 ;
 RECT 26.6 0.96 27.12 1.06 ;
 RECT 26.6 1.06 26.83 1.145 ;
 RECT 27.02 1.14 27.29 1.24 ;
 RECT 27.19 1.24 27.29 1.84 ;
 RECT 27.385 0.22 27.615 0.28 ;
 RECT 27.385 0.38 27.615 0.43 ;
 RECT 27.02 0.28 27.615 0.38 ;
 RECT 11.275 1.575 11.375 2.485 ;
 RECT 11.785 1.575 12.015 1.685 ;
 RECT 11.275 1.475 12.015 1.575 ;
 RECT 29.205 0.195 29.305 2.665 ;
 RECT 28.195 0.095 29.305 0.195 ;
 RECT 24.57 1.245 24.67 2.665 ;
 RECT 28.195 0.195 28.295 0.945 ;
 RECT 24.57 1.2 24.855 1.245 ;
 RECT 24.625 1.035 24.855 1.1 ;
 RECT 24.57 2.665 29.305 2.765 ;
 RECT 24.57 1.1 24.9 1.2 ;
 RECT 15.5 0.795 15.665 0.925 ;
 RECT 14.82 0.885 15.05 0.925 ;
 RECT 14.82 1.025 15.05 1.095 ;
 RECT 14.82 0.925 15.665 1.025 ;
 RECT 15.5 0.585 15.73 0.795 ;
 RECT 2.535 1.55 2.775 1.78 ;
 RECT 2.675 1.78 2.775 2.695 ;
 RECT 1.065 1.435 1.635 1.71 ;
 RECT 1.065 0.515 1.165 1.435 ;
 RECT 1.065 1.71 1.165 2.645 ;
 RECT 1.535 0.515 1.635 1.435 ;
 RECT 1.535 1.71 1.635 2.695 ;
 RECT 2.255 1.37 2.355 1.605 ;
 RECT 2.485 0.515 2.585 1.14 ;
 RECT 2.205 1.705 2.305 2.695 ;
 RECT 2.205 1.605 2.355 1.705 ;
 RECT 2.255 1.14 2.585 1.37 ;
 RECT 1.87 0.515 1.97 1.105 ;
 RECT 1.83 1.105 2.075 1.345 ;
 RECT 4.895 0.49 4.995 1.495 ;
 RECT 4.7 1.495 4.995 1.745 ;
 RECT 4.895 1.745 4.995 2.37 ;
 RECT 4.42 0.52 4.52 2.465 ;
 RECT 4.18 0.27 4.52 0.52 ;
 RECT 6.555 1.66 6.655 2.475 ;
 RECT 6.015 1.445 6.26 1.56 ;
 RECT 6.015 1.66 6.26 1.69 ;
 RECT 6.015 1.56 6.655 1.66 ;
 RECT 5.67 1.62 5.77 2.655 ;
 RECT 6.6 0.285 6.7 0.47 ;
 RECT 6.6 0.47 6.885 0.705 ;
 RECT 6.6 0.705 6.7 1.255 ;
 RECT 5.735 0.185 6.7 0.285 ;
 RECT 5.735 0.285 5.835 1.52 ;
 RECT 5.235 1.44 5.48 1.52 ;
 RECT 5.235 1.62 5.48 1.69 ;
 RECT 5.235 1.52 5.835 1.62 ;
 RECT 5.67 2.655 9.04 2.755 ;
 RECT 8.94 1.79 9.04 2.655 ;
 RECT 13.095 0.655 13.195 1.24 ;
 RECT 12.965 1.24 13.195 1.475 ;
 RECT 7.49 0.745 7.59 1.61 ;
 RECT 7.525 1.71 7.625 2.475 ;
 RECT 7.49 1.61 7.625 1.71 ;
 RECT 7.38 0.535 7.61 0.745 ;
 RECT 7.05 1.435 7.15 2.475 ;
 RECT 7.09 0.65 7.19 1.225 ;
 RECT 7.01 1.225 7.24 1.435 ;
 RECT 2.975 0.135 3.075 0.22 ;
 RECT 2.815 0.22 3.075 0.43 ;
 RECT 2.975 0.43 3.075 2.695 ;
 RECT 3.445 0.295 3.545 1.115 ;
 RECT 3.28 1.115 3.545 1.325 ;
 RECT 3.445 1.325 3.545 2.74 ;
 RECT 19.52 0.77 19.62 2.155 ;
 RECT 19.52 0.55 19.62 0.56 ;
 RECT 19.52 0.56 19.775 0.77 ;
 RECT 20.155 0.43 20.255 1.245 ;
 RECT 20.885 0.39 20.985 1.4 ;
 RECT 20.885 1.5 20.985 2.42 ;
 RECT 21.375 0.51 21.475 1.4 ;
 RECT 21.375 1.5 21.475 2.44 ;
 RECT 20.09 0.22 20.32 0.29 ;
 RECT 20.09 0.39 20.32 0.43 ;
 RECT 20.09 0.29 20.985 0.39 ;
 RECT 20.885 1.4 21.475 1.5 ;
 RECT 20.105 1.245 20.335 1.455 ;
 RECT 18.58 1.445 18.68 2.035 ;
 RECT 18.565 2.035 18.795 2.245 ;
 RECT 19.05 0.55 19.15 2.69 ;
 RECT 9.98 1.58 10.08 1.77 ;
 RECT 9.72 1.01 9.82 1.48 ;
 RECT 9.98 1.98 10.08 2.69 ;
 RECT 9.98 1.77 10.215 1.98 ;
 RECT 9.72 1.48 10.08 1.58 ;
 RECT 9.98 2.69 19.15 2.79 ;
 RECT 9.42 0.98 9.52 1.545 ;
 RECT 9.28 1.545 9.52 1.755 ;
 RECT 9.42 1.755 9.52 2.66 ;
 RECT 22.4 1.33 23.08 1.43 ;
 RECT 22.4 1.43 22.65 1.46 ;
 RECT 22.4 1.25 22.65 1.33 ;
 RECT 22.98 0.375 23.08 1.33 ;
 RECT 22.4 0.385 22.5 1.25 ;
 RECT 22.4 1.46 22.5 2.69 ;
 RECT 22.98 1.43 23.08 2.695 ;
 RECT 23.585 0.22 23.815 0.275 ;
 RECT 23.585 0.375 23.815 0.43 ;
 RECT 22.98 0.275 23.815 0.375 ;
 RECT 17.55 0.73 17.65 1.39 ;
 RECT 17.415 1.39 17.65 1.6 ;
 RECT 17.55 1.6 17.65 2.39 ;
 RECT 7.79 0.195 7.89 1.17 ;
 RECT 14.525 0.195 14.625 1.29 ;
 RECT 15.42 1.39 15.615 1.405 ;
 RECT 8.03 1.27 8.13 2.255 ;
 RECT 7.79 0.095 14.625 0.195 ;
 RECT 14.525 1.29 15.615 1.39 ;
 RECT 8.03 2.255 8.26 2.465 ;
 RECT 7.79 1.17 8.13 1.27 ;
 RECT 15.42 1.405 15.65 1.615 ;
 LAYER CO ;
 RECT 8.08 2.295 8.21 2.425 ;
 RECT 7.06 1.265 7.19 1.395 ;
 RECT 2.865 0.26 2.995 0.39 ;
 RECT 3.33 1.155 3.46 1.285 ;
 RECT 22.47 1.29 22.6 1.42 ;
 RECT 20.155 1.285 20.285 1.415 ;
 RECT 17.975 0.43 18.105 0.56 ;
 RECT 19.595 0.6 19.725 0.73 ;
 RECT 20.14 0.26 20.27 0.39 ;
 RECT 18.615 2.075 18.745 2.205 ;
 RECT 10.035 1.81 10.165 1.94 ;
 RECT 9.33 1.585 9.46 1.715 ;
 RECT 23.635 0.26 23.765 0.39 ;
 RECT 28.575 1.03 28.705 1.16 ;
 RECT 16.275 0.495 16.405 0.625 ;
 RECT 17.465 1.43 17.595 1.56 ;
 RECT 15.55 0.625 15.68 0.755 ;
 RECT 15.47 1.445 15.6 1.575 ;
 RECT 25.725 1.075 25.855 1.205 ;
 RECT 10.6 0.935 10.73 1.065 ;
 RECT 26.65 0.975 26.78 1.105 ;
 RECT 17.13 0.665 17.26 0.795 ;
 RECT 26.17 1.035 26.3 1.165 ;
 RECT 28.61 2.31 28.74 2.44 ;
 RECT 13.845 2.34 13.975 2.47 ;
 RECT 24.415 0.635 24.545 0.765 ;
 RECT 12.275 1.28 12.405 1.41 ;
 RECT 27.435 0.26 27.565 0.39 ;
 RECT 11.835 1.515 11.965 1.645 ;
 RECT 24.675 1.075 24.805 1.205 ;
 RECT 14.87 0.925 15 1.055 ;
 RECT 4.76 1.55 4.89 1.68 ;
 RECT 1.285 0.735 1.415 0.865 ;
 RECT 1.29 1.51 1.42 1.64 ;
 RECT 0.815 0.735 0.945 0.865 ;
 RECT 3.195 2.31 3.325 2.44 ;
 RECT 1.285 2.015 1.415 2.145 ;
 RECT 1.89 1.155 2.02 1.285 ;
 RECT 3.195 2.05 3.325 2.18 ;
 RECT 2.59 1.6 2.72 1.73 ;
 RECT 3.665 2.01 3.795 2.14 ;
 RECT 3.665 0.735 3.795 0.865 ;
 RECT 2.425 2.075 2.555 2.205 ;
 RECT 1.285 2.275 1.415 2.405 ;
 RECT 3.195 0.545 3.325 0.675 ;
 RECT 3.665 1.75 3.795 1.88 ;
 RECT 0.815 2.015 0.945 2.145 ;
 RECT 2.23 0.735 2.36 0.865 ;
 RECT 2.41 1.19 2.54 1.32 ;
 RECT 26.765 0.12 26.895 0.25 ;
 RECT 26.33 1.485 26.46 1.615 ;
 RECT 28.725 1.465 28.855 1.595 ;
 RECT 19.27 1.705 19.4 1.835 ;
 RECT 28.725 0.595 28.855 0.725 ;
 RECT 12.65 2.225 12.78 2.355 ;
 RECT 21.63 0.975 21.76 1.105 ;
 RECT 22.62 2.64 22.75 2.77 ;
 RECT 4.17 2.115 4.3 2.245 ;
 RECT 21.115 0.36 21.245 0.49 ;
 RECT 23.205 0.63 23.335 0.76 ;
 RECT 27.27 0.595 27.4 0.725 ;
 RECT 6.705 0.525 6.835 0.655 ;
 RECT 7.745 1.67 7.875 1.8 ;
 RECT 27.78 1.49 27.91 1.62 ;
 RECT 6.35 0.88 6.48 1.01 ;
 RECT 14.78 1.87 14.91 2 ;
 RECT 8.685 2.195 8.815 2.325 ;
 RECT 8.035 0.32 8.165 0.45 ;
 RECT 25.55 0.135 25.68 0.265 ;
 RECT 5.295 1.495 5.425 1.625 ;
 RECT 5.245 0.745 5.375 0.875 ;
 RECT 5.115 1.995 5.245 2.125 ;
 RECT 11.95 1.995 12.08 2.125 ;
 RECT 0.315 0.59 0.445 0.72 ;
 RECT 11.505 2.07 11.635 2.2 ;
 RECT 14.275 0.595 14.405 0.725 ;
 RECT 6.07 1.49 6.2 1.62 ;
 RECT 13.015 1.28 13.145 1.41 ;
 RECT 22.145 1.725 22.275 1.855 ;
 RECT 0.315 2.085 0.445 2.215 ;
 RECT 9.71 2.215 9.84 2.345 ;
 RECT 18.39 0.91 18.52 1.04 ;
 RECT 10.2 2.28 10.33 2.41 ;
 RECT 22.705 0.62 22.835 0.75 ;
 RECT 6.305 2.105 6.435 2.235 ;
 RECT 7.27 2.025 7.4 2.155 ;
 RECT 5.225 0.145 5.355 0.275 ;
 RECT 14.275 1.9 14.405 2.03 ;
 RECT 0.315 2.345 0.445 2.475 ;
 RECT 5.38 2.345 5.51 2.475 ;
 RECT 26.33 0.435 26.46 0.565 ;
 RECT 20.625 1.705 20.755 1.835 ;
 RECT 9.98 1.23 10.11 1.36 ;
 RECT 18.8 1.705 18.93 1.835 ;
 RECT 9.17 2.245 9.3 2.375 ;
 RECT 6.82 0.88 6.95 1.01 ;
 RECT 16.83 1.835 16.96 1.965 ;
 RECT 16.7 0.765 16.83 0.895 ;
 RECT 4.64 0.74 4.77 0.87 ;
 RECT 27.945 0.12 28.075 0.25 ;
 RECT 22.145 0.62 22.275 0.75 ;
 RECT 15.675 2.38 15.805 2.51 ;
 RECT 11.95 0.885 12.08 1.015 ;
 RECT 25.08 1.425 25.21 1.555 ;
 RECT 0.315 0.33 0.445 0.46 ;
 RECT 19.865 0.92 19.995 1.05 ;
 RECT 25.55 1.475 25.68 1.605 ;
 RECT 13.75 0.875 13.88 1.005 ;
 RECT 5.955 0.79 6.085 0.92 ;
 RECT 17.77 1.835 17.9 1.965 ;
 RECT 6.8 2.07 6.93 2.2 ;
 RECT 29.505 1.475 29.635 1.605 ;
 RECT 21.63 1.705 21.76 1.835 ;
 RECT 23.205 1.71 23.335 1.84 ;
 RECT 20.625 0.975 20.755 1.105 ;
 RECT 4.17 0.74 4.3 0.87 ;
 RECT 5.89 1.825 6.02 1.955 ;
 RECT 13.75 1.945 13.88 2.075 ;
 RECT 4.64 2.05 4.77 2.18 ;
 RECT 24.83 0.505 24.96 0.635 ;
 RECT 11.025 2.015 11.155 2.145 ;
 RECT 19.745 1.705 19.875 1.835 ;
 RECT 21.03 2.64 21.16 2.77 ;
 RECT 27.41 1.405 27.54 1.535 ;
 RECT 11.03 0.905 11.16 1.035 ;
 RECT 4.24 0.325 4.37 0.455 ;
 RECT 9.17 0.315 9.3 0.445 ;
 RECT 11.505 0.905 11.635 1.035 ;
 RECT 14.78 0.595 14.91 0.725 ;
 RECT 12.84 0.595 12.97 0.725 ;
 RECT 26.935 1.445 27.065 1.575 ;
 RECT 0.315 1.825 0.445 1.955 ;
 RECT 17.805 1.035 17.935 1.165 ;
 RECT 7.43 0.575 7.56 0.705 ;
 LAYER M1 ;
 RECT 5.195 0.88 5.335 1.475 ;
 RECT 5.045 1.99 5.295 2.13 ;
 RECT 5.195 0.74 5.515 0.88 ;
 RECT 6.64 0.875 6.955 1.08 ;
 RECT 6.64 1.08 6.78 1.665 ;
 RECT 6.64 1.805 6.78 2.015 ;
 RECT 6.64 1.685 7.95 1.805 ;
 RECT 6.765 0.8 6.955 0.875 ;
 RECT 6.64 2.015 7.005 2.215 ;
 RECT 9.28 1.685 9.51 1.755 ;
 RECT 6.64 1.665 9.51 1.685 ;
 RECT 7.68 1.545 9.51 1.665 ;
 RECT 2.88 0.87 3.02 1.15 ;
 RECT 2.88 1.29 3.02 2.07 ;
 RECT 2.175 0.73 3.02 0.87 ;
 RECT 2.37 2.07 3.02 2.21 ;
 RECT 2.88 1.15 3.51 1.29 ;
 RECT 3.28 1.115 3.51 1.15 ;
 RECT 3.28 1.29 3.51 1.325 ;
 RECT 26.645 1.145 26.785 1.345 ;
 RECT 26.325 1.485 26.465 1.76 ;
 RECT 26.645 0.73 26.785 0.935 ;
 RECT 26.325 0.355 26.465 0.59 ;
 RECT 26.325 1.345 26.785 1.485 ;
 RECT 26.6 0.935 26.83 1.145 ;
 RECT 26.325 0.59 26.785 0.73 ;
 RECT 27.265 0.73 27.405 1.04 ;
 RECT 27.405 1.18 27.545 1.605 ;
 RECT 27.2 0.59 27.475 0.73 ;
 RECT 28.525 0.99 28.755 1.04 ;
 RECT 27.265 1.04 28.755 1.18 ;
 RECT 28.525 1.18 28.755 1.2 ;
 RECT 27.385 0.29 27.755 0.43 ;
 RECT 27.615 0.43 27.755 0.71 ;
 RECT 27.385 0.22 27.615 0.29 ;
 RECT 29.035 0.85 29.175 1.385 ;
 RECT 28.72 1.525 28.86 1.73 ;
 RECT 27.615 0.71 29.175 0.85 ;
 RECT 28.72 0.51 28.86 0.71 ;
 RECT 28.72 1.385 29.175 1.525 ;
 RECT 24.625 1.225 24.855 1.245 ;
 RECT 24.625 1.195 25.215 1.225 ;
 RECT 24.765 1.015 25.075 1.035 ;
 RECT 24.625 1.035 25.075 1.055 ;
 RECT 24.9 0.64 25.04 1.015 ;
 RECT 25.075 1.225 25.215 1.75 ;
 RECT 24.78 0.5 25.04 0.64 ;
 RECT 25.675 1.035 25.905 1.055 ;
 RECT 25.675 1.195 25.905 1.245 ;
 RECT 24.625 1.055 25.905 1.195 ;
 RECT 23.585 0.36 23.815 0.43 ;
 RECT 25.18 0.36 25.32 0.565 ;
 RECT 23.585 0.22 25.32 0.36 ;
 RECT 25.92 0.705 26.06 0.75 ;
 RECT 26.045 0.995 26.35 1.205 ;
 RECT 26.045 0.89 26.185 0.995 ;
 RECT 25.92 0.75 26.185 0.89 ;
 RECT 25.18 0.565 26.06 0.705 ;
 RECT 18.82 0.775 18.96 1.405 ;
 RECT 19.545 0.56 19.775 0.635 ;
 RECT 17.8 1.405 18.96 1.545 ;
 RECT 17.8 1.545 17.94 1.83 ;
 RECT 16.755 1.83 18.005 1.97 ;
 RECT 17.8 1.17 17.94 1.405 ;
 RECT 17.73 1.03 18.01 1.17 ;
 RECT 21.74 0.36 21.88 0.635 ;
 RECT 18.82 0.635 21.88 0.775 ;
 RECT 22.42 0.36 22.56 1.25 ;
 RECT 22.42 1.25 22.65 1.46 ;
 RECT 21.74 0.22 22.56 0.36 ;
 RECT 17.925 0.28 20.32 0.42 ;
 RECT 17.925 0.42 18.155 0.6 ;
 RECT 20.09 0.22 20.32 0.28 ;
 RECT 20.09 0.42 20.32 0.43 ;
 RECT 17.08 0.57 17.31 0.95 ;
 RECT 14.775 0.525 14.915 0.885 ;
 RECT 14.775 1.095 14.915 2.065 ;
 RECT 14.775 0.885 15.05 1.095 ;
 RECT 11.5 1.04 11.64 2.34 ;
 RECT 11.5 0.895 11.64 0.9 ;
 RECT 11.43 0.9 11.705 1.04 ;
 RECT 12.295 2.055 12.435 2.34 ;
 RECT 11.5 2.34 12.435 2.48 ;
 RECT 12.295 1.915 14.41 2.055 ;
 RECT 13.745 0.765 13.885 1.915 ;
 RECT 13.745 2.055 13.885 2.145 ;
 RECT 14.27 0.525 14.41 1.915 ;
 RECT 14.27 2.055 14.41 2.11 ;
 RECT 15.5 0.585 16.455 0.63 ;
 RECT 16.225 0.63 16.455 0.665 ;
 RECT 16.225 0.455 16.455 0.49 ;
 RECT 15.525 0.49 16.455 0.585 ;
 RECT 15.5 0.63 15.73 0.795 ;
 RECT 5.95 1.67 6.09 1.82 ;
 RECT 5.95 1.96 6.09 2.51 ;
 RECT 5.95 0.5 6.09 1.44 ;
 RECT 5.95 1.44 6.205 1.67 ;
 RECT 5.82 1.82 6.13 1.96 ;
 RECT 8.03 2.255 8.26 2.51 ;
 RECT 5.95 2.51 8.26 2.65 ;
 RECT 3.945 0.875 4.085 1.195 ;
 RECT 3.945 1.335 4.085 2.11 ;
 RECT 3.945 2.25 4.085 2.255 ;
 RECT 3.945 0.735 4.37 0.875 ;
 RECT 3.945 2.11 4.37 2.25 ;
 RECT 3.945 1.195 5.055 1.335 ;
 RECT 4.915 0.6 5.055 1.195 ;
 RECT 6.345 0.36 6.485 2.035 ;
 RECT 5.66 0.36 5.8 0.46 ;
 RECT 5.66 0.22 6.485 0.36 ;
 RECT 6.3 2.17 6.44 2.305 ;
 RECT 4.915 0.46 5.8 0.6 ;
 RECT 6.3 2.035 6.485 2.17 ;
 RECT 7.095 0.66 7.235 0.895 ;
 RECT 6.635 0.52 7.235 0.66 ;
 RECT 7.095 0.895 10.78 1.035 ;
 RECT 10.55 1.035 10.78 1.105 ;
 RECT 3.66 0.46 3.8 2.21 ;
 RECT 4.13 0.22 4.495 0.32 ;
 RECT 4.13 0.46 4.495 0.525 ;
 RECT 3.66 0.32 4.495 0.46 ;
 RECT 0.81 0.68 0.95 1.155 ;
 RECT 0.81 1.295 0.95 2.23 ;
 RECT 1.595 0.36 1.735 1.155 ;
 RECT 0.81 1.155 1.735 1.295 ;
 RECT 2.815 0.36 3.045 0.43 ;
 RECT 1.595 0.22 3.045 0.36 ;
 RECT 19.63 1.7 19.925 1.84 ;
 RECT 19.63 1.84 19.77 2.075 ;
 RECT 18.935 1.84 19.075 2.075 ;
 RECT 18.74 1.7 19.075 1.84 ;
 RECT 18.935 2.075 19.77 2.215 ;
 RECT 19.825 1.055 19.965 1.245 ;
 RECT 19.265 1.385 19.405 1.625 ;
 RECT 20.105 1.385 20.335 1.455 ;
 RECT 19.265 1.245 20.335 1.385 ;
 RECT 19.795 0.915 20.095 1.055 ;
 RECT 19.235 1.625 19.49 1.92 ;
 RECT 20.335 2.205 20.475 2.39 ;
 RECT 16.19 1.895 16.33 2.39 ;
 RECT 16.19 2.39 20.475 2.53 ;
 RECT 15.065 1.755 16.33 1.895 ;
 RECT 15.065 1.895 15.205 2.34 ;
 RECT 13.795 2.3 14.025 2.34 ;
 RECT 13.795 2.48 14.025 2.51 ;
 RECT 13.795 2.34 15.205 2.48 ;
 RECT 20.335 2.065 24.36 2.205 ;
 RECT 24.22 2.205 24.36 2.52 ;
 RECT 28.56 2.48 28.7 2.52 ;
 RECT 24.22 2.52 28.7 2.66 ;
 RECT 28.56 2.27 28.79 2.48 ;
 RECT 11.945 1.02 12.085 1.475 ;
 RECT 11.785 1.475 12.085 1.635 ;
 RECT 11.945 1.775 12.085 2.18 ;
 RECT 11.875 0.88 12.15 1.02 ;
 RECT 11.945 1.685 13.15 1.775 ;
 RECT 13.01 1.415 13.15 1.635 ;
 RECT 11.785 1.635 13.15 1.685 ;
 RECT 12.96 1.275 13.215 1.415 ;
 RECT 16.47 1.56 16.61 2.11 ;
 RECT 15.42 1.405 15.65 1.42 ;
 RECT 15.42 1.56 15.65 1.615 ;
 RECT 15.42 1.42 16.61 1.56 ;
 RECT 16.47 2.11 18.795 2.245 ;
 RECT 16.47 2.245 18.79 2.25 ;
 RECT 18.565 2.035 18.795 2.11 ;
 RECT 7.2 2.115 7.475 2.205 ;
 RECT 8.61 2.115 8.885 2.375 ;
 RECT 7.2 1.975 8.885 2.115 ;
 RECT 9.705 1.365 9.845 2.41 ;
 RECT 7.01 1.365 7.24 1.435 ;
 RECT 11.02 1.04 11.16 1.25 ;
 RECT 11.02 1.39 11.16 2.215 ;
 RECT 11.02 0.885 11.16 0.9 ;
 RECT 7.01 1.25 11.16 1.365 ;
 RECT 7.01 1.225 10.41 1.25 ;
 RECT 10.27 1.365 11.16 1.39 ;
 RECT 10.955 0.9 11.23 1.04 ;
 RECT 5.155 1.475 5.5 1.63 ;
 RECT 5.155 1.63 5.295 1.99 ;
 END
END RSDFFSRASRX1

MACRO RSDFFSRASRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 33.6 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 26.695 0.59 27.065 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 31.925 1.435 32.265 1.8 ;
 RECT 30.245 1.99 32.11 2.13 ;
 RECT 28.015 2.22 30.385 2.36 ;
 RECT 31.97 1.8 32.11 1.99 ;
 RECT 30.245 1.435 30.385 1.99 ;
 RECT 28.015 1.39 28.155 2.22 ;
 RECT 29.4 1.37 29.54 2.22 ;
 RECT 30.245 2.13 30.385 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 33.6 0.08 ;
 RECT 9.075 0.31 9.365 0.45 ;
 RECT 12.76 0.59 13.03 0.73 ;
 RECT 16.685 0.275 17.71 0.415 ;
 RECT 22.01 0.335 22.275 0.495 ;
 RECT 21.015 0.335 21.28 0.495 ;
 RECT 17.57 0.75 18.515 0.89 ;
 RECT 4.515 0.08 4.655 0.97 ;
 RECT 3.18 0.08 3.32 0.74 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 0.93 ;
 RECT 5.145 0.08 5.425 0.295 ;
 RECT 7.97 0.08 8.205 0.46 ;
 RECT 23.815 0.08 23.955 0.82 ;
 RECT 28.015 0.08 28.155 0.36 ;
 RECT 24.87 0.08 25.01 0.82 ;
 RECT 30.365 0.08 30.605 0.26 ;
 RECT 29.23 0.08 29.37 0.35 ;
 RECT 9.155 0.08 9.295 0.31 ;
 RECT 12.825 0.08 12.965 0.59 ;
 RECT 16.685 0.415 16.825 0.945 ;
 RECT 16.685 0.08 16.825 0.275 ;
 RECT 22.065 0.08 22.205 0.335 ;
 RECT 21.07 0.08 21.21 0.335 ;
 RECT 18.375 0.89 18.515 1.11 ;
 RECT 17.57 0.415 17.71 0.75 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.6 1.475 4.93 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.215 1.16 12.615 1.49 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.365 0.485 7.68 0.605 ;
 RECT 7.365 0.625 11.72 0.745 ;
 RECT 11.58 0.485 12.425 0.605 ;
 RECT 7.365 0.605 12.425 0.625 ;
 RECT 12.285 0.875 13.34 1.015 ;
 RECT 13.2 0.245 15.345 0.255 ;
 RECT 13.2 0.255 15.35 0.385 ;
 RECT 15.21 1.09 17.2 1.23 ;
 RECT 17.405 1.56 17.635 1.6 ;
 RECT 17.06 1.42 17.635 1.56 ;
 RECT 17.405 1.39 17.635 1.42 ;
 RECT 12.285 0.625 12.425 0.875 ;
 RECT 13.2 0.385 13.34 0.875 ;
 RECT 15.21 0.385 15.35 1.09 ;
 RECT 17.06 1.23 17.2 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.975 1.765 10.415 2.06 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.435 1.615 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.78 1.59 2.725 1.75 ;
 RECT 1.875 1.09 2.015 1.44 ;
 RECT 1.78 1.44 2.025 1.59 ;
 RECT 2.575 1.75 2.715 1.805 ;
 RECT 2.575 1.53 2.715 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.24 1.115 2.66 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 33.6 2.96 ;
 RECT 12.57 2.215 12.845 2.355 ;
 RECT 1.27 1.965 1.41 2.8 ;
 RECT 3.18 1.99 3.32 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 4.49 1.98 4.63 2.8 ;
 RECT 5.18 2.34 5.43 2.8 ;
 RECT 9.155 2.16 9.295 2.8 ;
 RECT 10.185 2.2 10.325 2.8 ;
 RECT 15.595 2.335 15.865 2.8 ;
 RECT 21.92 2.6 22.185 2.8 ;
 RECT 20.925 2.6 21.19 2.8 ;
 RECT 23.67 2.6 23.935 2.8 ;
 RECT 24.725 2.6 24.99 2.8 ;
 RECT 12.635 2.355 12.775 2.8 ;
 RECT 12.635 2.195 12.775 2.215 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.47 1.205 20.72 1.445 ;
 RECT 20.58 0.915 20.72 1.205 ;
 RECT 21.585 1.84 21.725 1.885 ;
 RECT 21.585 0.915 21.725 1.7 ;
 RECT 22.58 1.84 22.72 1.885 ;
 RECT 22.58 0.915 22.72 1.7 ;
 RECT 20.58 1.7 22.77 1.84 ;
 RECT 20.58 1.84 20.72 1.885 ;
 RECT 20.58 1.445 20.72 1.7 ;
 END
 ANTENNADIFFAREA 0.883 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 23.135 1.095 23.395 1.335 ;
 RECT 23.255 0.51 23.395 1.095 ;
 RECT 24.315 1.905 24.455 1.91 ;
 RECT 24.315 0.56 24.455 1.765 ;
 RECT 25.37 1.905 25.51 1.91 ;
 RECT 25.37 0.56 25.51 1.765 ;
 RECT 23.255 1.905 23.395 1.915 ;
 RECT 23.255 1.335 23.395 1.765 ;
 RECT 23.255 1.765 25.51 1.905 ;
 END
 ANTENNADIFFAREA 0.854 ;
 END Q

 OBS
 LAYER PO ;
 RECT 15.905 0.205 16.005 1.91 ;
 RECT 18.63 0.205 18.73 1.265 ;
 RECT 15.085 1.71 15.185 1.91 ;
 RECT 14 1.61 15.185 1.71 ;
 RECT 14 0.475 14.1 1.61 ;
 RECT 14.55 1.71 14.65 2.425 ;
 RECT 10.665 0.475 10.765 0.895 ;
 RECT 15.085 1.91 16.005 2.01 ;
 RECT 10.665 0.375 14.1 0.475 ;
 RECT 10.54 0.895 10.77 1.105 ;
 RECT 16.215 0.455 18.145 0.535 ;
 RECT 17.915 0.535 18.145 0.6 ;
 RECT 17.915 0.39 18.145 0.435 ;
 RECT 16.295 0.435 18.145 0.455 ;
 RECT 16.215 0.535 16.445 0.665 ;
 RECT 17.07 0.535 17.3 0.835 ;
 RECT 17.07 0.835 17.17 2.39 ;
 RECT 28.58 0.215 28.68 0.995 ;
 RECT 28.58 0.995 28.82 1.205 ;
 RECT 28.58 1.205 28.68 2 ;
 RECT 30.975 0.375 31.075 0.99 ;
 RECT 30.975 0.99 31.225 1.2 ;
 RECT 30.975 1.2 31.075 2.27 ;
 RECT 30.975 2.27 31.26 2.48 ;
 RECT 13.48 0.655 13.58 2.305 ;
 RECT 13.785 2.3 14.015 2.305 ;
 RECT 13.785 2.405 14.015 2.51 ;
 RECT 13.48 2.305 14.015 2.405 ;
 RECT 27.8 0.855 27.9 2.2 ;
 RECT 30.665 1.125 30.765 2.2 ;
 RECT 26.835 0.755 28.37 0.84 ;
 RECT 26.835 0.84 28.365 0.855 ;
 RECT 28.27 0.215 28.37 0.755 ;
 RECT 27.8 0.21 27.9 0.755 ;
 RECT 26.835 0.595 27.065 0.755 ;
 RECT 27.8 2.2 30.765 2.3 ;
 RECT 12.19 1.28 12.445 1.45 ;
 RECT 12.19 1.45 12.29 1.655 ;
 RECT 12.19 0.655 12.29 1.18 ;
 RECT 12.19 1.655 13.15 1.755 ;
 RECT 13.05 1.755 13.15 2.355 ;
 RECT 11.275 0.66 11.375 1.18 ;
 RECT 12.19 1.755 12.29 2.51 ;
 RECT 11.275 1.24 12.445 1.28 ;
 RECT 11.275 1.18 12.29 1.24 ;
 RECT 29.49 0.38 29.59 0.96 ;
 RECT 29.49 1.06 29.59 1.14 ;
 RECT 29.07 0.935 29.3 0.96 ;
 RECT 29.07 0.96 29.59 1.06 ;
 RECT 29.07 1.06 29.3 1.145 ;
 RECT 29.49 1.14 29.76 1.24 ;
 RECT 29.66 1.24 29.76 1.84 ;
 RECT 29.855 0.22 30.085 0.28 ;
 RECT 29.855 0.38 30.085 0.43 ;
 RECT 29.49 0.28 30.085 0.38 ;
 RECT 11.265 1.575 11.365 2.485 ;
 RECT 11.775 1.575 12.005 1.685 ;
 RECT 11.265 1.475 12.005 1.575 ;
 RECT 31.675 0.195 31.775 2.665 ;
 RECT 30.665 0.095 31.775 0.195 ;
 RECT 27.04 1.245 27.14 2.665 ;
 RECT 30.665 0.195 30.765 0.945 ;
 RECT 27.04 1.2 27.325 1.245 ;
 RECT 27.095 1.035 27.325 1.1 ;
 RECT 27.04 2.665 31.775 2.765 ;
 RECT 27.04 1.1 27.37 1.2 ;
 RECT 15.49 0.795 15.655 0.925 ;
 RECT 14.81 0.885 15.04 0.925 ;
 RECT 14.81 1.025 15.04 1.095 ;
 RECT 14.81 0.925 15.655 1.025 ;
 RECT 15.49 0.585 15.72 0.795 ;
 RECT 2.525 1.55 2.765 1.78 ;
 RECT 2.665 1.78 2.765 2.695 ;
 RECT 1.055 1.435 1.625 1.71 ;
 RECT 1.055 0.515 1.155 1.435 ;
 RECT 1.055 1.71 1.155 2.645 ;
 RECT 1.525 0.515 1.625 1.435 ;
 RECT 1.525 1.71 1.625 2.695 ;
 RECT 2.245 1.37 2.345 1.605 ;
 RECT 2.475 0.515 2.575 1.14 ;
 RECT 2.195 1.705 2.295 2.695 ;
 RECT 2.195 1.605 2.345 1.705 ;
 RECT 2.245 1.14 2.575 1.37 ;
 RECT 1.86 0.515 1.96 1.105 ;
 RECT 1.82 1.105 2.065 1.345 ;
 RECT 7.48 0.715 7.58 1.61 ;
 RECT 7.515 1.71 7.615 2.475 ;
 RECT 7.48 1.61 7.615 1.71 ;
 RECT 7.36 0.485 7.6 0.715 ;
 RECT 4.275 0.52 4.375 2.465 ;
 RECT 4.13 0.27 4.375 0.52 ;
 RECT 13.085 0.655 13.185 1.24 ;
 RECT 12.955 1.24 13.185 1.475 ;
 RECT 4.81 0.49 4.91 1.495 ;
 RECT 4.615 1.495 4.91 1.745 ;
 RECT 4.81 1.745 4.91 2.37 ;
 RECT 5.635 0.285 5.735 1.52 ;
 RECT 5.635 1.62 5.735 2.655 ;
 RECT 6.48 0.285 6.58 0.485 ;
 RECT 5.635 2.655 9.03 2.755 ;
 RECT 8.93 1.79 9.03 2.655 ;
 RECT 5.18 1.44 5.425 1.52 ;
 RECT 5.18 1.52 5.735 1.62 ;
 RECT 5.18 1.62 5.425 1.69 ;
 RECT 5.635 0.185 6.58 0.285 ;
 RECT 6.48 0.485 6.795 0.695 ;
 RECT 6.48 0.695 6.58 1.255 ;
 RECT 6.545 1.66 6.645 2.475 ;
 RECT 5.915 1.45 6.145 1.56 ;
 RECT 5.915 1.56 6.645 1.66 ;
 RECT 7.04 1.435 7.14 2.475 ;
 RECT 7.08 0.65 7.18 1.225 ;
 RECT 7 1.225 7.23 1.435 ;
 RECT 2.965 0.135 3.065 0.22 ;
 RECT 2.805 0.22 3.065 0.43 ;
 RECT 2.965 0.43 3.065 2.695 ;
 RECT 3.435 0.295 3.535 1.115 ;
 RECT 3.27 1.115 3.535 1.325 ;
 RECT 3.435 1.325 3.535 2.74 ;
 RECT 19.51 0.77 19.61 2.155 ;
 RECT 19.51 0.55 19.61 0.56 ;
 RECT 19.51 0.56 19.765 0.77 ;
 RECT 20.08 0.195 20.31 0.43 ;
 RECT 20.845 0.195 20.945 1.4 ;
 RECT 20.845 1.5 20.945 2.42 ;
 RECT 21.84 0.54 21.94 1.4 ;
 RECT 20.845 1.4 22.43 1.5 ;
 RECT 22.33 0.51 22.43 1.4 ;
 RECT 22.33 1.5 22.43 2.44 ;
 RECT 21.84 1.5 21.94 2.42 ;
 RECT 21.335 0.51 21.435 1.4 ;
 RECT 21.335 1.5 21.435 2.44 ;
 RECT 20.145 0.43 20.245 1.245 ;
 RECT 20.095 1.245 20.325 1.455 ;
 RECT 20.08 0.095 20.945 0.195 ;
 RECT 18.57 1.445 18.67 2.035 ;
 RECT 18.555 2.035 18.785 2.245 ;
 RECT 19.04 0.55 19.14 2.69 ;
 RECT 9.97 1.58 10.07 1.78 ;
 RECT 9.71 1.01 9.81 1.48 ;
 RECT 9.97 1.99 10.07 2.69 ;
 RECT 9.97 1.78 10.205 1.99 ;
 RECT 9.71 1.48 10.07 1.58 ;
 RECT 9.97 2.69 19.14 2.79 ;
 RECT 9.41 0.98 9.51 1.545 ;
 RECT 9.27 1.545 9.51 1.755 ;
 RECT 9.41 1.755 9.51 2.64 ;
 RECT 23.515 1.33 25.25 1.43 ;
 RECT 23.515 1.43 23.765 1.46 ;
 RECT 23.515 1.25 23.765 1.33 ;
 RECT 24.57 1.43 24.67 2.69 ;
 RECT 25.15 0.375 25.25 1.33 ;
 RECT 23.515 0.385 23.615 1.25 ;
 RECT 23.515 1.46 23.615 2.69 ;
 RECT 24.095 0.385 24.195 1.33 ;
 RECT 24.095 1.43 24.195 2.695 ;
 RECT 24.57 0.385 24.67 1.33 ;
 RECT 25.15 1.43 25.25 2.695 ;
 RECT 26.055 0.22 26.285 0.275 ;
 RECT 26.055 0.375 26.285 0.43 ;
 RECT 25.15 0.275 26.285 0.375 ;
 RECT 17.54 0.73 17.64 1.39 ;
 RECT 17.405 1.39 17.64 1.6 ;
 RECT 17.54 1.6 17.64 2.39 ;
 RECT 7.78 0.195 7.88 1.17 ;
 RECT 14.515 0.195 14.615 1.29 ;
 RECT 15.41 1.39 15.605 1.405 ;
 RECT 8.02 1.27 8.12 2.265 ;
 RECT 7.78 0.095 14.615 0.195 ;
 RECT 14.515 1.29 15.605 1.39 ;
 RECT 8.02 2.265 8.25 2.475 ;
 RECT 7.78 1.17 8.12 1.27 ;
 RECT 15.41 1.405 15.64 1.615 ;
 RECT 28.275 1.245 28.375 2.02 ;
 RECT 28.145 1.035 28.375 1.245 ;
 RECT 15.905 0.105 18.73 0.205 ;
 LAYER CO ;
 RECT 18.605 2.075 18.735 2.205 ;
 RECT 10.025 1.82 10.155 1.95 ;
 RECT 9.32 1.585 9.45 1.715 ;
 RECT 26.105 0.26 26.235 0.39 ;
 RECT 31.045 1.03 31.175 1.16 ;
 RECT 16.265 0.495 16.395 0.625 ;
 RECT 17.455 1.43 17.585 1.56 ;
 RECT 15.54 0.625 15.67 0.755 ;
 RECT 15.46 1.445 15.59 1.575 ;
 RECT 28.195 1.075 28.325 1.205 ;
 RECT 10.59 0.935 10.72 1.065 ;
 RECT 29.12 0.975 29.25 1.105 ;
 RECT 17.12 0.665 17.25 0.795 ;
 RECT 28.64 1.035 28.77 1.165 ;
 RECT 31.08 2.31 31.21 2.44 ;
 RECT 13.835 2.34 13.965 2.47 ;
 RECT 26.885 0.635 27.015 0.765 ;
 RECT 12.265 1.28 12.395 1.41 ;
 RECT 29.905 0.26 30.035 0.39 ;
 RECT 11.825 1.515 11.955 1.645 ;
 RECT 27.145 1.075 27.275 1.205 ;
 RECT 14.86 0.925 14.99 1.055 ;
 RECT 4.675 1.55 4.805 1.68 ;
 RECT 20.585 1.705 20.715 1.835 ;
 RECT 21.59 1.705 21.72 1.835 ;
 RECT 20.585 0.975 20.715 1.105 ;
 RECT 21.59 0.975 21.72 1.105 ;
 RECT 21.075 0.36 21.205 0.49 ;
 RECT 1.275 0.735 1.405 0.865 ;
 RECT 1.28 1.51 1.41 1.64 ;
 RECT 0.805 0.735 0.935 0.865 ;
 RECT 3.185 2.31 3.315 2.44 ;
 RECT 1.275 2.015 1.405 2.145 ;
 RECT 1.88 1.155 2.01 1.285 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 2.58 1.6 2.71 1.73 ;
 RECT 3.655 2.01 3.785 2.14 ;
 RECT 3.655 0.735 3.785 0.865 ;
 RECT 2.415 2.075 2.545 2.205 ;
 RECT 1.275 2.275 1.405 2.405 ;
 RECT 3.185 0.545 3.315 0.675 ;
 RECT 3.655 1.75 3.785 1.88 ;
 RECT 0.805 2.015 0.935 2.145 ;
 RECT 2.22 0.735 2.35 0.865 ;
 RECT 2.4 1.19 2.53 1.32 ;
 RECT 30.25 1.49 30.38 1.62 ;
 RECT 6.23 0.88 6.36 1.01 ;
 RECT 14.77 1.87 14.9 2 ;
 RECT 8.675 2.185 8.805 2.315 ;
 RECT 8.025 0.32 8.155 0.45 ;
 RECT 28.02 0.135 28.15 0.265 ;
 RECT 5.24 1.495 5.37 1.625 ;
 RECT 5.145 0.745 5.275 0.875 ;
 RECT 5.03 1.995 5.16 2.125 ;
 RECT 11.94 1.995 12.07 2.125 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 11.495 2.07 11.625 2.2 ;
 RECT 14.265 0.595 14.395 0.725 ;
 RECT 13.005 1.28 13.135 1.41 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 23.26 1.725 23.39 1.855 ;
 RECT 23.82 0.62 23.95 0.75 ;
 RECT 23.26 0.62 23.39 0.75 ;
 RECT 24.32 1.71 24.45 1.84 ;
 RECT 23.735 2.64 23.865 2.77 ;
 RECT 24.32 0.63 24.45 0.76 ;
 RECT 20.99 2.64 21.12 2.77 ;
 RECT 9.7 2.205 9.83 2.335 ;
 RECT 18.79 1.705 18.92 1.835 ;
 RECT 9.16 2.235 9.29 2.365 ;
 RECT 6.7 0.88 6.83 1.01 ;
 RECT 16.82 1.835 16.95 1.965 ;
 RECT 16.69 0.765 16.82 0.895 ;
 RECT 4.52 0.74 4.65 0.87 ;
 RECT 30.415 0.12 30.545 0.25 ;
 RECT 7.415 0.53 7.545 0.66 ;
 RECT 15.665 2.38 15.795 2.51 ;
 RECT 11.94 0.885 12.07 1.015 ;
 RECT 27.55 1.425 27.68 1.555 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 19.855 0.92 19.985 1.05 ;
 RECT 28.02 1.475 28.15 1.605 ;
 RECT 13.74 0.875 13.87 1.005 ;
 RECT 5.855 0.79 5.985 0.92 ;
 RECT 17.76 1.835 17.89 1.965 ;
 RECT 6.79 2.07 6.92 2.2 ;
 RECT 31.975 1.475 32.105 1.605 ;
 RECT 22.585 1.705 22.715 1.835 ;
 RECT 25.375 1.71 25.505 1.84 ;
 RECT 4.025 0.74 4.155 0.87 ;
 RECT 5.86 1.825 5.99 1.955 ;
 RECT 13.74 1.945 13.87 2.075 ;
 RECT 4.495 2.05 4.625 2.18 ;
 RECT 27.3 0.505 27.43 0.635 ;
 RECT 11.015 2.015 11.145 2.145 ;
 RECT 29.235 0.12 29.365 0.25 ;
 RECT 28.8 1.485 28.93 1.615 ;
 RECT 31.195 1.465 31.325 1.595 ;
 RECT 19.26 1.705 19.39 1.835 ;
 RECT 31.195 0.595 31.325 0.725 ;
 RECT 12.64 2.225 12.77 2.355 ;
 RECT 22.585 0.975 22.715 1.105 ;
 RECT 24.79 2.64 24.92 2.77 ;
 RECT 4.025 2.115 4.155 2.245 ;
 RECT 22.07 0.36 22.2 0.49 ;
 RECT 25.375 0.63 25.505 0.76 ;
 RECT 29.74 0.595 29.87 0.725 ;
 RECT 7.74 1.675 7.87 1.805 ;
 RECT 19.735 1.705 19.865 1.835 ;
 RECT 21.985 2.64 22.115 2.77 ;
 RECT 29.88 1.405 30.01 1.535 ;
 RECT 11.02 0.905 11.15 1.035 ;
 RECT 4.19 0.325 4.32 0.455 ;
 RECT 9.16 0.315 9.29 0.445 ;
 RECT 11.495 0.905 11.625 1.035 ;
 RECT 14.77 0.595 14.9 0.725 ;
 RECT 12.83 0.595 12.96 0.725 ;
 RECT 29.405 1.445 29.535 1.575 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 17.795 1.035 17.925 1.165 ;
 RECT 18.38 0.91 18.51 1.04 ;
 RECT 10.19 2.27 10.32 2.4 ;
 RECT 24.875 0.62 25.005 0.75 ;
 RECT 6.29 2.105 6.42 2.235 ;
 RECT 7.26 2.025 7.39 2.155 ;
 RECT 5.215 0.145 5.345 0.275 ;
 RECT 14.265 1.9 14.395 2.03 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 5.23 2.345 5.36 2.475 ;
 RECT 28.8 0.435 28.93 0.565 ;
 RECT 9.97 1.23 10.1 1.36 ;
 RECT 23.585 1.29 23.715 1.42 ;
 RECT 6.615 0.525 6.745 0.655 ;
 RECT 5.965 1.49 6.095 1.62 ;
 RECT 8.07 2.305 8.2 2.435 ;
 RECT 7.05 1.265 7.18 1.395 ;
 RECT 2.855 0.26 2.985 0.39 ;
 RECT 3.32 1.155 3.45 1.285 ;
 RECT 20.145 1.285 20.275 1.415 ;
 RECT 17.965 0.43 18.095 0.56 ;
 RECT 19.585 0.6 19.715 0.73 ;
 RECT 20.13 0.26 20.26 0.39 ;
 LAYER M1 ;
 RECT 5.075 0.715 5.325 0.93 ;
 RECT 5.14 1.44 5.47 1.69 ;
 RECT 4.96 1.99 5.28 2.13 ;
 RECT 2.87 0.87 3.01 1.15 ;
 RECT 2.87 1.29 3.01 2.07 ;
 RECT 2.165 0.73 3.01 0.87 ;
 RECT 2.36 2.07 3.01 2.21 ;
 RECT 2.87 1.15 3.5 1.29 ;
 RECT 3.27 1.115 3.5 1.15 ;
 RECT 3.27 1.29 3.5 1.325 ;
 RECT 29.735 0.73 29.875 1.04 ;
 RECT 29.875 1.18 30.015 1.605 ;
 RECT 29.67 0.59 29.945 0.73 ;
 RECT 30.995 0.99 31.225 1.04 ;
 RECT 29.735 1.04 31.225 1.18 ;
 RECT 30.995 1.18 31.225 1.2 ;
 RECT 29.855 0.29 30.225 0.43 ;
 RECT 30.085 0.43 30.225 0.71 ;
 RECT 29.855 0.22 30.085 0.29 ;
 RECT 31.505 0.85 31.645 1.385 ;
 RECT 31.19 1.525 31.33 1.73 ;
 RECT 30.085 0.71 31.645 0.85 ;
 RECT 31.19 0.51 31.33 0.71 ;
 RECT 31.19 1.385 31.645 1.525 ;
 RECT 27.095 1.225 27.325 1.245 ;
 RECT 27.095 1.195 27.685 1.225 ;
 RECT 27.235 1.015 27.545 1.035 ;
 RECT 27.095 1.035 27.545 1.055 ;
 RECT 27.37 0.64 27.51 1.015 ;
 RECT 27.545 1.225 27.685 1.75 ;
 RECT 27.25 0.5 27.51 0.64 ;
 RECT 28.145 1.035 28.375 1.055 ;
 RECT 28.145 1.195 28.375 1.245 ;
 RECT 27.095 1.055 28.375 1.195 ;
 RECT 29.115 1.145 29.255 1.345 ;
 RECT 28.795 1.485 28.935 1.76 ;
 RECT 29.115 0.73 29.255 0.935 ;
 RECT 28.795 0.355 28.935 0.59 ;
 RECT 28.795 1.345 29.255 1.485 ;
 RECT 29.07 0.935 29.3 1.145 ;
 RECT 28.795 0.59 29.255 0.73 ;
 RECT 26.055 0.36 26.285 0.43 ;
 RECT 27.65 0.36 27.79 0.565 ;
 RECT 26.055 0.22 27.79 0.36 ;
 RECT 28.39 0.705 28.53 0.75 ;
 RECT 28.515 0.995 28.82 1.205 ;
 RECT 28.515 0.89 28.655 0.995 ;
 RECT 28.39 0.75 28.655 0.89 ;
 RECT 27.65 0.565 28.53 0.705 ;
 RECT 14.765 0.525 14.905 0.885 ;
 RECT 14.765 1.095 14.905 2.065 ;
 RECT 14.765 0.885 15.04 1.095 ;
 RECT 18.81 0.775 18.95 1.405 ;
 RECT 19.535 0.56 19.765 0.635 ;
 RECT 17.79 1.405 18.95 1.545 ;
 RECT 17.79 1.545 17.93 1.83 ;
 RECT 16.745 1.83 17.995 1.97 ;
 RECT 17.79 1.17 17.93 1.405 ;
 RECT 17.72 1.03 18 1.17 ;
 RECT 22.835 0.36 22.975 0.635 ;
 RECT 18.81 0.635 22.975 0.775 ;
 RECT 23.535 0.36 23.675 1.25 ;
 RECT 23.535 1.25 23.765 1.46 ;
 RECT 22.835 0.22 23.675 0.36 ;
 RECT 20.08 0.22 20.31 0.28 ;
 RECT 20.08 0.42 20.31 0.43 ;
 RECT 17.915 0.28 20.31 0.42 ;
 RECT 17.915 0.42 18.145 0.6 ;
 RECT 15.49 0.585 16.445 0.63 ;
 RECT 16.215 0.63 16.445 0.665 ;
 RECT 16.215 0.455 16.445 0.49 ;
 RECT 15.515 0.49 16.445 0.585 ;
 RECT 15.49 0.63 15.72 0.795 ;
 RECT 17.07 0.57 17.3 0.95 ;
 RECT 11.49 1.04 11.63 2.34 ;
 RECT 11.49 0.895 11.63 0.9 ;
 RECT 11.42 0.9 11.695 1.04 ;
 RECT 12.285 2.055 12.425 2.34 ;
 RECT 11.49 2.34 12.425 2.48 ;
 RECT 13.42 1.66 13.56 1.915 ;
 RECT 12.285 1.915 13.56 2.055 ;
 RECT 13.735 0.765 13.875 1.52 ;
 RECT 13.735 1.66 13.875 2.145 ;
 RECT 14.26 0.525 14.4 1.52 ;
 RECT 14.26 1.66 14.4 2.11 ;
 RECT 13.42 1.52 14.4 1.66 ;
 RECT 7.085 0.66 7.225 0.895 ;
 RECT 6.565 0.485 6.795 0.52 ;
 RECT 6.565 0.66 6.795 0.695 ;
 RECT 6.565 0.52 7.225 0.66 ;
 RECT 7.085 0.895 10.77 1.035 ;
 RECT 10.54 1.035 10.77 1.105 ;
 RECT 3.935 0.875 4.075 1.195 ;
 RECT 3.935 1.335 4.075 2.11 ;
 RECT 3.935 0.735 4.225 0.875 ;
 RECT 3.935 2.11 4.225 2.25 ;
 RECT 4.795 0.575 4.935 1.195 ;
 RECT 3.935 1.195 4.935 1.335 ;
 RECT 6.285 0.36 6.425 0.875 ;
 RECT 6.285 1.015 6.425 2.305 ;
 RECT 5.65 0.36 5.79 0.435 ;
 RECT 6.175 0.875 6.49 1.015 ;
 RECT 5.65 0.22 6.425 0.36 ;
 RECT 4.795 0.435 5.79 0.575 ;
 RECT 3.65 0.46 3.79 2.21 ;
 RECT 4.05 0.22 4.375 0.32 ;
 RECT 4.05 0.46 4.375 0.525 ;
 RECT 3.65 0.32 4.375 0.46 ;
 RECT 0.8 0.68 0.94 1.155 ;
 RECT 0.8 1.295 0.94 2.23 ;
 RECT 1.585 0.36 1.725 1.155 ;
 RECT 0.8 1.155 1.725 1.295 ;
 RECT 2.805 0.36 3.035 0.43 ;
 RECT 1.585 0.22 3.035 0.36 ;
 RECT 16.18 1.895 16.32 2.39 ;
 RECT 20.105 2.205 20.245 2.39 ;
 RECT 16.18 2.39 20.245 2.53 ;
 RECT 15.055 1.755 16.32 1.895 ;
 RECT 15.055 1.895 15.195 2.34 ;
 RECT 13.785 2.3 14.015 2.34 ;
 RECT 13.785 2.48 14.015 2.51 ;
 RECT 13.785 2.34 15.195 2.48 ;
 RECT 20.105 2.065 26.83 2.205 ;
 RECT 26.69 2.205 26.83 2.52 ;
 RECT 31.03 2.48 31.17 2.52 ;
 RECT 26.69 2.52 31.17 2.66 ;
 RECT 31.03 2.27 31.26 2.48 ;
 RECT 19.62 1.7 19.915 1.84 ;
 RECT 19.62 1.84 19.76 2.075 ;
 RECT 18.925 1.84 19.065 2.075 ;
 RECT 18.73 1.7 19.065 1.84 ;
 RECT 18.925 2.075 19.76 2.215 ;
 RECT 19.815 1.055 19.955 1.245 ;
 RECT 19.255 1.385 19.395 1.625 ;
 RECT 19.255 1.245 20.325 1.385 ;
 RECT 20.095 1.385 20.325 1.455 ;
 RECT 19.785 0.915 20.085 1.055 ;
 RECT 19.225 1.625 19.48 1.92 ;
 RECT 16.46 1.56 16.6 2.11 ;
 RECT 15.41 1.405 15.64 1.42 ;
 RECT 15.41 1.56 15.64 1.615 ;
 RECT 15.41 1.42 16.6 1.56 ;
 RECT 16.46 2.11 18.785 2.245 ;
 RECT 16.46 2.245 18.78 2.25 ;
 RECT 18.555 2.035 18.785 2.11 ;
 RECT 11.935 1.02 12.075 1.475 ;
 RECT 11.775 1.475 12.075 1.635 ;
 RECT 11.935 1.775 12.075 2.18 ;
 RECT 11.87 0.88 12.145 1.02 ;
 RECT 13 1.415 13.14 1.635 ;
 RECT 11.935 1.685 13.14 1.775 ;
 RECT 11.775 1.635 13.14 1.685 ;
 RECT 12.95 1.275 13.205 1.415 ;
 RECT 7.19 2.125 7.465 2.205 ;
 RECT 8.6 2.125 8.875 2.365 ;
 RECT 7.19 1.985 8.875 2.125 ;
 RECT 5.875 1.67 6.015 1.82 ;
 RECT 5.875 1.96 6.015 2.52 ;
 RECT 5.875 0.96 6.015 1.44 ;
 RECT 8.02 2.265 8.25 2.52 ;
 RECT 5.81 1.82 6.08 1.96 ;
 RECT 5.875 1.44 6.145 1.67 ;
 RECT 5.78 0.75 6.035 0.96 ;
 RECT 5.875 2.52 8.25 2.66 ;
 RECT 9.695 1.365 9.835 2.41 ;
 RECT 7 1.365 7.23 1.435 ;
 RECT 11.01 1.04 11.15 1.25 ;
 RECT 11.01 1.39 11.15 2.215 ;
 RECT 11.01 0.885 11.15 0.9 ;
 RECT 7 1.25 11.15 1.365 ;
 RECT 7 1.225 10.4 1.25 ;
 RECT 10.26 1.365 11.15 1.39 ;
 RECT 10.945 0.9 11.22 1.04 ;
 RECT 6.63 1.015 6.77 1.7 ;
 RECT 6.63 1.84 6.77 2.015 ;
 RECT 6.63 1.7 7.945 1.84 ;
 RECT 7.67 1.685 7.945 1.7 ;
 RECT 6.63 0.875 6.945 1.015 ;
 RECT 6.63 2.015 6.995 2.215 ;
 RECT 9.27 1.685 9.5 1.755 ;
 RECT 7.67 1.545 9.5 1.685 ;
 RECT 5.14 0.93 5.28 1.44 ;
 RECT 5.14 1.69 5.28 1.99 ;
 END
END RSDFFSRASRX2

MACRO RSDFFSRASX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 31.36 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 24.54 0.59 24.91 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 29.77 1.435 30.11 1.8 ;
 RECT 28.09 1.99 29.955 2.13 ;
 RECT 25.86 2.22 28.23 2.36 ;
 RECT 29.815 1.8 29.955 1.99 ;
 RECT 28.09 1.435 28.23 1.99 ;
 RECT 25.86 1.39 26 2.22 ;
 RECT 27.245 1.37 27.385 2.22 ;
 RECT 28.09 2.13 28.23 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 31.36 0.08 ;
 RECT 5.155 0.08 5.435 0.295 ;
 RECT 28.21 0.08 28.45 0.26 ;
 RECT 9.4 0.31 9.69 0.45 ;
 RECT 17.01 0.275 18.035 0.415 ;
 RECT 13.085 0.595 13.355 0.735 ;
 RECT 21.37 0.335 21.635 0.495 ;
 RECT 17.895 0.75 18.84 0.89 ;
 RECT 3.19 0.08 3.33 0.74 ;
 RECT 0.31 0.08 0.45 0.775 ;
 RECT 1.28 0.08 1.42 0.93 ;
 RECT 4.635 0.08 4.775 0.97 ;
 RECT 7.98 0.08 8.215 0.46 ;
 RECT 25.86 0.08 26 0.36 ;
 RECT 23.015 0.08 23.155 0.82 ;
 RECT 27.075 0.08 27.215 0.35 ;
 RECT 9.48 0.08 9.62 0.31 ;
 RECT 17.01 0.415 17.15 0.945 ;
 RECT 17.01 0.08 17.15 0.275 ;
 RECT 13.15 0.08 13.29 0.595 ;
 RECT 21.425 0.08 21.565 0.335 ;
 RECT 18.7 0.89 18.84 1.11 ;
 RECT 17.895 0.415 18.035 0.75 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.825 1.205 21.18 1.445 ;
 RECT 20.935 0.915 21.075 1.205 ;
 RECT 20.935 1.7 22.08 1.84 ;
 RECT 20.935 1.84 21.075 1.885 ;
 RECT 20.935 1.445 21.075 1.7 ;
 RECT 21.94 1.84 22.08 1.885 ;
 RECT 21.94 0.915 22.08 1.7 ;
 END
 ANTENNADIFFAREA 0.464 ;
 END QN

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.685 1.475 5.015 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.335 1.095 22.595 1.335 ;
 RECT 22.455 0.51 22.595 1.095 ;
 RECT 23.515 1.905 23.655 1.91 ;
 RECT 22.455 1.765 23.655 1.905 ;
 RECT 23.515 0.56 23.655 1.765 ;
 RECT 22.455 1.905 22.595 1.915 ;
 RECT 22.455 1.335 22.595 1.765 ;
 END
 ANTENNADIFFAREA 0.674 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.32 2.12 13.62 2.475 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.3 1.76 10.69 2.04 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.1 1.435 1.625 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.79 1.44 2.035 1.59 ;
 RECT 1.79 1.59 2.735 1.75 ;
 RECT 2.585 1.75 2.725 1.805 ;
 RECT 2.585 1.53 2.725 1.59 ;
 RECT 1.885 1.09 2.025 1.44 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.25 1.115 2.67 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 31.36 2.96 ;
 RECT 21.28 2.6 21.545 2.8 ;
 RECT 22.87 2.6 23.135 2.8 ;
 RECT 8.545 2.255 8.775 2.465 ;
 RECT 12.895 2.215 13.17 2.355 ;
 RECT 1.28 1.965 1.42 2.8 ;
 RECT 3.19 1.99 3.33 2.8 ;
 RECT 0.31 1.74 0.45 2.8 ;
 RECT 5.31 2.34 5.56 2.8 ;
 RECT 4.635 1.98 4.775 2.8 ;
 RECT 9.48 2.17 9.62 2.8 ;
 RECT 10.51 2.21 10.65 2.8 ;
 RECT 15.92 2.335 16.19 2.8 ;
 RECT 8.59 2.465 8.73 2.8 ;
 RECT 12.96 2.355 13.1 2.8 ;
 RECT 12.96 2.195 13.1 2.215 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 14.875 1.71 14.975 2.425 ;
 RECT 10.99 0.475 11.09 0.895 ;
 RECT 15.41 1.91 16.33 2.01 ;
 RECT 10.99 0.375 14.425 0.475 ;
 RECT 10.865 0.895 11.095 1.105 ;
 RECT 16.54 0.455 18.47 0.535 ;
 RECT 18.24 0.535 18.47 0.6 ;
 RECT 18.24 0.39 18.47 0.435 ;
 RECT 16.62 0.435 18.47 0.455 ;
 RECT 16.54 0.535 16.77 0.665 ;
 RECT 17.395 0.535 17.625 0.835 ;
 RECT 17.395 0.835 17.495 2.39 ;
 RECT 26.425 0.215 26.525 0.995 ;
 RECT 26.425 0.995 26.665 1.205 ;
 RECT 26.425 1.205 26.525 2 ;
 RECT 28.82 0.375 28.92 0.99 ;
 RECT 28.82 0.99 29.07 1.2 ;
 RECT 28.82 1.2 28.92 2.27 ;
 RECT 28.82 2.27 29.105 2.48 ;
 RECT 13.805 0.655 13.905 2.305 ;
 RECT 14.11 2.3 14.34 2.305 ;
 RECT 14.11 2.405 14.34 2.51 ;
 RECT 13.805 2.305 14.34 2.405 ;
 RECT 25.645 0.21 25.745 0.755 ;
 RECT 25.645 0.855 25.745 2.2 ;
 RECT 28.51 1.125 28.61 2.2 ;
 RECT 24.68 0.755 26.215 0.84 ;
 RECT 24.68 0.84 26.21 0.855 ;
 RECT 26.115 0.215 26.215 0.755 ;
 RECT 24.68 0.595 24.91 0.755 ;
 RECT 25.645 2.2 28.61 2.3 ;
 RECT 27.335 0.38 27.435 0.96 ;
 RECT 27.335 1.06 27.435 1.14 ;
 RECT 26.915 0.935 27.145 0.96 ;
 RECT 26.915 0.96 27.435 1.06 ;
 RECT 26.915 1.06 27.145 1.145 ;
 RECT 27.335 1.14 27.605 1.24 ;
 RECT 27.505 1.24 27.605 1.84 ;
 RECT 27.7 0.22 27.93 0.28 ;
 RECT 27.7 0.38 27.93 0.43 ;
 RECT 27.335 0.28 27.93 0.38 ;
 RECT 11.59 1.575 11.69 2.485 ;
 RECT 12.1 1.365 12.33 1.475 ;
 RECT 11.59 1.475 12.33 1.575 ;
 RECT 29.52 0.195 29.62 2.665 ;
 RECT 28.51 0.095 29.62 0.195 ;
 RECT 24.885 1.245 24.985 2.665 ;
 RECT 28.51 0.195 28.61 0.945 ;
 RECT 24.885 1.2 25.17 1.245 ;
 RECT 24.94 1.035 25.17 1.1 ;
 RECT 24.885 2.665 29.62 2.765 ;
 RECT 24.885 1.1 25.215 1.2 ;
 RECT 15.815 0.795 15.98 0.925 ;
 RECT 15.135 0.885 15.365 0.925 ;
 RECT 15.135 1.025 15.365 1.095 ;
 RECT 15.135 0.925 15.98 1.025 ;
 RECT 15.815 0.585 16.045 0.795 ;
 RECT 2.535 1.55 2.775 1.78 ;
 RECT 2.675 1.78 2.775 2.695 ;
 RECT 1.065 1.435 1.635 1.71 ;
 RECT 1.065 0.515 1.165 1.435 ;
 RECT 1.065 1.71 1.165 2.645 ;
 RECT 1.535 0.515 1.635 1.435 ;
 RECT 1.535 1.71 1.635 2.695 ;
 RECT 2.255 1.37 2.355 1.605 ;
 RECT 2.485 0.515 2.585 1.14 ;
 RECT 2.205 1.705 2.305 2.695 ;
 RECT 2.205 1.605 2.355 1.705 ;
 RECT 2.255 1.14 2.585 1.37 ;
 RECT 1.87 0.515 1.97 1.105 ;
 RECT 1.83 1.105 2.075 1.345 ;
 RECT 4.895 0.49 4.995 1.495 ;
 RECT 4.7 1.495 4.995 1.745 ;
 RECT 4.895 1.745 4.995 2.37 ;
 RECT 4.42 0.52 4.52 2.465 ;
 RECT 4.18 0.27 4.52 0.52 ;
 RECT 6.555 1.66 6.655 2.475 ;
 RECT 6.015 1.445 6.26 1.56 ;
 RECT 6.015 1.66 6.26 1.69 ;
 RECT 6.015 1.56 6.655 1.66 ;
 RECT 5.67 1.62 5.77 2.655 ;
 RECT 6.6 0.285 6.7 0.47 ;
 RECT 6.6 0.47 6.885 0.705 ;
 RECT 6.6 0.705 6.7 1.255 ;
 RECT 5.735 0.185 6.7 0.285 ;
 RECT 5.735 0.285 5.835 1.52 ;
 RECT 5.235 1.44 5.48 1.52 ;
 RECT 5.235 1.62 5.48 1.69 ;
 RECT 5.235 1.52 5.835 1.62 ;
 RECT 5.67 2.655 9.355 2.755 ;
 RECT 9.255 1.79 9.355 2.655 ;
 RECT 13.41 0.655 13.51 1.19 ;
 RECT 13.28 1.19 13.51 1.425 ;
 RECT 12.515 0.755 12.615 1.62 ;
 RECT 11.6 0.755 11.7 1.255 ;
 RECT 13.375 1.72 13.475 2.255 ;
 RECT 12.515 1.72 12.615 2.51 ;
 RECT 11.6 0.655 12.615 0.755 ;
 RECT 12.515 1.62 13.475 1.72 ;
 RECT 13.375 2.255 13.605 2.465 ;
 RECT 8.62 0.745 8.72 2.255 ;
 RECT 8.545 2.255 8.775 2.465 ;
 RECT 8.555 0.535 8.785 0.745 ;
 RECT 7.49 0.745 7.59 1.61 ;
 RECT 7.525 1.71 7.625 2.475 ;
 RECT 7.49 1.61 7.625 1.71 ;
 RECT 7.38 0.535 7.61 0.745 ;
 RECT 7.05 1.435 7.15 2.475 ;
 RECT 7.09 0.65 7.19 1.225 ;
 RECT 7.01 1.225 7.24 1.435 ;
 RECT 2.975 0.135 3.075 0.22 ;
 RECT 2.815 0.22 3.075 0.43 ;
 RECT 2.975 0.43 3.075 2.695 ;
 RECT 3.445 0.295 3.545 1.115 ;
 RECT 3.28 1.115 3.545 1.325 ;
 RECT 3.445 1.325 3.545 2.74 ;
 RECT 19.835 0.77 19.935 2.155 ;
 RECT 19.835 0.55 19.935 0.56 ;
 RECT 19.835 0.56 20.09 0.77 ;
 RECT 20.47 0.43 20.57 1.245 ;
 RECT 21.2 0.39 21.3 1.4 ;
 RECT 21.2 1.5 21.3 2.42 ;
 RECT 21.69 0.51 21.79 1.4 ;
 RECT 21.69 1.5 21.79 2.44 ;
 RECT 20.405 0.22 20.635 0.29 ;
 RECT 20.405 0.39 20.635 0.43 ;
 RECT 20.405 0.29 21.3 0.39 ;
 RECT 21.2 1.4 21.79 1.5 ;
 RECT 20.42 1.245 20.65 1.455 ;
 RECT 18.895 1.445 18.995 2.035 ;
 RECT 18.88 2.035 19.11 2.245 ;
 RECT 19.365 0.55 19.465 2.69 ;
 RECT 10.295 1.58 10.395 1.77 ;
 RECT 10.035 1.01 10.135 1.48 ;
 RECT 10.295 1.98 10.395 2.69 ;
 RECT 10.295 1.77 10.53 1.98 ;
 RECT 10.035 1.48 10.395 1.58 ;
 RECT 10.295 2.69 19.465 2.79 ;
 RECT 9.735 0.98 9.835 1.545 ;
 RECT 9.595 1.545 9.835 1.755 ;
 RECT 9.735 1.755 9.835 2.655 ;
 RECT 22.715 1.33 23.395 1.43 ;
 RECT 22.715 1.43 22.965 1.46 ;
 RECT 22.715 1.25 22.965 1.33 ;
 RECT 23.295 0.375 23.395 1.33 ;
 RECT 22.715 0.385 22.815 1.25 ;
 RECT 22.715 1.46 22.815 2.69 ;
 RECT 23.295 1.43 23.395 2.695 ;
 RECT 23.9 0.22 24.13 0.275 ;
 RECT 23.9 0.375 24.13 0.43 ;
 RECT 23.295 0.275 24.13 0.375 ;
 RECT 17.865 0.73 17.965 1.39 ;
 RECT 17.73 1.39 17.965 1.6 ;
 RECT 17.865 1.6 17.965 2.39 ;
 RECT 7.79 0.195 7.89 1.17 ;
 RECT 14.84 0.195 14.94 1.29 ;
 RECT 15.735 1.39 15.93 1.405 ;
 RECT 8.03 1.27 8.13 2.255 ;
 RECT 7.79 0.095 14.945 0.195 ;
 RECT 14.84 1.29 15.93 1.39 ;
 RECT 8.03 2.255 8.26 2.465 ;
 RECT 7.79 1.17 8.13 1.27 ;
 RECT 15.735 1.405 15.965 1.615 ;
 RECT 26.12 1.245 26.22 2.02 ;
 RECT 25.99 1.035 26.22 1.245 ;
 RECT 16.23 0.105 19.055 0.205 ;
 RECT 16.23 0.205 16.33 1.91 ;
 RECT 18.955 0.205 19.055 1.265 ;
 RECT 15.41 1.71 15.51 1.91 ;
 RECT 14.325 1.61 15.51 1.71 ;
 RECT 14.325 0.475 14.425 1.61 ;
 LAYER CO ;
 RECT 15.785 1.445 15.915 1.575 ;
 RECT 26.04 1.075 26.17 1.205 ;
 RECT 10.915 0.935 11.045 1.065 ;
 RECT 26.965 0.975 27.095 1.105 ;
 RECT 17.445 0.665 17.575 0.795 ;
 RECT 26.485 1.035 26.615 1.165 ;
 RECT 28.925 2.31 29.055 2.44 ;
 RECT 14.16 2.34 14.29 2.47 ;
 RECT 24.73 0.635 24.86 0.765 ;
 RECT 27.75 0.26 27.88 0.39 ;
 RECT 12.15 1.405 12.28 1.535 ;
 RECT 24.99 1.075 25.12 1.205 ;
 RECT 15.185 0.925 15.315 1.055 ;
 RECT 4.76 1.55 4.89 1.68 ;
 RECT 1.285 0.735 1.415 0.865 ;
 RECT 1.29 1.51 1.42 1.64 ;
 RECT 0.815 0.735 0.945 0.865 ;
 RECT 3.195 2.31 3.325 2.44 ;
 RECT 1.285 2.015 1.415 2.145 ;
 RECT 1.89 1.155 2.02 1.285 ;
 RECT 3.195 2.05 3.325 2.18 ;
 RECT 2.59 1.6 2.72 1.73 ;
 RECT 3.665 2.01 3.795 2.14 ;
 RECT 3.665 0.735 3.795 0.865 ;
 RECT 2.425 2.075 2.555 2.205 ;
 RECT 1.285 2.275 1.415 2.405 ;
 RECT 3.195 0.545 3.325 0.675 ;
 RECT 3.665 1.75 3.795 1.88 ;
 RECT 0.815 2.015 0.945 2.145 ;
 RECT 2.23 0.735 2.36 0.865 ;
 RECT 2.41 1.19 2.54 1.32 ;
 RECT 11.34 2.015 11.47 2.145 ;
 RECT 27.08 0.12 27.21 0.25 ;
 RECT 26.645 1.485 26.775 1.615 ;
 RECT 29.04 1.465 29.17 1.595 ;
 RECT 19.585 1.705 19.715 1.835 ;
 RECT 29.04 0.595 29.17 0.725 ;
 RECT 12.965 2.225 13.095 2.355 ;
 RECT 21.945 0.975 22.075 1.105 ;
 RECT 22.935 2.64 23.065 2.77 ;
 RECT 4.17 2.115 4.3 2.245 ;
 RECT 21.43 0.36 21.56 0.49 ;
 RECT 23.52 0.63 23.65 0.76 ;
 RECT 27.585 0.595 27.715 0.725 ;
 RECT 6.705 0.525 6.835 0.655 ;
 RECT 7.745 1.67 7.875 1.8 ;
 RECT 28.095 1.49 28.225 1.62 ;
 RECT 6.35 0.88 6.48 1.01 ;
 RECT 15.095 1.87 15.225 2 ;
 RECT 9 2.195 9.13 2.325 ;
 RECT 8.035 0.32 8.165 0.45 ;
 RECT 25.865 0.135 25.995 0.265 ;
 RECT 5.295 1.495 5.425 1.625 ;
 RECT 5.245 0.745 5.375 0.875 ;
 RECT 5.115 1.995 5.245 2.125 ;
 RECT 12.265 1.995 12.395 2.125 ;
 RECT 0.315 0.59 0.445 0.72 ;
 RECT 11.82 2.07 11.95 2.2 ;
 RECT 14.59 0.595 14.72 0.725 ;
 RECT 6.07 1.49 6.2 1.62 ;
 RECT 13.33 1.235 13.46 1.365 ;
 RECT 22.46 1.725 22.59 1.855 ;
 RECT 0.315 2.085 0.445 2.215 ;
 RECT 10.025 2.215 10.155 2.345 ;
 RECT 18.12 1.035 18.25 1.165 ;
 RECT 18.705 0.91 18.835 1.04 ;
 RECT 10.515 2.28 10.645 2.41 ;
 RECT 23.02 0.62 23.15 0.75 ;
 RECT 6.305 2.105 6.435 2.235 ;
 RECT 7.27 2.025 7.4 2.155 ;
 RECT 5.225 0.145 5.355 0.275 ;
 RECT 14.59 1.9 14.72 2.03 ;
 RECT 0.315 2.345 0.445 2.475 ;
 RECT 5.38 2.345 5.51 2.475 ;
 RECT 26.645 0.435 26.775 0.565 ;
 RECT 20.94 1.705 21.07 1.835 ;
 RECT 10.295 1.23 10.425 1.36 ;
 RECT 19.115 1.705 19.245 1.835 ;
 RECT 9.485 2.245 9.615 2.375 ;
 RECT 6.82 0.88 6.95 1.01 ;
 RECT 17.145 1.835 17.275 1.965 ;
 RECT 17.015 0.765 17.145 0.895 ;
 RECT 4.64 0.74 4.77 0.87 ;
 RECT 28.26 0.12 28.39 0.25 ;
 RECT 22.46 0.62 22.59 0.75 ;
 RECT 15.99 2.38 16.12 2.51 ;
 RECT 12.265 0.885 12.395 1.015 ;
 RECT 25.395 1.425 25.525 1.555 ;
 RECT 0.315 0.33 0.445 0.46 ;
 RECT 20.18 0.92 20.31 1.05 ;
 RECT 25.865 1.475 25.995 1.605 ;
 RECT 14.065 0.875 14.195 1.005 ;
 RECT 5.955 0.79 6.085 0.92 ;
 RECT 18.085 1.835 18.215 1.965 ;
 RECT 6.8 2.07 6.93 2.2 ;
 RECT 29.82 1.475 29.95 1.605 ;
 RECT 21.945 1.705 22.075 1.835 ;
 RECT 23.52 1.71 23.65 1.84 ;
 RECT 20.94 0.975 21.07 1.105 ;
 RECT 4.17 0.74 4.3 0.87 ;
 RECT 5.89 1.825 6.02 1.955 ;
 RECT 14.065 1.945 14.195 2.075 ;
 RECT 4.64 2.05 4.77 2.18 ;
 RECT 25.145 0.505 25.275 0.635 ;
 RECT 20.06 1.705 20.19 1.835 ;
 RECT 21.345 2.64 21.475 2.77 ;
 RECT 27.725 1.405 27.855 1.535 ;
 RECT 11.345 0.905 11.475 1.035 ;
 RECT 4.24 0.325 4.37 0.455 ;
 RECT 9.485 0.315 9.615 0.445 ;
 RECT 11.82 0.905 11.95 1.035 ;
 RECT 15.095 0.595 15.225 0.725 ;
 RECT 13.155 0.595 13.285 0.725 ;
 RECT 27.25 1.445 27.38 1.575 ;
 RECT 0.315 1.825 0.445 1.955 ;
 RECT 13.425 2.295 13.555 2.425 ;
 RECT 8.595 2.295 8.725 2.425 ;
 RECT 8.605 0.575 8.735 0.705 ;
 RECT 7.43 0.575 7.56 0.705 ;
 RECT 8.08 2.295 8.21 2.425 ;
 RECT 7.06 1.265 7.19 1.395 ;
 RECT 2.865 0.26 2.995 0.39 ;
 RECT 3.33 1.155 3.46 1.285 ;
 RECT 22.785 1.29 22.915 1.42 ;
 RECT 20.47 1.285 20.6 1.415 ;
 RECT 18.29 0.43 18.42 0.56 ;
 RECT 19.91 0.6 20.04 0.73 ;
 RECT 20.455 0.26 20.585 0.39 ;
 RECT 18.93 2.075 19.06 2.205 ;
 RECT 10.35 1.81 10.48 1.94 ;
 RECT 9.645 1.585 9.775 1.715 ;
 RECT 23.95 0.26 24.08 0.39 ;
 RECT 28.89 1.03 29.02 1.16 ;
 RECT 16.59 0.495 16.72 0.625 ;
 RECT 17.78 1.43 17.91 1.56 ;
 RECT 15.865 0.625 15.995 0.755 ;
 LAYER M1 ;
 RECT 3.28 1.29 3.51 1.325 ;
 RECT 27.58 0.73 27.72 1.04 ;
 RECT 27.72 1.18 27.86 1.605 ;
 RECT 27.515 0.59 27.79 0.73 ;
 RECT 28.84 0.99 29.07 1.04 ;
 RECT 27.58 1.04 29.07 1.18 ;
 RECT 28.84 1.18 29.07 1.2 ;
 RECT 27.7 0.29 28.07 0.43 ;
 RECT 27.93 0.43 28.07 0.71 ;
 RECT 27.7 0.22 27.93 0.29 ;
 RECT 29.35 0.85 29.49 1.385 ;
 RECT 29.035 1.525 29.175 1.73 ;
 RECT 27.93 0.71 29.49 0.85 ;
 RECT 29.035 0.51 29.175 0.71 ;
 RECT 29.035 1.385 29.49 1.525 ;
 RECT 24.94 1.225 25.17 1.245 ;
 RECT 24.94 1.195 25.53 1.225 ;
 RECT 25.08 1.015 25.39 1.035 ;
 RECT 24.94 1.035 25.39 1.055 ;
 RECT 25.215 0.64 25.355 1.015 ;
 RECT 25.39 1.225 25.53 1.75 ;
 RECT 25.095 0.5 25.355 0.64 ;
 RECT 25.99 1.035 26.22 1.055 ;
 RECT 25.99 1.195 26.22 1.245 ;
 RECT 24.94 1.055 26.22 1.195 ;
 RECT 26.96 1.145 27.1 1.345 ;
 RECT 26.64 1.485 26.78 1.76 ;
 RECT 26.96 0.73 27.1 0.935 ;
 RECT 26.64 0.355 26.78 0.59 ;
 RECT 26.64 1.345 27.1 1.485 ;
 RECT 26.915 0.935 27.145 1.145 ;
 RECT 26.64 0.59 27.1 0.73 ;
 RECT 23.9 0.36 24.13 0.43 ;
 RECT 25.495 0.36 25.635 0.565 ;
 RECT 23.9 0.22 25.635 0.36 ;
 RECT 26.235 0.705 26.375 0.75 ;
 RECT 26.36 0.995 26.665 1.205 ;
 RECT 26.36 0.89 26.5 0.995 ;
 RECT 26.235 0.75 26.5 0.89 ;
 RECT 25.495 0.565 26.375 0.705 ;
 RECT 19.135 0.775 19.275 1.405 ;
 RECT 19.86 0.56 20.09 0.635 ;
 RECT 18.115 1.405 19.275 1.545 ;
 RECT 18.115 1.545 18.255 1.83 ;
 RECT 18.115 1.17 18.255 1.405 ;
 RECT 17.07 1.83 18.32 1.97 ;
 RECT 18.045 1.03 18.325 1.17 ;
 RECT 22.055 0.36 22.195 0.635 ;
 RECT 19.135 0.635 22.195 0.775 ;
 RECT 22.735 0.36 22.875 1.25 ;
 RECT 22.735 1.25 22.965 1.46 ;
 RECT 22.055 0.22 22.875 0.36 ;
 RECT 18.24 0.28 20.635 0.42 ;
 RECT 18.24 0.42 18.47 0.6 ;
 RECT 20.405 0.22 20.635 0.28 ;
 RECT 20.405 0.42 20.635 0.43 ;
 RECT 17.395 0.57 17.625 0.95 ;
 RECT 15.09 0.525 15.23 0.885 ;
 RECT 15.09 1.095 15.23 2.065 ;
 RECT 15.09 0.885 15.365 1.095 ;
 RECT 11.815 1.04 11.955 2.34 ;
 RECT 11.815 0.895 11.955 0.9 ;
 RECT 12.61 1.845 12.75 2.34 ;
 RECT 11.745 0.9 12.02 1.04 ;
 RECT 11.815 2.34 12.75 2.48 ;
 RECT 14.06 1.845 14.2 2.145 ;
 RECT 14.06 0.765 14.2 1.705 ;
 RECT 12.61 1.72 14.725 1.845 ;
 RECT 12.63 1.705 14.725 1.72 ;
 RECT 14.585 0.525 14.725 1.705 ;
 RECT 14.585 1.845 14.725 2.11 ;
 RECT 15.815 0.585 16.77 0.63 ;
 RECT 16.54 0.63 16.77 0.665 ;
 RECT 16.54 0.455 16.77 0.49 ;
 RECT 15.84 0.49 16.77 0.585 ;
 RECT 15.815 0.63 16.045 0.795 ;
 RECT 8.03 2.255 8.26 2.51 ;
 RECT 5.95 1.67 6.09 1.82 ;
 RECT 5.95 1.96 6.09 2.51 ;
 RECT 5.95 0.5 6.09 1.44 ;
 RECT 5.95 1.44 6.205 1.67 ;
 RECT 5.82 1.82 6.13 1.96 ;
 RECT 5.95 2.51 8.26 2.65 ;
 RECT 3.945 0.875 4.085 1.195 ;
 RECT 3.945 1.335 4.085 2.11 ;
 RECT 3.945 2.25 4.085 2.255 ;
 RECT 3.945 0.735 4.37 0.875 ;
 RECT 3.945 2.11 4.37 2.25 ;
 RECT 3.945 1.195 5.055 1.335 ;
 RECT 4.915 0.6 5.055 1.195 ;
 RECT 6.345 0.36 6.485 2.035 ;
 RECT 5.66 0.36 5.8 0.46 ;
 RECT 5.66 0.22 6.485 0.36 ;
 RECT 6.3 2.17 6.44 2.305 ;
 RECT 4.915 0.46 5.8 0.6 ;
 RECT 6.3 2.035 6.485 2.17 ;
 RECT 7.095 0.895 11.095 1.035 ;
 RECT 10.865 1.035 11.095 1.105 ;
 RECT 7.095 0.66 7.235 0.895 ;
 RECT 6.635 0.52 7.235 0.66 ;
 RECT 3.66 0.46 3.8 2.21 ;
 RECT 4.13 0.22 4.495 0.32 ;
 RECT 4.13 0.46 4.495 0.525 ;
 RECT 3.66 0.32 4.495 0.46 ;
 RECT 17.385 1.23 17.525 1.42 ;
 RECT 15.535 1.09 17.525 1.23 ;
 RECT 15.535 0.385 15.675 1.09 ;
 RECT 13.525 0.385 13.665 0.88 ;
 RECT 13.525 0.255 15.675 0.385 ;
 RECT 13.525 0.245 15.67 0.255 ;
 RECT 12.61 0.88 13.665 1.01 ;
 RECT 12.61 1.01 13.645 1.02 ;
 RECT 12.61 0.675 12.75 0.88 ;
 RECT 7.38 0.605 12.75 0.675 ;
 RECT 7.38 0.675 12.04 0.745 ;
 RECT 11.9 0.535 12.75 0.605 ;
 RECT 8.555 0.535 8.785 0.605 ;
 RECT 7.38 0.535 7.61 0.605 ;
 RECT 17.73 1.39 17.96 1.42 ;
 RECT 17.385 1.42 17.96 1.56 ;
 RECT 17.73 1.56 17.96 1.6 ;
 RECT 0.81 0.68 0.95 1.155 ;
 RECT 0.81 1.295 0.95 2.23 ;
 RECT 1.595 0.36 1.735 1.155 ;
 RECT 0.81 1.155 1.735 1.295 ;
 RECT 2.815 0.36 3.045 0.43 ;
 RECT 1.595 0.22 3.045 0.36 ;
 RECT 19.945 1.7 20.24 1.84 ;
 RECT 19.945 1.84 20.085 2.075 ;
 RECT 19.25 1.84 19.39 2.075 ;
 RECT 19.055 1.7 19.39 1.84 ;
 RECT 19.25 2.075 20.085 2.215 ;
 RECT 20.14 1.055 20.28 1.245 ;
 RECT 19.58 1.385 19.72 1.625 ;
 RECT 20.42 1.385 20.65 1.455 ;
 RECT 19.58 1.245 20.65 1.385 ;
 RECT 20.11 0.915 20.41 1.055 ;
 RECT 19.55 1.625 19.805 1.92 ;
 RECT 16.785 1.56 16.925 2.11 ;
 RECT 16.785 2.11 19.11 2.245 ;
 RECT 16.785 2.245 19.105 2.25 ;
 RECT 18.88 2.035 19.11 2.11 ;
 RECT 15.735 1.405 15.965 1.42 ;
 RECT 15.735 1.56 15.965 1.615 ;
 RECT 15.735 1.42 16.925 1.56 ;
 RECT 20.65 2.205 20.79 2.39 ;
 RECT 16.505 1.895 16.645 2.39 ;
 RECT 16.505 2.39 20.79 2.53 ;
 RECT 15.38 1.755 16.645 1.895 ;
 RECT 15.38 1.895 15.52 2.34 ;
 RECT 14.11 2.3 14.34 2.34 ;
 RECT 14.11 2.48 14.34 2.51 ;
 RECT 14.11 2.34 15.52 2.48 ;
 RECT 20.65 2.065 24.675 2.205 ;
 RECT 24.535 2.205 24.675 2.52 ;
 RECT 28.875 2.48 29.015 2.52 ;
 RECT 24.535 2.52 29.015 2.66 ;
 RECT 28.875 2.27 29.105 2.48 ;
 RECT 12.1 1.365 12.4 1.42 ;
 RECT 12.1 1.56 12.4 1.575 ;
 RECT 12.26 1.02 12.4 1.365 ;
 RECT 12.26 1.575 12.4 2.18 ;
 RECT 12.19 0.88 12.465 1.02 ;
 RECT 12.1 1.42 13.465 1.56 ;
 RECT 13.325 1.165 13.465 1.42 ;
 RECT 5.155 1.475 5.5 1.63 ;
 RECT 5.155 1.63 5.295 1.99 ;
 RECT 5.195 0.88 5.335 1.475 ;
 RECT 5.045 1.99 5.295 2.13 ;
 RECT 5.195 0.74 5.515 0.88 ;
 RECT 7.2 2.115 7.475 2.205 ;
 RECT 8.925 2.115 9.2 2.375 ;
 RECT 7.2 1.975 9.2 2.115 ;
 RECT 6.64 0.875 6.955 1.08 ;
 RECT 6.64 1.08 6.78 1.665 ;
 RECT 6.64 1.805 6.78 2.015 ;
 RECT 6.64 1.685 7.95 1.805 ;
 RECT 6.765 0.8 6.955 0.875 ;
 RECT 6.64 2.015 7.005 2.215 ;
 RECT 9.595 1.685 9.825 1.755 ;
 RECT 6.64 1.665 9.825 1.685 ;
 RECT 7.68 1.545 9.825 1.665 ;
 RECT 10.02 1.365 10.16 2.415 ;
 RECT 7.01 1.365 7.24 1.435 ;
 RECT 11.335 1.04 11.475 1.25 ;
 RECT 11.335 1.39 11.475 2.215 ;
 RECT 11.335 0.885 11.475 0.9 ;
 RECT 7.01 1.25 11.475 1.365 ;
 RECT 7.01 1.225 10.725 1.25 ;
 RECT 10.585 1.365 11.475 1.39 ;
 RECT 11.27 0.9 11.545 1.04 ;
 RECT 2.88 0.87 3.02 1.15 ;
 RECT 2.88 1.29 3.02 2.07 ;
 RECT 2.175 0.73 3.02 0.87 ;
 RECT 2.37 2.07 3.02 2.21 ;
 RECT 2.88 1.15 3.51 1.29 ;
 RECT 3.28 1.115 3.51 1.15 ;
 END
END RSDFFSRASX1

MACRO RSDFFSRASX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 34.24 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 27.395 0.59 27.765 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 32.625 1.435 32.965 1.8 ;
 RECT 30.945 1.99 32.81 2.13 ;
 RECT 28.715 2.22 31.085 2.36 ;
 RECT 30.945 1.435 31.085 1.99 ;
 RECT 32.67 1.8 32.81 1.99 ;
 RECT 28.715 1.39 28.855 2.22 ;
 RECT 30.1 1.37 30.24 2.22 ;
 RECT 30.945 2.13 31.085 2.22 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 34.24 0.08 ;
 RECT 9.775 0.31 10.065 0.45 ;
 RECT 13.46 0.595 13.73 0.735 ;
 RECT 17.385 0.275 18.41 0.415 ;
 RECT 22.71 0.335 22.975 0.495 ;
 RECT 21.715 0.335 21.98 0.495 ;
 RECT 18.27 0.75 19.215 0.89 ;
 RECT 4.515 0.08 4.655 0.97 ;
 RECT 3.18 0.08 3.32 0.74 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 0.93 ;
 RECT 5.145 0.08 5.425 0.295 ;
 RECT 7.97 0.08 8.205 0.46 ;
 RECT 28.715 0.08 28.855 0.36 ;
 RECT 24.515 0.08 24.655 0.82 ;
 RECT 25.57 0.08 25.71 0.82 ;
 RECT 31.065 0.08 31.305 0.26 ;
 RECT 29.93 0.08 30.07 0.35 ;
 RECT 9.855 0.08 9.995 0.31 ;
 RECT 13.525 0.08 13.665 0.595 ;
 RECT 17.385 0.415 17.525 0.945 ;
 RECT 17.385 0.08 17.525 0.275 ;
 RECT 22.765 0.08 22.905 0.335 ;
 RECT 21.77 0.08 21.91 0.335 ;
 RECT 19.075 0.89 19.215 1.11 ;
 RECT 18.27 0.415 18.41 0.75 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.6 1.475 4.93 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.915 1.16 13.325 1.485 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.675 1.615 11 2.04 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.435 1.615 1.71 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.78 1.59 2.725 1.75 ;
 RECT 1.875 1.09 2.015 1.44 ;
 RECT 1.78 1.44 2.025 1.59 ;
 RECT 2.575 1.75 2.715 1.805 ;
 RECT 2.575 1.53 2.715 1.59 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.24 1.115 2.66 1.375 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 34.24 2.96 ;
 RECT 8.78 2.265 9.01 2.475 ;
 RECT 13.27 2.215 13.545 2.355 ;
 RECT 1.27 1.965 1.41 2.8 ;
 RECT 3.18 1.99 3.32 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 4.49 1.98 4.63 2.8 ;
 RECT 5.18 2.34 5.43 2.8 ;
 RECT 9.855 1.98 9.995 2.8 ;
 RECT 10.885 2.33 11.025 2.8 ;
 RECT 16.295 2.335 16.565 2.8 ;
 RECT 22.62 2.6 22.885 2.8 ;
 RECT 21.625 2.6 21.89 2.8 ;
 RECT 24.37 2.6 24.635 2.8 ;
 RECT 25.425 2.6 25.69 2.8 ;
 RECT 8.825 2.475 8.965 2.8 ;
 RECT 13.335 2.355 13.475 2.8 ;
 RECT 13.335 2.195 13.475 2.215 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 21.17 1.205 21.47 1.445 ;
 RECT 21.28 0.915 21.42 1.205 ;
 RECT 22.285 1.84 22.425 1.885 ;
 RECT 22.285 0.915 22.425 1.7 ;
 RECT 23.28 1.84 23.42 1.885 ;
 RECT 23.28 0.915 23.42 1.7 ;
 RECT 21.28 1.7 23.47 1.84 ;
 RECT 21.28 1.84 21.42 1.885 ;
 RECT 21.28 1.445 21.42 1.7 ;
 END
 ANTENNADIFFAREA 0.883 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 23.835 1.095 24.095 1.335 ;
 RECT 23.955 0.51 24.095 1.095 ;
 RECT 25.015 1.905 25.155 1.91 ;
 RECT 25.015 0.56 25.155 1.765 ;
 RECT 26.07 1.905 26.21 1.91 ;
 RECT 26.07 0.56 26.21 1.765 ;
 RECT 23.955 1.905 24.095 1.915 ;
 RECT 23.955 1.335 24.095 1.765 ;
 RECT 23.955 1.765 26.21 1.905 ;
 END
 ANTENNADIFFAREA 0.827 ;
 END Q

 OBS
 LAYER PO ;
 RECT 16.915 0.535 17.145 0.665 ;
 RECT 17.77 0.535 18 0.835 ;
 RECT 17.77 0.835 17.87 2.39 ;
 RECT 29.28 0.215 29.38 0.995 ;
 RECT 29.28 0.995 29.52 1.205 ;
 RECT 29.28 1.205 29.38 2 ;
 RECT 31.675 0.375 31.775 0.99 ;
 RECT 31.675 0.99 31.925 1.2 ;
 RECT 31.675 1.2 31.775 2.27 ;
 RECT 31.675 2.27 31.96 2.48 ;
 RECT 14.18 0.655 14.28 2.305 ;
 RECT 14.485 2.3 14.715 2.305 ;
 RECT 14.485 2.405 14.715 2.51 ;
 RECT 14.18 2.305 14.715 2.405 ;
 RECT 28.5 0.855 28.6 2.2 ;
 RECT 31.365 1.125 31.465 2.2 ;
 RECT 27.535 0.755 29.07 0.84 ;
 RECT 27.535 0.84 29.065 0.855 ;
 RECT 28.97 0.215 29.07 0.755 ;
 RECT 28.5 0.21 28.6 0.755 ;
 RECT 27.535 0.595 27.765 0.755 ;
 RECT 28.5 2.2 31.465 2.3 ;
 RECT 12.89 1.44 12.99 1.62 ;
 RECT 12.89 1.72 12.99 2.51 ;
 RECT 12.89 0.755 12.99 1.23 ;
 RECT 11.975 0.755 12.075 1.255 ;
 RECT 12.89 1.62 13.85 1.72 ;
 RECT 13.75 1.72 13.85 2.355 ;
 RECT 12.89 1.23 13.145 1.44 ;
 RECT 11.975 0.655 12.99 0.755 ;
 RECT 30.19 0.38 30.29 0.96 ;
 RECT 30.19 1.06 30.29 1.14 ;
 RECT 29.77 0.935 30 0.96 ;
 RECT 29.77 0.96 30.29 1.06 ;
 RECT 29.77 1.06 30 1.145 ;
 RECT 30.19 1.14 30.46 1.24 ;
 RECT 30.36 1.24 30.46 1.84 ;
 RECT 30.555 0.22 30.785 0.28 ;
 RECT 30.555 0.38 30.785 0.43 ;
 RECT 30.19 0.28 30.785 0.38 ;
 RECT 11.965 1.685 12.065 2.485 ;
 RECT 12.48 1.48 12.71 1.585 ;
 RECT 12.48 1.685 12.71 1.69 ;
 RECT 11.965 1.585 12.71 1.685 ;
 RECT 32.375 0.195 32.475 2.665 ;
 RECT 31.365 0.095 32.475 0.195 ;
 RECT 27.74 1.245 27.84 2.665 ;
 RECT 31.365 0.195 31.465 0.945 ;
 RECT 27.74 1.2 28.025 1.245 ;
 RECT 27.795 1.035 28.025 1.1 ;
 RECT 27.74 2.665 32.475 2.765 ;
 RECT 27.74 1.1 28.07 1.2 ;
 RECT 16.19 0.795 16.355 0.925 ;
 RECT 15.51 0.885 15.74 0.925 ;
 RECT 15.51 1.025 15.74 1.095 ;
 RECT 15.51 0.925 16.355 1.025 ;
 RECT 16.19 0.585 16.42 0.795 ;
 RECT 2.525 1.55 2.765 1.78 ;
 RECT 2.665 1.78 2.765 2.695 ;
 RECT 1.055 1.435 1.625 1.71 ;
 RECT 1.055 0.515 1.155 1.435 ;
 RECT 1.055 1.71 1.155 2.645 ;
 RECT 1.525 0.515 1.625 1.435 ;
 RECT 1.525 1.71 1.625 2.695 ;
 RECT 2.245 1.37 2.345 1.605 ;
 RECT 2.475 0.515 2.575 1.14 ;
 RECT 2.195 1.705 2.295 2.695 ;
 RECT 2.195 1.605 2.345 1.705 ;
 RECT 2.245 1.14 2.575 1.37 ;
 RECT 1.86 0.515 1.96 1.105 ;
 RECT 1.82 1.105 2.065 1.345 ;
 RECT 7.48 0.715 7.58 1.61 ;
 RECT 7.515 1.71 7.615 2.475 ;
 RECT 7.48 1.61 7.615 1.71 ;
 RECT 7.36 0.485 7.6 0.715 ;
 RECT 4.275 0.52 4.375 2.465 ;
 RECT 4.13 0.27 4.375 0.52 ;
 RECT 13.785 0.655 13.885 1.195 ;
 RECT 13.655 1.195 13.885 1.43 ;
 RECT 4.81 0.49 4.91 1.495 ;
 RECT 4.615 1.495 4.91 1.745 ;
 RECT 4.81 1.745 4.91 2.37 ;
 RECT 8.785 0.735 8.885 2.265 ;
 RECT 8.78 2.265 9.01 2.475 ;
 RECT 8.72 0.525 8.95 0.735 ;
 RECT 5.635 2.655 9.73 2.755 ;
 RECT 5.635 1.62 5.735 2.655 ;
 RECT 5.635 0.285 5.735 1.52 ;
 RECT 6.48 0.285 6.58 0.485 ;
 RECT 9.63 1.79 9.73 2.655 ;
 RECT 5.18 1.44 5.425 1.52 ;
 RECT 5.18 1.52 5.735 1.62 ;
 RECT 5.18 1.62 5.425 1.69 ;
 RECT 5.635 0.185 6.58 0.285 ;
 RECT 6.48 0.485 6.795 0.695 ;
 RECT 6.48 0.695 6.58 1.255 ;
 RECT 6.545 1.66 6.645 2.475 ;
 RECT 5.915 1.45 6.145 1.56 ;
 RECT 5.915 1.56 6.645 1.66 ;
 RECT 7.04 1.435 7.14 2.475 ;
 RECT 7.08 0.65 7.18 1.225 ;
 RECT 7 1.225 7.23 1.435 ;
 RECT 2.965 0.135 3.065 0.22 ;
 RECT 2.805 0.22 3.065 0.43 ;
 RECT 2.965 0.43 3.065 2.695 ;
 RECT 3.435 0.295 3.535 1.115 ;
 RECT 3.27 1.115 3.535 1.325 ;
 RECT 3.435 1.325 3.535 2.74 ;
 RECT 20.21 0.77 20.31 2.155 ;
 RECT 20.21 0.55 20.31 0.56 ;
 RECT 20.21 0.56 20.465 0.77 ;
 RECT 20.78 0.195 21.01 0.43 ;
 RECT 21.545 0.195 21.645 1.4 ;
 RECT 21.545 1.5 21.645 2.42 ;
 RECT 22.54 0.54 22.64 1.4 ;
 RECT 21.545 1.4 23.13 1.5 ;
 RECT 23.03 0.51 23.13 1.4 ;
 RECT 23.03 1.5 23.13 2.44 ;
 RECT 22.54 1.5 22.64 2.42 ;
 RECT 22.035 0.51 22.135 1.4 ;
 RECT 22.035 1.5 22.135 2.44 ;
 RECT 20.845 0.43 20.945 1.245 ;
 RECT 20.795 1.245 21.025 1.455 ;
 RECT 20.78 0.095 21.645 0.195 ;
 RECT 19.27 1.445 19.37 2.035 ;
 RECT 19.255 2.035 19.485 2.245 ;
 RECT 19.74 0.55 19.84 2.69 ;
 RECT 10.67 1.58 10.77 1.62 ;
 RECT 10.41 1.01 10.51 1.48 ;
 RECT 10.67 1.83 10.77 2.69 ;
 RECT 10.67 1.62 10.915 1.83 ;
 RECT 10.41 1.48 10.77 1.58 ;
 RECT 10.67 2.69 19.84 2.79 ;
 RECT 10.11 0.98 10.21 1.545 ;
 RECT 9.97 1.545 10.21 1.755 ;
 RECT 10.11 1.755 10.21 2.51 ;
 RECT 25.85 0.335 25.95 1.33 ;
 RECT 24.215 1.25 24.465 1.33 ;
 RECT 24.215 1.43 24.465 1.46 ;
 RECT 24.215 1.33 25.95 1.43 ;
 RECT 24.215 0.385 24.315 1.25 ;
 RECT 24.215 1.46 24.315 2.69 ;
 RECT 24.795 0.385 24.895 1.33 ;
 RECT 24.795 1.43 24.895 2.695 ;
 RECT 25.27 0.385 25.37 1.33 ;
 RECT 25.27 1.43 25.37 2.69 ;
 RECT 25.85 1.43 25.95 2.695 ;
 RECT 26.755 0.22 26.985 0.235 ;
 RECT 26.755 0.335 26.985 0.43 ;
 RECT 25.85 0.235 26.985 0.335 ;
 RECT 18.24 0.73 18.34 1.39 ;
 RECT 18.105 1.39 18.34 1.6 ;
 RECT 18.24 1.6 18.34 2.39 ;
 RECT 7.78 0.195 7.88 1.17 ;
 RECT 15.215 0.195 15.315 1.29 ;
 RECT 16.11 1.39 16.305 1.405 ;
 RECT 8.02 1.27 8.12 2.265 ;
 RECT 7.78 0.095 15.315 0.195 ;
 RECT 15.215 1.29 16.305 1.39 ;
 RECT 8.02 2.265 8.25 2.475 ;
 RECT 7.78 1.17 8.12 1.27 ;
 RECT 16.11 1.405 16.34 1.615 ;
 RECT 28.975 1.245 29.075 2.02 ;
 RECT 28.845 1.035 29.075 1.245 ;
 RECT 16.605 0.105 19.43 0.205 ;
 RECT 16.605 0.205 16.705 1.91 ;
 RECT 19.33 0.205 19.43 1.265 ;
 RECT 15.785 1.71 15.885 1.91 ;
 RECT 14.7 1.61 15.885 1.71 ;
 RECT 14.7 0.475 14.8 1.61 ;
 RECT 15.25 1.71 15.35 2.425 ;
 RECT 11.365 0.475 11.465 0.895 ;
 RECT 15.785 1.91 16.705 2.01 ;
 RECT 11.365 0.375 14.8 0.475 ;
 RECT 11.24 0.895 11.47 1.105 ;
 RECT 16.915 0.455 18.845 0.535 ;
 RECT 18.615 0.535 18.845 0.6 ;
 RECT 18.615 0.39 18.845 0.435 ;
 RECT 16.995 0.435 18.845 0.455 ;
 LAYER CO ;
 RECT 12.965 1.27 13.095 1.4 ;
 RECT 30.605 0.26 30.735 0.39 ;
 RECT 12.53 1.52 12.66 1.65 ;
 RECT 27.845 1.075 27.975 1.205 ;
 RECT 15.56 0.925 15.69 1.055 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 2.58 1.6 2.71 1.73 ;
 RECT 3.655 2.01 3.785 2.14 ;
 RECT 3.655 0.735 3.785 0.865 ;
 RECT 2.415 2.075 2.545 2.205 ;
 RECT 1.275 2.275 1.405 2.405 ;
 RECT 3.185 0.545 3.315 0.675 ;
 RECT 3.655 1.75 3.785 1.88 ;
 RECT 0.805 2.015 0.935 2.145 ;
 RECT 2.22 0.735 2.35 0.865 ;
 RECT 2.4 1.19 2.53 1.32 ;
 RECT 30.95 1.49 31.08 1.62 ;
 RECT 6.23 0.88 6.36 1.01 ;
 RECT 15.47 1.87 15.6 2 ;
 RECT 9.375 2.025 9.505 2.155 ;
 RECT 8.025 0.32 8.155 0.45 ;
 RECT 28.72 0.135 28.85 0.265 ;
 RECT 5.24 1.495 5.37 1.625 ;
 RECT 5.145 0.745 5.275 0.875 ;
 RECT 5.03 1.995 5.16 2.125 ;
 RECT 12.64 1.995 12.77 2.125 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 12.195 2.07 12.325 2.2 ;
 RECT 14.965 0.595 15.095 0.725 ;
 RECT 13.705 1.24 13.835 1.37 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 23.96 1.725 24.09 1.855 ;
 RECT 24.52 0.62 24.65 0.75 ;
 RECT 23.96 0.62 24.09 0.75 ;
 RECT 25.02 1.71 25.15 1.84 ;
 RECT 24.435 2.64 24.565 2.77 ;
 RECT 25.02 0.63 25.15 0.76 ;
 RECT 21.69 2.64 21.82 2.77 ;
 RECT 10.4 2.045 10.53 2.175 ;
 RECT 10.67 1.23 10.8 1.36 ;
 RECT 19.49 1.705 19.62 1.835 ;
 RECT 9.86 2.075 9.99 2.205 ;
 RECT 6.7 0.88 6.83 1.01 ;
 RECT 17.52 1.835 17.65 1.965 ;
 RECT 17.39 0.765 17.52 0.895 ;
 RECT 4.52 0.74 4.65 0.87 ;
 RECT 31.115 0.12 31.245 0.25 ;
 RECT 7.415 0.53 7.545 0.66 ;
 RECT 16.365 2.38 16.495 2.51 ;
 RECT 12.64 0.905 12.77 1.035 ;
 RECT 28.25 1.425 28.38 1.555 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 20.555 0.92 20.685 1.05 ;
 RECT 28.72 1.475 28.85 1.605 ;
 RECT 14.44 0.875 14.57 1.005 ;
 RECT 5.855 0.79 5.985 0.92 ;
 RECT 18.46 1.835 18.59 1.965 ;
 RECT 6.79 2.07 6.92 2.2 ;
 RECT 32.675 1.475 32.805 1.605 ;
 RECT 23.285 1.705 23.415 1.835 ;
 RECT 26.075 1.71 26.205 1.84 ;
 RECT 4.025 0.74 4.155 0.87 ;
 RECT 5.86 1.825 5.99 1.955 ;
 RECT 14.44 1.945 14.57 2.075 ;
 RECT 4.495 2.05 4.625 2.18 ;
 RECT 28 0.505 28.13 0.635 ;
 RECT 11.715 2.015 11.845 2.145 ;
 RECT 29.935 0.12 30.065 0.25 ;
 RECT 29.5 1.485 29.63 1.615 ;
 RECT 31.895 1.465 32.025 1.595 ;
 RECT 19.96 1.705 20.09 1.835 ;
 RECT 31.895 0.595 32.025 0.725 ;
 RECT 13.34 2.225 13.47 2.355 ;
 RECT 23.285 0.975 23.415 1.105 ;
 RECT 25.49 2.64 25.62 2.77 ;
 RECT 4.025 2.115 4.155 2.245 ;
 RECT 22.77 0.36 22.9 0.49 ;
 RECT 26.075 0.63 26.205 0.76 ;
 RECT 30.44 0.595 30.57 0.725 ;
 RECT 7.74 1.675 7.87 1.805 ;
 RECT 20.435 1.705 20.565 1.835 ;
 RECT 22.685 2.64 22.815 2.77 ;
 RECT 30.58 1.405 30.71 1.535 ;
 RECT 11.72 0.905 11.85 1.035 ;
 RECT 4.19 0.325 4.32 0.455 ;
 RECT 9.86 0.315 9.99 0.445 ;
 RECT 12.195 0.905 12.325 1.035 ;
 RECT 15.47 0.595 15.6 0.725 ;
 RECT 13.53 0.595 13.66 0.725 ;
 RECT 30.105 1.445 30.235 1.575 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 18.495 1.035 18.625 1.165 ;
 RECT 19.08 0.91 19.21 1.04 ;
 RECT 10.89 2.405 11.02 2.535 ;
 RECT 25.575 0.62 25.705 0.75 ;
 RECT 6.29 2.105 6.42 2.235 ;
 RECT 7.26 2.025 7.39 2.155 ;
 RECT 5.215 0.145 5.345 0.275 ;
 RECT 14.965 1.9 15.095 2.03 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 5.23 2.345 5.36 2.475 ;
 RECT 29.5 0.435 29.63 0.565 ;
 RECT 8.83 2.305 8.96 2.435 ;
 RECT 8.77 0.565 8.9 0.695 ;
 RECT 24.285 1.29 24.415 1.42 ;
 RECT 6.615 0.525 6.745 0.655 ;
 RECT 5.965 1.49 6.095 1.62 ;
 RECT 8.07 2.305 8.2 2.435 ;
 RECT 7.05 1.265 7.18 1.395 ;
 RECT 2.855 0.26 2.985 0.39 ;
 RECT 3.32 1.155 3.45 1.285 ;
 RECT 20.845 1.285 20.975 1.415 ;
 RECT 18.665 0.43 18.795 0.56 ;
 RECT 20.285 0.6 20.415 0.73 ;
 RECT 20.83 0.26 20.96 0.39 ;
 RECT 19.305 2.075 19.435 2.205 ;
 RECT 10.735 1.66 10.865 1.79 ;
 RECT 10.02 1.585 10.15 1.715 ;
 RECT 26.805 0.26 26.935 0.39 ;
 RECT 31.745 1.03 31.875 1.16 ;
 RECT 16.965 0.495 17.095 0.625 ;
 RECT 18.155 1.43 18.285 1.56 ;
 RECT 16.24 0.625 16.37 0.755 ;
 RECT 16.16 1.445 16.29 1.575 ;
 RECT 28.895 1.075 29.025 1.205 ;
 RECT 11.29 0.935 11.42 1.065 ;
 RECT 29.82 0.975 29.95 1.105 ;
 RECT 17.82 0.665 17.95 0.795 ;
 RECT 29.34 1.035 29.47 1.165 ;
 RECT 31.78 2.31 31.91 2.44 ;
 RECT 14.535 2.34 14.665 2.47 ;
 RECT 27.585 0.635 27.715 0.765 ;
 RECT 4.675 1.55 4.805 1.68 ;
 RECT 21.285 1.705 21.415 1.835 ;
 RECT 22.29 1.705 22.42 1.835 ;
 RECT 21.285 0.975 21.415 1.105 ;
 RECT 22.29 0.975 22.42 1.105 ;
 RECT 21.775 0.36 21.905 0.49 ;
 RECT 1.275 0.735 1.405 0.865 ;
 RECT 1.28 1.51 1.41 1.64 ;
 RECT 0.805 0.735 0.935 0.865 ;
 RECT 3.185 2.31 3.315 2.44 ;
 RECT 1.275 2.015 1.405 2.145 ;
 RECT 1.88 1.155 2.01 1.285 ;
 LAYER M1 ;
 RECT 29.495 1.345 29.955 1.485 ;
 RECT 29.77 0.935 30 1.145 ;
 RECT 29.495 0.59 29.955 0.73 ;
 RECT 30.435 0.73 30.575 1.04 ;
 RECT 30.575 1.18 30.715 1.605 ;
 RECT 30.37 0.59 30.645 0.73 ;
 RECT 31.695 0.99 31.925 1.04 ;
 RECT 30.435 1.04 31.925 1.18 ;
 RECT 31.695 1.18 31.925 1.2 ;
 RECT 30.555 0.29 30.925 0.43 ;
 RECT 30.785 0.43 30.925 0.71 ;
 RECT 30.555 0.22 30.785 0.29 ;
 RECT 32.205 0.85 32.345 1.385 ;
 RECT 31.89 1.525 32.03 1.73 ;
 RECT 30.785 0.71 32.345 0.85 ;
 RECT 31.89 0.51 32.03 0.71 ;
 RECT 31.89 1.385 32.345 1.525 ;
 RECT 27.795 1.225 28.025 1.245 ;
 RECT 27.795 1.195 28.385 1.225 ;
 RECT 27.935 1.015 28.245 1.035 ;
 RECT 27.795 1.035 28.245 1.055 ;
 RECT 28.07 0.64 28.21 1.015 ;
 RECT 28.245 1.225 28.385 1.75 ;
 RECT 27.95 0.5 28.21 0.64 ;
 RECT 28.845 1.035 29.075 1.055 ;
 RECT 28.845 1.195 29.075 1.245 ;
 RECT 27.795 1.055 29.075 1.195 ;
 RECT 26.755 0.36 26.985 0.43 ;
 RECT 28.35 0.36 28.49 0.565 ;
 RECT 26.755 0.22 28.49 0.36 ;
 RECT 29.09 0.705 29.23 0.75 ;
 RECT 29.215 0.995 29.52 1.205 ;
 RECT 29.215 0.89 29.355 0.995 ;
 RECT 29.09 0.75 29.355 0.89 ;
 RECT 28.35 0.565 29.23 0.705 ;
 RECT 15.465 0.525 15.605 0.885 ;
 RECT 15.465 1.095 15.605 2.065 ;
 RECT 15.465 0.885 15.74 1.095 ;
 RECT 12.19 1.04 12.33 2.34 ;
 RECT 12.19 0.895 12.33 0.9 ;
 RECT 12.12 0.9 12.395 1.04 ;
 RECT 12.985 2.055 13.125 2.34 ;
 RECT 12.19 2.34 13.125 2.48 ;
 RECT 14.12 1.66 14.26 1.915 ;
 RECT 12.985 1.915 14.26 2.055 ;
 RECT 14.435 0.765 14.575 1.52 ;
 RECT 14.435 1.66 14.575 2.145 ;
 RECT 14.96 0.525 15.1 1.52 ;
 RECT 14.96 1.66 15.1 2.11 ;
 RECT 14.12 1.52 15.1 1.66 ;
 RECT 19.51 0.775 19.65 1.405 ;
 RECT 20.235 0.56 20.465 0.635 ;
 RECT 18.49 1.405 19.65 1.545 ;
 RECT 18.49 1.545 18.63 1.83 ;
 RECT 17.445 1.83 18.695 1.97 ;
 RECT 18.49 1.17 18.63 1.405 ;
 RECT 18.42 1.03 18.7 1.17 ;
 RECT 23.535 0.36 23.675 0.635 ;
 RECT 19.51 0.635 23.675 0.775 ;
 RECT 24.235 0.36 24.375 1.25 ;
 RECT 24.235 1.25 24.465 1.46 ;
 RECT 23.535 0.22 24.375 0.36 ;
 RECT 20.78 0.22 21.01 0.28 ;
 RECT 20.78 0.42 21.01 0.43 ;
 RECT 18.615 0.28 21.01 0.42 ;
 RECT 18.615 0.42 18.845 0.6 ;
 RECT 16.19 0.585 17.145 0.63 ;
 RECT 16.915 0.63 17.145 0.665 ;
 RECT 16.915 0.455 17.145 0.49 ;
 RECT 16.215 0.49 17.145 0.585 ;
 RECT 16.19 0.63 16.42 0.795 ;
 RECT 17.77 0.57 18 0.95 ;
 RECT 8.72 0.525 8.95 0.605 ;
 RECT 7.365 0.485 7.68 0.605 ;
 RECT 17.76 1.23 17.9 1.42 ;
 RECT 15.91 1.09 17.9 1.23 ;
 RECT 15.91 0.385 16.05 1.09 ;
 RECT 13.9 0.385 14.04 0.875 ;
 RECT 13.9 0.255 16.05 0.385 ;
 RECT 13.9 0.245 16.045 0.255 ;
 RECT 12.985 0.875 14.04 1.015 ;
 RECT 12.985 0.745 13.125 0.875 ;
 RECT 7.365 0.605 13.125 0.745 ;
 RECT 18.105 1.39 18.335 1.42 ;
 RECT 17.76 1.42 18.335 1.56 ;
 RECT 18.105 1.56 18.335 1.6 ;
 RECT 7.085 0.895 11.47 1.035 ;
 RECT 11.24 1.035 11.47 1.105 ;
 RECT 7.085 0.66 7.225 0.895 ;
 RECT 6.565 0.485 6.795 0.52 ;
 RECT 6.565 0.66 6.795 0.695 ;
 RECT 6.565 0.52 7.225 0.66 ;
 RECT 3.935 0.875 4.075 1.195 ;
 RECT 3.935 1.335 4.075 2.11 ;
 RECT 3.935 0.735 4.225 0.875 ;
 RECT 3.935 2.11 4.225 2.25 ;
 RECT 4.795 0.575 4.935 1.195 ;
 RECT 3.935 1.195 4.935 1.335 ;
 RECT 6.285 0.36 6.425 0.875 ;
 RECT 6.285 1.015 6.425 2.305 ;
 RECT 5.65 0.36 5.79 0.435 ;
 RECT 6.175 0.875 6.49 1.015 ;
 RECT 5.65 0.22 6.425 0.36 ;
 RECT 4.795 0.435 5.79 0.575 ;
 RECT 3.65 0.46 3.79 2.21 ;
 RECT 4.05 0.22 4.375 0.32 ;
 RECT 4.05 0.46 4.375 0.525 ;
 RECT 3.65 0.32 4.375 0.46 ;
 RECT 0.8 0.68 0.94 1.155 ;
 RECT 0.8 1.295 0.94 2.23 ;
 RECT 1.585 0.36 1.725 1.155 ;
 RECT 0.8 1.155 1.725 1.295 ;
 RECT 2.805 0.36 3.035 0.43 ;
 RECT 1.585 0.22 3.035 0.36 ;
 RECT 16.88 1.895 17.02 2.39 ;
 RECT 20.805 2.205 20.945 2.39 ;
 RECT 16.88 2.39 20.945 2.53 ;
 RECT 15.755 1.755 17.02 1.895 ;
 RECT 15.755 1.895 15.895 2.34 ;
 RECT 14.485 2.3 14.715 2.34 ;
 RECT 14.485 2.48 14.715 2.51 ;
 RECT 14.485 2.34 15.895 2.48 ;
 RECT 20.805 2.065 27.53 2.205 ;
 RECT 27.39 2.205 27.53 2.52 ;
 RECT 31.73 2.48 31.87 2.52 ;
 RECT 27.39 2.52 31.87 2.66 ;
 RECT 31.73 2.27 31.96 2.48 ;
 RECT 20.515 1.055 20.655 1.245 ;
 RECT 19.955 1.385 20.095 1.625 ;
 RECT 20.795 1.385 21.025 1.455 ;
 RECT 19.955 1.245 21.025 1.385 ;
 RECT 20.485 0.915 20.785 1.055 ;
 RECT 19.925 1.625 20.18 1.92 ;
 RECT 20.32 1.7 20.615 1.84 ;
 RECT 20.32 1.84 20.46 2.075 ;
 RECT 19.625 1.84 19.765 2.075 ;
 RECT 19.43 1.7 19.765 1.84 ;
 RECT 19.625 2.075 20.46 2.215 ;
 RECT 17.16 1.56 17.3 2.11 ;
 RECT 17.16 2.11 19.485 2.245 ;
 RECT 17.16 2.245 19.48 2.25 ;
 RECT 19.255 2.035 19.485 2.11 ;
 RECT 16.11 1.405 16.34 1.42 ;
 RECT 16.11 1.56 16.34 1.615 ;
 RECT 16.11 1.42 17.3 1.56 ;
 RECT 12.635 1.04 12.775 1.48 ;
 RECT 12.48 1.48 12.775 1.635 ;
 RECT 12.635 1.775 12.775 2.18 ;
 RECT 12.565 0.9 12.84 1.04 ;
 RECT 13.675 1.375 13.815 1.635 ;
 RECT 12.635 1.69 13.82 1.775 ;
 RECT 12.48 1.635 13.82 1.69 ;
 RECT 13.635 1.235 13.905 1.375 ;
 RECT 5.14 1.69 5.28 1.99 ;
 RECT 5.14 0.93 5.28 1.44 ;
 RECT 4.96 1.99 5.28 2.13 ;
 RECT 5.075 0.715 5.325 0.93 ;
 RECT 5.14 1.44 5.47 1.69 ;
 RECT 7.19 2.125 7.465 2.205 ;
 RECT 9.3 2.125 9.575 2.205 ;
 RECT 7.19 1.985 9.575 2.125 ;
 RECT 6.63 1.84 6.77 2.015 ;
 RECT 7.67 1.685 7.945 1.7 ;
 RECT 6.63 1.015 6.77 1.7 ;
 RECT 6.63 1.7 7.945 1.84 ;
 RECT 6.63 0.875 6.945 1.015 ;
 RECT 6.63 2.015 6.995 2.215 ;
 RECT 9.97 1.685 10.2 1.755 ;
 RECT 7.67 1.545 10.2 1.685 ;
 RECT 5.875 1.67 6.015 1.82 ;
 RECT 5.875 1.96 6.015 2.52 ;
 RECT 5.875 0.96 6.015 1.44 ;
 RECT 8.02 2.265 8.25 2.52 ;
 RECT 5.81 1.82 6.08 1.96 ;
 RECT 5.875 1.44 6.145 1.67 ;
 RECT 5.78 0.75 6.035 0.96 ;
 RECT 5.875 2.52 8.25 2.66 ;
 RECT 7 1.365 7.23 1.435 ;
 RECT 10.395 1.365 10.535 2.25 ;
 RECT 11.71 1.04 11.85 1.25 ;
 RECT 11.71 1.39 11.85 2.215 ;
 RECT 11.71 0.885 11.85 0.9 ;
 RECT 7 1.25 11.85 1.365 ;
 RECT 7 1.225 11.1 1.25 ;
 RECT 10.96 1.365 11.85 1.39 ;
 RECT 11.645 0.9 11.92 1.04 ;
 RECT 2.87 0.87 3.01 1.15 ;
 RECT 2.87 1.29 3.01 2.07 ;
 RECT 2.165 0.73 3.01 0.87 ;
 RECT 2.36 2.07 3.01 2.21 ;
 RECT 2.87 1.15 3.5 1.29 ;
 RECT 3.27 1.115 3.5 1.15 ;
 RECT 3.27 1.29 3.5 1.325 ;
 RECT 29.815 1.145 29.955 1.345 ;
 RECT 29.495 1.485 29.635 1.76 ;
 RECT 29.815 0.73 29.955 0.935 ;
 RECT 29.495 0.355 29.635 0.59 ;
 END
END RSDFFSRASX2

MACRO RSDFFSRSSRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 30.08 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 30.08 0.08 ;
 RECT 26.88 0.08 27.12 0.26 ;
 RECT 20.165 0.335 20.47 0.475 ;
 RECT 3.15 0.08 3.29 0.685 ;
 RECT 6.595 0.08 6.735 1.055 ;
 RECT 4.115 0.08 4.255 0.565 ;
 RECT 7.34 0.08 7.48 0.39 ;
 RECT 9.94 0.08 10.175 0.515 ;
 RECT 12.815 0.08 12.955 0.815 ;
 RECT 16.375 0.08 16.515 0.5 ;
 RECT 18.18 0.08 18.32 0.525 ;
 RECT 24.53 0.08 24.67 0.36 ;
 RECT 21.945 0.08 22.085 0.82 ;
 RECT 25.745 0.08 25.885 0.35 ;
 RECT 0.65 0.08 0.92 0.245 ;
 RECT 20.25 0.08 20.39 0.335 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 30.08 2.96 ;
 RECT 2.83 1.87 2.97 2.8 ;
 RECT 9.33 2.29 9.59 2.545 ;
 RECT 0.925 1.89 1.065 2.8 ;
 RECT 7.27 2.59 7.52 2.8 ;
 RECT 6.53 2.59 6.78 2.8 ;
 RECT 4.115 2.365 4.255 2.8 ;
 RECT 10.525 2.07 10.665 2.8 ;
 RECT 12.625 2.375 12.765 2.8 ;
 RECT 16.85 2.57 16.99 2.8 ;
 RECT 20.27 2.57 20.41 2.8 ;
 RECT 18.175 2.57 18.315 2.8 ;
 RECT 21.86 2.57 22 2.8 ;
 RECT 9.405 2.545 9.545 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.6 1.475 6.975 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 21.32 1.765 22.585 1.905 ;
 RECT 21.385 0.55 21.525 1.71 ;
 RECT 21.32 1.905 21.585 2.04 ;
 RECT 21.32 1.71 21.585 1.765 ;
 RECT 22.445 1.905 22.585 1.93 ;
 RECT 22.445 1.64 22.585 1.765 ;
 END
 ANTENNADIFFAREA 0.59 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.68 1.165 20.92 1.465 ;
 RECT 20.72 0.915 20.86 1.165 ;
 RECT 19.78 1.765 20.86 1.905 ;
 RECT 20.72 1.465 20.86 1.765 ;
 RECT 19.78 0.905 19.92 1.765 ;
 END
 ANTENNADIFFAREA 0.59 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13 2.12 13.265 2.475 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 28.44 1.435 28.78 1.8 ;
 RECT 26.76 1.99 28.625 2.13 ;
 RECT 24.53 2.22 26.9 2.36 ;
 RECT 26.76 1.435 26.9 1.99 ;
 RECT 28.485 1.8 28.625 1.99 ;
 RECT 24.53 1.39 24.67 2.22 ;
 RECT 25.915 1.37 26.055 2.22 ;
 RECT 26.76 2.13 26.9 2.22 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 23.21 0.59 23.58 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.035 1.365 4.455 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.96 2.12 6.2 2.395 ;
 RECT 5.405 2.395 6.2 2.535 ;
 RECT 5.405 2.535 5.635 2.57 ;
 RECT 5.405 2.36 5.635 2.395 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.905 0.825 3.27 1.08 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END RSTB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.155 1.45 1.7 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.52 1.15 0.96 1.4 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SETB

 OBS
 LAYER PO ;
 RECT 11.265 1.13 12.28 1.23 ;
 RECT 13.025 2.255 13.255 2.465 ;
 RECT 15.715 0.685 15.945 0.875 ;
 RECT 15.045 0.82 15.275 0.875 ;
 RECT 15.045 0.975 15.275 1.03 ;
 RECT 15.045 0.875 15.95 0.975 ;
 RECT 18.43 1.635 18.53 1.66 ;
 RECT 18.43 1.66 18.685 1.87 ;
 RECT 18.43 1.87 18.53 2.565 ;
 RECT 19.09 0.19 19.19 0.22 ;
 RECT 20.035 0.19 20.135 1.435 ;
 RECT 20.035 1.535 20.135 2.37 ;
 RECT 20.505 0.5 20.605 1.435 ;
 RECT 20.505 1.535 20.605 2.37 ;
 RECT 19.09 0.09 20.135 0.19 ;
 RECT 20.03 1.435 20.605 1.535 ;
 RECT 18.96 0.22 19.19 0.43 ;
 RECT 18.705 1.25 18.965 1.3 ;
 RECT 18.865 0.61 18.965 1.25 ;
 RECT 18.705 1.4 18.965 1.46 ;
 RECT 18.865 1.46 18.965 2.56 ;
 RECT 19.395 0.68 19.495 1.3 ;
 RECT 18.705 1.3 19.495 1.4 ;
 RECT 19.38 0.47 19.61 0.68 ;
 RECT 17.105 0.51 17.205 0.53 ;
 RECT 17.105 0.74 17.205 2.21 ;
 RECT 17.065 0.53 17.295 0.74 ;
 RECT 16.635 0.54 16.885 0.695 ;
 RECT 16.635 0.695 16.735 2.21 ;
 RECT 16.655 0.485 16.885 0.54 ;
 RECT 13.47 2.69 15.38 2.695 ;
 RECT 15.28 2.54 15.38 2.69 ;
 RECT 14.26 2.695 15.38 2.79 ;
 RECT 13.47 0.66 13.57 2.595 ;
 RECT 13.47 2.595 14.36 2.69 ;
 RECT 15.28 2.33 15.51 2.54 ;
 RECT 14.505 1.355 15.6 1.39 ;
 RECT 14.505 0.19 14.605 1.29 ;
 RECT 14.505 1.29 15.595 1.355 ;
 RECT 8.015 0.19 8.115 0.51 ;
 RECT 9.75 0.19 9.85 1.24 ;
 RECT 15.37 1.39 15.6 1.565 ;
 RECT 7.975 0.51 8.22 0.755 ;
 RECT 8.015 0.09 14.605 0.19 ;
 RECT 15.075 1.71 15.175 1.76 ;
 RECT 10.8 0.48 10.985 0.5 ;
 RECT 18.435 0.19 18.535 1.18 ;
 RECT 16.135 0.19 16.235 1.76 ;
 RECT 15.075 1.76 16.235 1.86 ;
 RECT 13.99 0.48 14.09 1.61 ;
 RECT 14.54 1.71 14.64 2.445 ;
 RECT 16.135 0.09 18.535 0.19 ;
 RECT 13.99 1.61 15.175 1.71 ;
 RECT 10.8 0.38 14.09 0.48 ;
 RECT 10.755 0.5 10.985 0.71 ;
 RECT 11.255 1.575 11.355 2.485 ;
 RECT 11.765 1.41 11.995 1.475 ;
 RECT 11.765 1.575 11.995 1.62 ;
 RECT 11.255 1.475 11.995 1.575 ;
 RECT 3.515 2.15 3.615 2.69 ;
 RECT 3.515 2.69 5.03 2.79 ;
 RECT 4.93 1.495 5.03 2.69 ;
 RECT 3.385 1.88 3.615 2.15 ;
 RECT 1.65 0.66 1.75 1.45 ;
 RECT 1.46 1.45 1.75 1.685 ;
 RECT 1.65 1.685 1.75 2.38 ;
 RECT 1.18 1.69 1.28 2.59 ;
 RECT 0.265 2.29 0.495 2.59 ;
 RECT 0.265 2.59 1.28 2.69 ;
 RECT 4.46 0.555 4.56 1.365 ;
 RECT 4.46 1.6 4.56 2.185 ;
 RECT 4.18 1.365 4.56 1.6 ;
 RECT 2.815 0.48 2.915 0.835 ;
 RECT 1.18 0.48 1.28 1.24 ;
 RECT 2.815 1.07 2.915 1.625 ;
 RECT 2.12 1.725 2.22 2.73 ;
 RECT 2.815 0.835 3.22 1.07 ;
 RECT 1.18 0.38 2.915 0.48 ;
 RECT 2.12 1.625 2.915 1.725 ;
 RECT 0.71 0.48 0.81 1.155 ;
 RECT 0.71 1.155 0.95 1.39 ;
 RECT 0.71 1.39 0.81 2.38 ;
 RECT 5.325 0.16 5.59 0.465 ;
 RECT 5.49 0.465 5.59 1.13 ;
 RECT 10.615 1.61 10.88 1.82 ;
 RECT 10.78 1.82 10.88 2.49 ;
 RECT 10.41 0.66 10.51 1.51 ;
 RECT 10.41 1.51 10.88 1.61 ;
 RECT 13.075 0.66 13.175 1.24 ;
 RECT 12.945 1.24 13.175 1.475 ;
 RECT 6.855 0.655 6.955 1.495 ;
 RECT 6.66 1.495 6.955 1.745 ;
 RECT 6.855 1.745 6.955 2.19 ;
 RECT 6.14 0.27 6.48 0.52 ;
 RECT 6.38 0.52 6.48 2.31 ;
 RECT 8.515 1.595 8.615 2.33 ;
 RECT 7.975 1.445 8.22 1.495 ;
 RECT 7.975 1.495 8.615 1.595 ;
 RECT 7.975 1.595 8.22 1.69 ;
 RECT 7.695 1.265 7.795 1.52 ;
 RECT 7.195 1.52 7.795 1.62 ;
 RECT 7.63 1.62 7.73 2.69 ;
 RECT 10.31 1.79 10.41 2.69 ;
 RECT 8.56 0.375 8.845 0.61 ;
 RECT 8.56 0.61 8.66 1.165 ;
 RECT 7.195 1.44 7.44 1.52 ;
 RECT 7.195 1.62 7.44 1.69 ;
 RECT 7.695 0.585 7.795 1.165 ;
 RECT 7.63 2.69 10.41 2.79 ;
 RECT 7.695 1.165 8.66 1.265 ;
 RECT 5.4 1.41 5.5 2.36 ;
 RECT 5.21 1.31 5.5 1.41 ;
 RECT 4.93 0.23 5.03 1.21 ;
 RECT 3.9 0.23 4 2.185 ;
 RECT 4.93 1.21 5.31 1.31 ;
 RECT 5.4 2.36 5.635 2.57 ;
 RECT 3.9 0.13 5.03 0.23 ;
 RECT 9.05 0.65 9.15 1.23 ;
 RECT 9.01 1.44 9.11 2.33 ;
 RECT 9 1.23 9.23 1.44 ;
 RECT 2.12 0.66 2.22 1.195 ;
 RECT 2.385 1.43 2.615 1.435 ;
 RECT 2.12 1.195 2.63 1.43 ;
 RECT 9.45 0.6 9.55 1.61 ;
 RECT 9.485 1.71 9.585 2.285 ;
 RECT 9.33 0.37 9.57 0.6 ;
 RECT 9.45 1.61 9.585 1.71 ;
 RECT 9.36 2.285 9.59 2.5 ;
 RECT 24.79 1.245 24.89 2.02 ;
 RECT 24.66 1.035 24.89 1.245 ;
 RECT 21.645 0.385 21.745 1.2 ;
 RECT 22.225 0.375 22.325 1.33 ;
 RECT 21.63 1.2 21.84 1.33 ;
 RECT 21.63 1.43 21.84 1.435 ;
 RECT 21.63 1.33 22.325 1.43 ;
 RECT 21.645 1.435 21.745 2.555 ;
 RECT 22.225 1.43 22.325 2.565 ;
 RECT 22.77 0.22 23 0.275 ;
 RECT 22.77 0.375 23 0.43 ;
 RECT 22.225 0.275 23 0.375 ;
 RECT 26.005 0.38 26.105 0.96 ;
 RECT 26.005 1.06 26.105 1.14 ;
 RECT 25.585 0.935 25.815 0.96 ;
 RECT 25.585 0.96 26.105 1.06 ;
 RECT 25.585 1.06 25.815 1.145 ;
 RECT 26.005 1.14 26.275 1.24 ;
 RECT 26.175 1.24 26.275 1.84 ;
 RECT 26.37 0.22 26.6 0.28 ;
 RECT 26.37 0.38 26.6 0.43 ;
 RECT 26.005 0.28 26.6 0.38 ;
 RECT 28.19 0.195 28.29 2.665 ;
 RECT 27.18 0.095 28.29 0.195 ;
 RECT 23.555 1.245 23.655 2.665 ;
 RECT 23.555 1.2 23.84 1.245 ;
 RECT 27.18 0.195 27.28 0.945 ;
 RECT 23.61 1.035 23.84 1.1 ;
 RECT 23.555 2.665 28.29 2.765 ;
 RECT 23.555 1.1 23.885 1.2 ;
 RECT 25.095 0.215 25.195 0.995 ;
 RECT 25.095 0.995 25.335 1.205 ;
 RECT 25.095 1.205 25.195 2 ;
 RECT 27.49 0.375 27.59 0.99 ;
 RECT 27.49 0.99 27.74 1.2 ;
 RECT 27.49 1.2 27.59 2.27 ;
 RECT 27.49 2.27 27.775 2.48 ;
 RECT 24.315 0.855 24.415 2.2 ;
 RECT 27.18 1.125 27.28 2.2 ;
 RECT 23.35 0.755 24.885 0.84 ;
 RECT 23.35 0.84 24.88 0.855 ;
 RECT 24.785 0.215 24.885 0.755 ;
 RECT 24.315 0.21 24.415 0.755 ;
 RECT 23.35 0.595 23.58 0.755 ;
 RECT 24.315 2.2 27.28 2.3 ;
 RECT 12.18 0.66 12.28 1.13 ;
 RECT 12.18 1.23 12.28 1.655 ;
 RECT 11.265 0.66 11.365 1.13 ;
 RECT 12.18 1.655 13.14 1.755 ;
 RECT 13.04 1.755 13.14 2.255 ;
 RECT 12.18 1.755 12.28 2.57 ;
 LAYER CO ;
 RECT 18.755 1.29 18.885 1.42 ;
 RECT 17.115 0.57 17.245 0.7 ;
 RECT 16.705 0.525 16.835 0.655 ;
 RECT 15.33 2.37 15.46 2.5 ;
 RECT 15.42 1.395 15.55 1.525 ;
 RECT 10.805 0.54 10.935 0.67 ;
 RECT 11.815 1.45 11.945 1.58 ;
 RECT 17.325 0.975 17.455 1.105 ;
 RECT 17.325 1.705 17.455 1.835 ;
 RECT 16.855 2.64 16.985 2.77 ;
 RECT 16.385 1.7 16.515 1.83 ;
 RECT 12.63 2.445 12.76 2.575 ;
 RECT 2.835 2.255 2.965 2.385 ;
 RECT 4.265 1.42 4.395 1.55 ;
 RECT 5.62 1.8 5.75 1.93 ;
 RECT 1.4 1.965 1.53 2.095 ;
 RECT 5.71 0.85 5.84 0.98 ;
 RECT 0.72 0.11 0.85 0.24 ;
 RECT 5.15 0.78 5.28 0.91 ;
 RECT 1.87 1.965 2 2.095 ;
 RECT 0.93 1.965 1.06 2.095 ;
 RECT 4.12 2.435 4.25 2.565 ;
 RECT 3.56 1.49 3.69 1.62 ;
 RECT 1.51 1.505 1.64 1.635 ;
 RECT 4.68 0.78 4.81 0.91 ;
 RECT 4.12 0.35 4.25 0.48 ;
 RECT 3.445 1.94 3.575 2.07 ;
 RECT 4.68 1.725 4.81 1.855 ;
 RECT 26.395 1.405 26.525 1.535 ;
 RECT 23.815 0.505 23.945 0.635 ;
 RECT 25.315 1.485 25.445 1.615 ;
 RECT 25.75 0.12 25.88 0.25 ;
 RECT 26.765 1.49 26.895 1.62 ;
 RECT 24.535 1.475 24.665 1.605 ;
 RECT 25.92 1.445 26.05 1.575 ;
 RECT 26.93 0.12 27.06 0.25 ;
 RECT 27.71 1.465 27.84 1.595 ;
 RECT 24.535 0.135 24.665 0.265 ;
 RECT 28.49 1.475 28.62 1.605 ;
 RECT 25.315 0.435 25.445 0.565 ;
 RECT 27.71 0.595 27.84 0.725 ;
 RECT 24.065 1.425 24.195 1.555 ;
 RECT 26.255 0.595 26.385 0.725 ;
 RECT 20.255 0.34 20.385 0.47 ;
 RECT 20.275 2.64 20.405 2.77 ;
 RECT 20.725 1.705 20.855 1.835 ;
 RECT 20.725 0.975 20.855 1.105 ;
 RECT 19.785 0.975 19.915 1.105 ;
 RECT 14.76 0.595 14.89 0.725 ;
 RECT 14.76 1.87 14.89 2 ;
 RECT 14.255 0.595 14.385 0.725 ;
 RECT 14.255 1.9 14.385 2.03 ;
 RECT 19.785 1.705 19.915 1.835 ;
 RECT 21.39 0.625 21.52 0.755 ;
 RECT 22.45 1.71 22.58 1.84 ;
 RECT 21.865 2.64 21.995 2.77 ;
 RECT 21.39 1.725 21.52 1.855 ;
 RECT 21.67 1.25 21.8 1.38 ;
 RECT 21.95 0.62 22.08 0.75 ;
 RECT 6.6 2.64 6.73 2.77 ;
 RECT 3.04 0.89 3.17 1.02 ;
 RECT 0.77 1.21 0.9 1.34 ;
 RECT 3.645 0.78 3.775 0.91 ;
 RECT 2.34 1.965 2.47 2.095 ;
 RECT 2.835 1.995 2.965 2.125 ;
 RECT 0.46 0.705 0.59 0.835 ;
 RECT 1.87 0.885 2 1.015 ;
 RECT 1.4 0.885 1.53 1.015 ;
 RECT 0.315 2.345 0.445 2.475 ;
 RECT 3.155 0.5 3.285 0.63 ;
 RECT 5.375 0.26 5.505 0.39 ;
 RECT 2.34 0.885 2.47 1.015 ;
 RECT 3.155 0.24 3.285 0.37 ;
 RECT 5.15 1.725 5.28 1.855 ;
 RECT 0.46 1.965 0.59 2.095 ;
 RECT 19.085 0.83 19.215 0.96 ;
 RECT 18.185 0.33 18.315 0.46 ;
 RECT 19.085 1.78 19.215 1.91 ;
 RECT 18.18 2.64 18.31 2.77 ;
 RECT 7.85 1.825 7.98 1.955 ;
 RECT 12.995 1.28 13.125 1.41 ;
 RECT 11 2.015 11.13 2.145 ;
 RECT 11.93 0.88 12.06 1.01 ;
 RECT 13.73 1.945 13.86 2.075 ;
 RECT 12.82 0.62 12.95 0.75 ;
 RECT 9.385 0.42 9.515 0.55 ;
 RECT 8.76 1.925 8.89 2.055 ;
 RECT 6.6 0.875 6.73 1.005 ;
 RECT 9.99 0.325 10.12 0.455 ;
 RECT 8.03 1.49 8.16 1.62 ;
 RECT 8.03 0.555 8.16 0.685 ;
 RECT 8.78 0.88 8.91 1.01 ;
 RECT 6.2 0.325 6.33 0.455 ;
 RECT 6.13 0.875 6.26 1.005 ;
 RECT 10.53 2.135 10.66 2.265 ;
 RECT 7.34 2.64 7.47 2.77 ;
 RECT 11.485 2.07 11.615 2.2 ;
 RECT 6.125 1.675 6.255 1.805 ;
 RECT 9.23 1.98 9.36 2.11 ;
 RECT 7.915 0.905 8.045 1.035 ;
 RECT 8.265 1.96 8.395 2.09 ;
 RECT 7.205 0.875 7.335 1.005 ;
 RECT 9.705 1.675 9.835 1.805 ;
 RECT 6.72 1.55 6.85 1.68 ;
 RECT 7.345 0.21 7.475 0.34 ;
 RECT 10.06 2.125 10.19 2.255 ;
 RECT 7.075 1.92 7.205 2.05 ;
 RECT 8.31 0.88 8.44 1.01 ;
 RECT 11 0.93 11.13 1.06 ;
 RECT 8.665 0.43 8.795 0.56 ;
 RECT 11.93 1.995 12.06 2.125 ;
 RECT 11.485 0.88 11.615 1.01 ;
 RECT 7.255 1.495 7.385 1.625 ;
 RECT 13.73 0.88 13.86 1.01 ;
 RECT 10.67 1.63 10.8 1.76 ;
 RECT 5.455 2.4 5.585 2.53 ;
 RECT 9.05 1.27 9.18 1.4 ;
 RECT 2.435 1.265 2.565 1.395 ;
 RECT 9.41 2.33 9.54 2.46 ;
 RECT 24.71 1.075 24.84 1.205 ;
 RECT 27.56 1.03 27.69 1.16 ;
 RECT 22.82 0.26 22.95 0.39 ;
 RECT 25.635 0.975 25.765 1.105 ;
 RECT 26.42 0.26 26.55 0.39 ;
 RECT 23.66 1.075 23.79 1.205 ;
 RECT 25.155 1.035 25.285 1.165 ;
 RECT 27.595 2.31 27.725 2.44 ;
 RECT 23.4 0.635 23.53 0.765 ;
 RECT 13.075 2.295 13.205 2.425 ;
 RECT 15.765 0.725 15.895 0.855 ;
 RECT 15.095 0.86 15.225 0.99 ;
 RECT 19.43 0.51 19.56 0.64 ;
 RECT 18.505 1.7 18.635 1.83 ;
 RECT 19.01 0.26 19.14 0.39 ;
 RECT 16.38 0.3 16.51 0.43 ;
 LAYER M1 ;
 RECT 25.63 0.73 25.77 0.935 ;
 RECT 25.31 0.355 25.45 0.59 ;
 RECT 25.31 1.345 25.77 1.485 ;
 RECT 25.585 0.935 25.815 1.145 ;
 RECT 25.31 0.59 25.77 0.73 ;
 RECT 23.61 1.225 23.84 1.245 ;
 RECT 23.61 1.195 24.2 1.225 ;
 RECT 23.75 1.015 24.06 1.035 ;
 RECT 23.61 1.035 24.06 1.055 ;
 RECT 23.885 0.64 24.025 1.015 ;
 RECT 24.06 1.225 24.2 1.75 ;
 RECT 23.765 0.5 24.025 0.64 ;
 RECT 24.66 1.035 24.89 1.055 ;
 RECT 24.66 1.195 24.89 1.245 ;
 RECT 23.61 1.055 24.89 1.195 ;
 RECT 22.77 0.36 23 0.43 ;
 RECT 24.165 0.36 24.305 0.565 ;
 RECT 22.77 0.22 24.305 0.36 ;
 RECT 24.905 0.705 25.045 0.75 ;
 RECT 25.03 0.995 25.335 1.205 ;
 RECT 25.03 0.89 25.17 0.995 ;
 RECT 24.905 0.75 25.17 0.89 ;
 RECT 24.165 0.565 25.045 0.705 ;
 RECT 19.38 0.475 19.985 0.625 ;
 RECT 19.38 0.47 19.61 0.475 ;
 RECT 19.38 0.635 19.61 0.68 ;
 RECT 20.765 0.37 20.905 0.625 ;
 RECT 19.38 0.625 20.905 0.635 ;
 RECT 19.845 0.635 20.905 0.765 ;
 RECT 20.765 0.765 20.905 0.77 ;
 RECT 21.665 0.37 21.805 1.46 ;
 RECT 20.765 0.23 21.805 0.37 ;
 RECT 15.045 0.82 15.275 0.855 ;
 RECT 15.045 0.995 15.275 1.03 ;
 RECT 14.755 0.525 14.895 0.855 ;
 RECT 14.755 0.995 14.895 2.065 ;
 RECT 14.755 0.855 15.275 0.995 ;
 RECT 11.48 0.82 11.62 2.33 ;
 RECT 12.33 1.975 12.47 2.33 ;
 RECT 12.33 2.47 12.47 2.475 ;
 RECT 11.48 2.47 11.62 2.475 ;
 RECT 11.48 2.33 12.47 2.47 ;
 RECT 13.41 1.975 13.55 2.295 ;
 RECT 13.725 0.765 13.865 2.295 ;
 RECT 14.25 0.525 14.39 2.295 ;
 RECT 12.33 1.835 13.55 1.975 ;
 RECT 13.41 2.295 14.39 2.435 ;
 RECT 16.655 0.22 18.035 0.36 ;
 RECT 16.655 0.36 16.885 0.68 ;
 RECT 17.895 0.36 18.035 0.675 ;
 RECT 15.72 0.68 16.885 0.685 ;
 RECT 15.72 0.895 16.885 0.91 ;
 RECT 15.715 0.685 16.885 0.895 ;
 RECT 17.895 0.675 19.22 0.815 ;
 RECT 18.96 0.23 19.22 0.43 ;
 RECT 18.96 0.22 19.19 0.23 ;
 RECT 19.08 0.43 19.22 0.675 ;
 RECT 19.08 0.815 19.22 1.98 ;
 RECT 15.42 0.385 15.56 1.05 ;
 RECT 13.19 0.385 13.33 0.99 ;
 RECT 12.215 0.99 13.33 1.13 ;
 RECT 13.19 0.245 15.56 0.385 ;
 RECT 12.215 0.36 12.355 0.99 ;
 RECT 10.315 0.22 12.355 0.36 ;
 RECT 10.315 0.36 10.455 0.655 ;
 RECT 9.38 0.655 10.455 0.795 ;
 RECT 9.38 0.35 9.71 0.655 ;
 RECT 17.03 0.555 17.295 0.74 ;
 RECT 17.065 0.53 17.295 0.555 ;
 RECT 17.03 0.74 17.17 1.05 ;
 RECT 15.42 1.05 17.17 1.19 ;
 RECT 8.595 0.565 8.845 0.66 ;
 RECT 9.1 0.565 9.24 0.945 ;
 RECT 8.595 0.425 9.24 0.565 ;
 RECT 10.6 0.505 10.985 0.71 ;
 RECT 10.6 0.71 10.74 0.945 ;
 RECT 10.755 0.5 10.985 0.505 ;
 RECT 9.1 0.945 10.74 1.085 ;
 RECT 4.675 0.59 4.815 1.925 ;
 RECT 7.91 0.5 8.165 0.965 ;
 RECT 7.91 1.67 8.05 1.82 ;
 RECT 7.91 0.965 8.05 1.44 ;
 RECT 7.91 1.44 8.165 1.67 ;
 RECT 7.78 1.82 8.05 1.96 ;
 RECT 6.125 1.01 6.265 1.195 ;
 RECT 6.125 1.335 6.265 1.67 ;
 RECT 6.06 0.87 6.33 1.01 ;
 RECT 6.05 1.67 6.33 1.81 ;
 RECT 6.125 1.195 7.015 1.335 ;
 RECT 6.875 0.67 7.015 1.195 ;
 RECT 8.305 0.36 8.445 1.895 ;
 RECT 7.62 0.22 8.445 0.36 ;
 RECT 6.875 0.53 7.76 0.67 ;
 RECT 8.26 1.895 8.445 2.17 ;
 RECT 7.62 0.36 7.76 0.53 ;
 RECT 5.145 0.685 5.285 1.925 ;
 RECT 5.145 0.545 6.455 0.615 ;
 RECT 6.09 0.22 6.455 0.545 ;
 RECT 5.145 0.615 6.45 0.685 ;
 RECT 3.555 0.915 3.695 1.875 ;
 RECT 3.44 1.875 3.695 2.175 ;
 RECT 3.555 0.845 3.845 0.915 ;
 RECT 3.555 0.705 4.535 0.845 ;
 RECT 4.395 0.37 4.535 0.705 ;
 RECT 5.305 0.37 5.585 0.395 ;
 RECT 4.395 0.23 5.585 0.37 ;
 RECT 1.32 0.88 1.65 1.01 ;
 RECT 1.32 1.01 1.605 1.02 ;
 RECT 1.51 0.74 1.65 0.88 ;
 RECT 2.335 0.74 2.475 1.075 ;
 RECT 1.51 0.6 2.475 0.74 ;
 RECT 0.24 0.84 0.38 1.96 ;
 RECT 0.31 2.1 0.45 2.545 ;
 RECT 0.465 0.56 0.605 0.7 ;
 RECT 0.24 1.96 0.65 2.1 ;
 RECT 0.24 0.7 0.66 0.84 ;
 RECT 0.465 0.42 2.755 0.455 ;
 RECT 2.615 0.455 2.755 1.215 ;
 RECT 0.465 0.455 1.37 0.56 ;
 RECT 1.215 0.315 2.755 0.42 ;
 RECT 2.385 1.215 2.755 1.435 ;
 RECT 15.28 2.42 15.51 2.54 ;
 RECT 22.76 2.42 22.9 2.52 ;
 RECT 15.28 2.28 22.9 2.42 ;
 RECT 27.545 2.48 27.685 2.52 ;
 RECT 27.545 2.27 27.775 2.48 ;
 RECT 22.76 2.52 27.685 2.66 ;
 RECT 17.32 0.905 17.46 1.37 ;
 RECT 17.32 1.51 17.46 1.7 ;
 RECT 16.38 1.51 16.52 1.695 ;
 RECT 18.705 1.25 18.935 1.37 ;
 RECT 16.38 1.37 18.935 1.51 ;
 RECT 17.255 1.7 17.53 1.84 ;
 RECT 16.31 1.695 16.59 1.835 ;
 RECT 15.415 1.565 15.555 1.985 ;
 RECT 15.415 1.985 18.685 2.125 ;
 RECT 18.455 1.66 18.685 1.985 ;
 RECT 15.37 1.355 15.6 1.565 ;
 RECT 10.055 2.115 10.195 2.325 ;
 RECT 9.16 1.975 10.26 2.115 ;
 RECT 8.685 1.81 8.965 2.115 ;
 RECT 8.6 1.015 8.74 1.67 ;
 RECT 8.595 0.875 8.96 1.015 ;
 RECT 8.6 1.67 10.855 1.81 ;
 RECT 10.615 1.58 10.855 1.67 ;
 RECT 10.615 1.81 10.855 1.835 ;
 RECT 11.765 1.41 12.065 1.455 ;
 RECT 11.925 0.81 12.065 1.41 ;
 RECT 11.765 1.595 12.065 1.62 ;
 RECT 11.925 1.62 12.065 2.18 ;
 RECT 12.675 1.415 12.815 1.455 ;
 RECT 11.765 1.455 12.815 1.595 ;
 RECT 12.675 1.275 13.195 1.415 ;
 RECT 9 1.37 9.23 1.44 ;
 RECT 10.995 0.865 11.135 1.23 ;
 RECT 8.99 1.23 11.135 1.37 ;
 RECT 10.995 1.37 11.135 2.215 ;
 RECT 7.115 1.63 7.255 1.915 ;
 RECT 7.2 0.825 7.34 1.475 ;
 RECT 7.115 1.475 7.46 1.63 ;
 RECT 7.005 1.915 7.255 2.055 ;
 RECT 1.395 1.895 1.535 2.38 ;
 RECT 1.395 2.38 2.475 2.52 ;
 RECT 2.335 1.895 2.475 2.38 ;
 RECT 2.055 1.02 2.195 1.585 ;
 RECT 2.055 1.725 2.195 1.815 ;
 RECT 1.865 1.955 2.005 2.17 ;
 RECT 1.79 0.88 2.195 1.02 ;
 RECT 1.865 1.815 2.195 1.955 ;
 RECT 3.835 2.22 3.975 2.315 ;
 RECT 2.055 1.585 3.285 1.725 ;
 RECT 3.145 1.725 3.285 2.315 ;
 RECT 3.145 2.315 3.975 2.455 ;
 RECT 3.835 2.08 5.565 2.22 ;
 RECT 5.615 0.835 5.755 0.845 ;
 RECT 5.615 0.845 5.91 0.985 ;
 RECT 5.615 0.985 5.755 1.795 ;
 RECT 5.425 1.795 5.82 1.935 ;
 RECT 5.425 1.935 5.565 2.08 ;
 RECT 26.25 0.73 26.39 1.04 ;
 RECT 26.39 1.18 26.53 1.605 ;
 RECT 26.185 0.59 26.46 0.73 ;
 RECT 27.51 0.99 27.74 1.04 ;
 RECT 26.25 1.04 27.74 1.18 ;
 RECT 27.51 1.18 27.74 1.2 ;
 RECT 26.37 0.29 26.74 0.43 ;
 RECT 26.6 0.43 26.74 0.71 ;
 RECT 26.37 0.22 26.6 0.29 ;
 RECT 28.02 0.85 28.16 1.385 ;
 RECT 27.705 1.525 27.845 1.73 ;
 RECT 26.6 0.71 28.16 0.85 ;
 RECT 27.705 0.51 27.845 0.71 ;
 RECT 27.705 1.385 28.16 1.525 ;
 RECT 25.63 1.145 25.77 1.345 ;
 RECT 25.31 1.485 25.45 1.76 ;
 END
END RSDFFSRSSRX1

MACRO RSDFFSRSSRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 31.68 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 31.68 0.08 ;
 RECT 28.545 0.08 28.785 0.26 ;
 RECT 20.215 0.345 20.48 0.485 ;
 RECT 21.155 0.345 21.46 0.485 ;
 RECT 4.115 0.08 4.255 0.565 ;
 RECT 3.15 0.08 3.29 0.445 ;
 RECT 6.595 0.08 6.735 1.055 ;
 RECT 7.34 0.08 7.48 0.39 ;
 RECT 9.94 0.08 10.175 0.515 ;
 RECT 12.815 0.08 12.955 0.815 ;
 RECT 16.375 0.08 16.515 0.5 ;
 RECT 18.18 0.08 18.32 0.525 ;
 RECT 26.195 0.08 26.335 0.36 ;
 RECT 22.935 0.08 23.075 0.815 ;
 RECT 27.41 0.08 27.55 0.35 ;
 RECT 0.65 0.08 0.92 0.245 ;
 RECT 20.29 0.08 20.43 0.345 ;
 RECT 21.24 0.08 21.38 0.345 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 31.68 2.96 ;
 RECT 2.83 1.87 2.97 2.8 ;
 RECT 9.33 2.29 9.59 2.545 ;
 RECT 4.115 1.975 4.255 2.8 ;
 RECT 0.925 1.89 1.065 2.8 ;
 RECT 7.27 2.59 7.52 2.8 ;
 RECT 6.53 2.59 6.78 2.8 ;
 RECT 10.525 2.07 10.665 2.8 ;
 RECT 16.85 2.57 16.99 2.8 ;
 RECT 20.26 2.565 20.4 2.8 ;
 RECT 21.26 2.565 21.4 2.8 ;
 RECT 18.175 2.57 18.315 2.8 ;
 RECT 22.85 2.565 22.99 2.8 ;
 RECT 23.905 2.565 24.045 2.8 ;
 RECT 12.565 2.625 12.83 2.8 ;
 RECT 9.405 2.545 9.545 2.8 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.58 1.475 6.975 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.905 1.55 13.24 2.04 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 29.995 1.58 30.445 1.8 ;
 RECT 30.105 1.435 30.445 1.58 ;
 RECT 26.195 1.9 28.565 1.99 ;
 RECT 28.27 2.04 30.135 2.13 ;
 RECT 26.195 1.99 30.135 2.04 ;
 RECT 28.425 1.435 28.565 1.9 ;
 RECT 26.195 1.39 26.335 1.9 ;
 RECT 27.58 1.37 27.72 1.9 ;
 RECT 29.995 1.8 30.135 1.99 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 24.805 0.59 25.09 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.985 1.03 4.52 1.525 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.955 2.12 6.205 2.41 ;
 RECT 5.4 2.55 5.63 2.585 ;
 RECT 5.4 2.41 6.205 2.55 ;
 RECT 5.4 2.375 5.63 2.41 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.905 0.84 3.325 1.09 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END RSTB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 1.47 1.915 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 2.285 0.775 2.505 ;
 RECT 0.2 2.115 0.445 2.285 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.215 1.47 22.52 1.77 ;
 RECT 22.375 0.545 22.515 1.47 ;
 RECT 22.375 1.995 24.515 2.135 ;
 RECT 23.365 1.705 23.64 1.845 ;
 RECT 22.375 1.77 22.515 1.995 ;
 RECT 24.375 1.695 24.515 1.995 ;
 RECT 23.435 1.845 23.575 1.995 ;
 RECT 23.435 0.555 23.575 1.705 ;
 END
 ANTENNADIFFAREA 0.848 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 21.64 1.16 21.88 1.4 ;
 RECT 21.71 0.91 21.85 1.16 ;
 RECT 19.81 1.955 21.85 2.095 ;
 RECT 21.71 1.4 21.85 1.955 ;
 RECT 19.81 2.095 19.95 2.1 ;
 RECT 19.81 0.91 19.95 1.955 ;
 RECT 20.77 0.91 20.91 1.955 ;
 END
 ANTENNADIFFAREA 0.886 ;
 END Q

 OBS
 LAYER PO ;
 RECT 15.045 0.82 15.275 0.875 ;
 RECT 15.045 0.975 15.275 1.03 ;
 RECT 15.045 0.875 15.95 0.975 ;
 RECT 18.43 1.635 18.53 1.66 ;
 RECT 18.43 1.66 18.685 1.87 ;
 RECT 18.43 1.87 18.53 2.565 ;
 RECT 20.075 0.19 20.175 1.27 ;
 RECT 21.025 0.48 21.125 1.27 ;
 RECT 21.025 1.37 21.125 2.265 ;
 RECT 20.555 0.495 20.655 1.27 ;
 RECT 20.555 1.37 20.655 2.305 ;
 RECT 21.495 0.49 21.595 1.27 ;
 RECT 21.495 1.37 21.595 2.265 ;
 RECT 20.075 1.37 20.175 2.315 ;
 RECT 19.09 0.19 19.19 0.22 ;
 RECT 20.075 1.27 21.595 1.37 ;
 RECT 19.09 0.09 20.175 0.19 ;
 RECT 18.96 0.22 19.19 0.43 ;
 RECT 18.705 1.25 18.965 1.3 ;
 RECT 18.865 0.61 18.965 1.25 ;
 RECT 18.705 1.4 18.965 1.46 ;
 RECT 18.865 1.46 18.965 2.56 ;
 RECT 19.395 0.68 19.495 1.3 ;
 RECT 18.705 1.3 19.495 1.4 ;
 RECT 19.38 0.47 19.61 0.68 ;
 RECT 17.105 0.51 17.205 0.53 ;
 RECT 17.105 0.74 17.205 2.21 ;
 RECT 17.065 0.53 17.295 0.74 ;
 RECT 16.635 0.54 16.885 0.695 ;
 RECT 16.635 0.695 16.735 2.21 ;
 RECT 16.655 0.485 16.885 0.54 ;
 RECT 13.47 2.69 15.38 2.695 ;
 RECT 15.28 2.54 15.38 2.69 ;
 RECT 14.26 2.695 15.38 2.79 ;
 RECT 13.47 0.66 13.57 2.595 ;
 RECT 13.47 2.595 14.36 2.69 ;
 RECT 15.28 2.33 15.51 2.54 ;
 RECT 14.505 1.355 15.6 1.39 ;
 RECT 14.505 0.19 14.605 1.29 ;
 RECT 14.505 1.29 15.595 1.355 ;
 RECT 8.015 0.19 8.115 0.51 ;
 RECT 9.75 0.19 9.85 1.24 ;
 RECT 15.37 1.39 15.6 1.565 ;
 RECT 7.975 0.51 8.22 0.755 ;
 RECT 8.015 0.09 14.605 0.19 ;
 RECT 15.075 1.71 15.175 1.76 ;
 RECT 10.8 0.48 10.985 0.5 ;
 RECT 18.435 0.19 18.535 1.18 ;
 RECT 16.135 0.19 16.235 1.76 ;
 RECT 15.075 1.76 16.235 1.86 ;
 RECT 13.99 0.48 14.09 1.61 ;
 RECT 14.54 1.71 14.64 2.445 ;
 RECT 16.135 0.09 18.535 0.19 ;
 RECT 13.99 1.61 15.175 1.71 ;
 RECT 10.8 0.38 14.09 0.48 ;
 RECT 10.755 0.5 10.985 0.71 ;
 RECT 11.255 1.575 11.355 2.485 ;
 RECT 11.765 1.41 11.995 1.475 ;
 RECT 11.765 1.575 11.995 1.62 ;
 RECT 11.255 1.475 11.995 1.575 ;
 RECT 4.93 1.495 5.03 2.365 ;
 RECT 3.385 2.365 5.03 2.465 ;
 RECT 3.385 1.88 3.615 2.365 ;
 RECT 1.65 0.66 1.75 1.48 ;
 RECT 1.65 1.715 1.75 2.38 ;
 RECT 1.605 1.48 1.835 1.715 ;
 RECT 4.46 0.555 4.56 1.035 ;
 RECT 4.46 1.27 4.56 2.185 ;
 RECT 4.18 1.035 4.56 1.27 ;
 RECT 5.325 0.16 5.59 0.465 ;
 RECT 5.49 0.465 5.59 1.13 ;
 RECT 10.615 1.61 10.88 1.82 ;
 RECT 10.78 1.82 10.88 2.49 ;
 RECT 10.41 0.66 10.51 1.51 ;
 RECT 10.41 1.51 10.88 1.61 ;
 RECT 13.075 0.66 13.175 1.205 ;
 RECT 12.46 1.305 12.69 1.475 ;
 RECT 12.46 1.205 13.175 1.305 ;
 RECT 6.855 0.655 6.955 1.495 ;
 RECT 6.66 1.495 6.955 1.745 ;
 RECT 6.855 1.745 6.955 2.19 ;
 RECT 6.14 0.27 6.48 0.52 ;
 RECT 6.38 0.52 6.48 2.31 ;
 RECT 8.515 1.595 8.615 2.33 ;
 RECT 7.975 1.445 8.22 1.495 ;
 RECT 7.975 1.495 8.615 1.595 ;
 RECT 7.975 1.595 8.22 1.69 ;
 RECT 7.695 1.265 7.795 1.52 ;
 RECT 7.195 1.52 7.795 1.62 ;
 RECT 7.63 1.62 7.73 2.69 ;
 RECT 10.31 1.79 10.41 2.69 ;
 RECT 7.195 1.44 7.44 1.52 ;
 RECT 7.195 1.62 7.44 1.69 ;
 RECT 8.56 0.375 8.845 0.61 ;
 RECT 8.56 0.61 8.66 1.165 ;
 RECT 7.695 0.585 7.795 1.165 ;
 RECT 7.63 2.69 10.41 2.79 ;
 RECT 7.695 1.165 8.66 1.265 ;
 RECT 5.4 1.41 5.5 2.375 ;
 RECT 5.21 1.31 5.5 1.41 ;
 RECT 4.93 0.23 5.03 1.21 ;
 RECT 3.9 0.23 4 2.185 ;
 RECT 4.93 1.21 5.31 1.31 ;
 RECT 3.9 0.13 5.03 0.23 ;
 RECT 5.4 2.375 5.63 2.585 ;
 RECT 13.04 1.76 13.14 2.48 ;
 RECT 12.18 1.23 12.28 1.655 ;
 RECT 12.18 1.755 12.28 2.57 ;
 RECT 11.265 0.66 11.365 1.13 ;
 RECT 12.18 0.66 12.28 1.13 ;
 RECT 12.91 1.55 13.14 1.655 ;
 RECT 12.91 1.755 13.14 1.76 ;
 RECT 12.18 1.655 13.14 1.755 ;
 RECT 11.265 1.13 12.28 1.23 ;
 RECT 0.545 2.285 0.81 2.495 ;
 RECT 0.71 0.48 0.81 2.285 ;
 RECT 1.18 1.75 1.28 2.69 ;
 RECT 1.05 1.54 1.28 1.75 ;
 RECT 2.815 0.48 2.915 0.87 ;
 RECT 1.18 0.48 1.28 1.24 ;
 RECT 2.815 1.08 2.915 1.625 ;
 RECT 2.12 1.725 2.22 2.775 ;
 RECT 2.815 0.87 3.135 1.08 ;
 RECT 1.18 0.38 2.915 0.48 ;
 RECT 2.12 1.625 2.915 1.725 ;
 RECT 22.635 1.325 24.26 1.425 ;
 RECT 23.215 1.425 23.315 2.645 ;
 RECT 23.855 0.45 23.955 1.325 ;
 RECT 23.215 0.375 23.315 1.325 ;
 RECT 22.635 1.425 22.735 2.62 ;
 RECT 24.16 1.425 24.26 2.645 ;
 RECT 23.69 1.425 23.79 2.64 ;
 RECT 22.635 0.38 22.735 1.12 ;
 RECT 22.635 1.12 22.885 1.325 ;
 RECT 23.7 0.22 24.11 0.45 ;
 RECT 9.05 0.65 9.15 1.23 ;
 RECT 9.01 1.44 9.11 2.33 ;
 RECT 9 1.23 9.23 1.44 ;
 RECT 2.12 0.66 2.22 1.195 ;
 RECT 2.385 1.43 2.615 1.435 ;
 RECT 2.12 1.195 2.63 1.43 ;
 RECT 9.45 0.6 9.55 1.61 ;
 RECT 9.485 1.71 9.585 2.285 ;
 RECT 9.33 0.37 9.57 0.6 ;
 RECT 9.45 1.61 9.585 1.71 ;
 RECT 9.36 2.285 9.59 2.5 ;
 RECT 26.455 1.245 26.555 2.02 ;
 RECT 26.325 1.035 26.555 1.245 ;
 RECT 27.67 0.38 27.77 0.96 ;
 RECT 27.67 1.06 27.77 1.14 ;
 RECT 27.25 0.935 27.48 0.96 ;
 RECT 27.25 0.96 27.77 1.06 ;
 RECT 27.25 1.06 27.48 1.145 ;
 RECT 27.67 1.14 27.94 1.24 ;
 RECT 27.84 1.24 27.94 1.84 ;
 RECT 28.035 0.22 28.265 0.28 ;
 RECT 28.035 0.38 28.265 0.43 ;
 RECT 27.67 0.28 28.265 0.38 ;
 RECT 29.85 0.195 29.95 2.665 ;
 RECT 28.845 0.095 29.95 0.195 ;
 RECT 25.065 1.245 25.165 2.665 ;
 RECT 25.065 1.2 25.35 1.245 ;
 RECT 28.845 0.195 28.945 0.945 ;
 RECT 25.065 2.665 29.95 2.765 ;
 RECT 25.12 1.035 25.35 1.1 ;
 RECT 25.065 1.1 25.395 1.2 ;
 RECT 26.76 0.215 26.86 0.995 ;
 RECT 26.76 0.995 27 1.205 ;
 RECT 26.76 1.205 26.86 2 ;
 RECT 29.155 0.375 29.255 0.99 ;
 RECT 29.155 0.99 29.405 1.2 ;
 RECT 29.155 1.2 29.255 2.27 ;
 RECT 29 2.27 29.285 2.48 ;
 RECT 25.975 1.87 26.08 1.97 ;
 RECT 25.98 0.855 26.08 1.87 ;
 RECT 25.975 1.97 26.075 2.2 ;
 RECT 28.69 1.125 28.79 2.2 ;
 RECT 25.975 2.2 28.79 2.3 ;
 RECT 26.45 0.215 26.55 0.755 ;
 RECT 25.98 0.21 26.08 0.755 ;
 RECT 24.86 0.595 25.09 0.755 ;
 RECT 24.86 0.755 26.55 0.855 ;
 RECT 15.715 0.685 15.945 0.875 ;
 LAYER CO ;
 RECT 15.33 2.37 15.46 2.5 ;
 RECT 15.42 1.395 15.55 1.525 ;
 RECT 10.805 0.54 10.935 0.67 ;
 RECT 11.815 1.45 11.945 1.58 ;
 RECT 0.72 0.11 0.85 0.24 ;
 RECT 5.15 0.78 5.28 0.91 ;
 RECT 1.87 1.965 2 2.095 ;
 RECT 0.93 1.965 1.06 2.095 ;
 RECT 3.56 1.49 3.69 1.62 ;
 RECT 1.655 1.535 1.785 1.665 ;
 RECT 4.68 0.78 4.81 0.91 ;
 RECT 4.12 0.35 4.25 0.48 ;
 RECT 3.445 1.94 3.575 2.07 ;
 RECT 4.68 1.725 4.81 1.855 ;
 RECT 28.06 1.405 28.19 1.535 ;
 RECT 25.325 0.505 25.455 0.635 ;
 RECT 26.98 1.485 27.11 1.615 ;
 RECT 27.415 0.12 27.545 0.25 ;
 RECT 28.43 1.49 28.56 1.62 ;
 RECT 26.2 1.475 26.33 1.605 ;
 RECT 27.585 1.445 27.715 1.575 ;
 RECT 28.595 0.12 28.725 0.25 ;
 RECT 29.375 1.465 29.505 1.595 ;
 RECT 26.2 0.135 26.33 0.265 ;
 RECT 30.155 1.475 30.285 1.605 ;
 RECT 26.98 0.435 27.11 0.565 ;
 RECT 29.375 0.595 29.505 0.725 ;
 RECT 25.73 1.425 25.86 1.555 ;
 RECT 27.92 0.595 28.05 0.725 ;
 RECT 14.76 1.87 14.89 2 ;
 RECT 14.255 0.595 14.385 0.725 ;
 RECT 14.255 1.9 14.385 2.03 ;
 RECT 21.265 2.635 21.395 2.765 ;
 RECT 20.775 0.97 20.905 1.1 ;
 RECT 21.715 1.705 21.845 1.835 ;
 RECT 19.815 1.705 19.945 1.835 ;
 RECT 23.44 1.705 23.57 1.835 ;
 RECT 4.12 2.045 4.25 2.175 ;
 RECT 23.44 0.625 23.57 0.755 ;
 RECT 22.38 0.62 22.51 0.75 ;
 RECT 21.245 0.35 21.375 0.48 ;
 RECT 20.265 2.635 20.395 2.765 ;
 RECT 22.38 1.72 22.51 1.85 ;
 RECT 20.775 1.705 20.905 1.835 ;
 RECT 20.295 0.35 20.425 0.48 ;
 RECT 23.91 2.635 24.04 2.765 ;
 RECT 19.815 0.97 19.945 1.1 ;
 RECT 22.855 2.635 22.985 2.765 ;
 RECT 6.6 2.64 6.73 2.77 ;
 RECT 3.645 0.78 3.775 0.91 ;
 RECT 2.34 1.965 2.47 2.095 ;
 RECT 2.835 1.995 2.965 2.125 ;
 RECT 0.46 0.705 0.59 0.835 ;
 RECT 1.87 0.885 2 1.015 ;
 RECT 1.4 0.885 1.53 1.015 ;
 RECT 5.375 0.26 5.505 0.39 ;
 RECT 2.34 0.885 2.47 1.015 ;
 RECT 3.155 0.24 3.285 0.37 ;
 RECT 5.15 1.725 5.28 1.855 ;
 RECT 0.46 1.735 0.59 1.865 ;
 RECT 19.085 0.83 19.215 0.96 ;
 RECT 18.185 0.33 18.315 0.46 ;
 RECT 19.085 1.78 19.215 1.91 ;
 RECT 18.18 2.64 18.31 2.77 ;
 RECT 16.38 0.3 16.51 0.43 ;
 RECT 17.325 0.975 17.455 1.105 ;
 RECT 17.325 1.705 17.455 1.835 ;
 RECT 16.855 2.64 16.985 2.77 ;
 RECT 7.85 1.825 7.98 1.955 ;
 RECT 12.51 1.28 12.64 1.41 ;
 RECT 11 2.015 11.13 2.145 ;
 RECT 11.93 0.88 12.06 1.01 ;
 RECT 13.73 1.945 13.86 2.075 ;
 RECT 12.82 0.62 12.95 0.75 ;
 RECT 9.385 0.42 9.515 0.55 ;
 RECT 8.76 1.925 8.89 2.055 ;
 RECT 6.6 0.875 6.73 1.005 ;
 RECT 9.99 0.325 10.12 0.455 ;
 RECT 8.03 1.49 8.16 1.62 ;
 RECT 8.03 0.555 8.16 0.685 ;
 RECT 8.78 0.88 8.91 1.01 ;
 RECT 6.2 0.325 6.33 0.455 ;
 RECT 6.13 0.875 6.26 1.005 ;
 RECT 10.53 2.135 10.66 2.265 ;
 RECT 7.34 2.64 7.47 2.77 ;
 RECT 11.485 2.07 11.615 2.2 ;
 RECT 6.13 1.675 6.26 1.805 ;
 RECT 9.23 1.98 9.36 2.11 ;
 RECT 7.915 0.905 8.045 1.035 ;
 RECT 8.265 1.96 8.395 2.09 ;
 RECT 7.205 0.875 7.335 1.005 ;
 RECT 9.705 1.675 9.835 1.805 ;
 RECT 6.72 1.55 6.85 1.68 ;
 RECT 7.345 0.21 7.475 0.34 ;
 RECT 10.06 2.125 10.19 2.255 ;
 RECT 7.075 1.92 7.205 2.05 ;
 RECT 8.31 0.88 8.44 1.01 ;
 RECT 11 0.93 11.13 1.06 ;
 RECT 8.665 0.43 8.795 0.56 ;
 RECT 11.93 1.935 12.06 2.065 ;
 RECT 11.485 0.88 11.615 1.01 ;
 RECT 7.255 1.495 7.385 1.625 ;
 RECT 13.73 0.88 13.86 1.01 ;
 RECT 10.67 1.63 10.8 1.76 ;
 RECT 14.76 0.595 14.89 0.725 ;
 RECT 5.45 2.415 5.58 2.545 ;
 RECT 12.96 1.59 13.09 1.72 ;
 RECT 0.595 2.325 0.725 2.455 ;
 RECT 1.1 1.58 1.23 1.71 ;
 RECT 2.955 0.91 3.085 1.04 ;
 RECT 22.705 1.16 22.835 1.29 ;
 RECT 23.93 0.27 24.06 0.4 ;
 RECT 9.05 1.27 9.18 1.4 ;
 RECT 2.435 1.265 2.565 1.395 ;
 RECT 9.41 2.33 9.54 2.46 ;
 RECT 26.375 1.075 26.505 1.205 ;
 RECT 29.225 1.03 29.355 1.16 ;
 RECT 27.3 0.975 27.43 1.105 ;
 RECT 28.085 0.26 28.215 0.39 ;
 RECT 25.17 1.075 25.3 1.205 ;
 RECT 26.82 1.035 26.95 1.165 ;
 RECT 29.105 2.31 29.235 2.44 ;
 RECT 24.91 0.635 25.04 0.765 ;
 RECT 15.765 0.725 15.895 0.855 ;
 RECT 15.095 0.86 15.225 0.99 ;
 RECT 19.43 0.51 19.56 0.64 ;
 RECT 18.505 1.7 18.635 1.83 ;
 RECT 19.01 0.26 19.14 0.39 ;
 RECT 18.755 1.29 18.885 1.42 ;
 RECT 17.115 0.57 17.245 0.7 ;
 RECT 16.705 0.525 16.835 0.655 ;
 RECT 16.385 1.7 16.515 1.83 ;
 RECT 12.63 2.63 12.76 2.76 ;
 RECT 21.715 0.97 21.845 1.1 ;
 RECT 22.94 0.615 23.07 0.745 ;
 RECT 24.38 1.765 24.51 1.895 ;
 RECT 2.835 2.255 2.965 2.385 ;
 RECT 4.265 1.09 4.395 1.22 ;
 RECT 5.62 1.8 5.75 1.93 ;
 RECT 1.4 2.02 1.53 2.15 ;
 RECT 5.71 0.85 5.84 0.98 ;
 LAYER M1 ;
 RECT 29.37 1.385 29.825 1.525 ;
 RECT 27.295 1.145 27.435 1.345 ;
 RECT 26.975 1.485 27.115 1.76 ;
 RECT 27.295 0.73 27.435 0.935 ;
 RECT 26.975 0.355 27.115 0.59 ;
 RECT 26.975 1.345 27.435 1.485 ;
 RECT 27.25 0.935 27.48 1.145 ;
 RECT 26.975 0.59 27.435 0.73 ;
 RECT 25.26 1.015 25.57 1.035 ;
 RECT 25.12 1.035 25.57 1.055 ;
 RECT 25.12 1.195 25.57 1.225 ;
 RECT 25.12 1.225 25.35 1.245 ;
 RECT 25.395 0.64 25.535 1.015 ;
 RECT 25.725 1.195 25.865 1.75 ;
 RECT 25.275 0.5 25.535 0.64 ;
 RECT 26.325 1.035 26.555 1.055 ;
 RECT 26.325 1.195 26.555 1.245 ;
 RECT 25.12 1.055 26.555 1.195 ;
 RECT 23.74 0.36 24.11 0.445 ;
 RECT 25.83 0.36 25.97 0.565 ;
 RECT 23.74 0.22 25.97 0.36 ;
 RECT 26.57 0.705 26.71 0.75 ;
 RECT 26.695 0.995 27 1.205 ;
 RECT 26.695 0.89 26.835 0.995 ;
 RECT 26.57 0.75 26.835 0.89 ;
 RECT 25.83 0.565 26.71 0.705 ;
 RECT 19.38 0.475 19.955 0.63 ;
 RECT 19.38 0.47 19.61 0.475 ;
 RECT 19.38 0.635 19.61 0.68 ;
 RECT 21.78 0.365 21.92 0.63 ;
 RECT 19.38 0.63 21.92 0.635 ;
 RECT 19.75 0.635 21.92 0.77 ;
 RECT 22.655 0.365 22.795 1.12 ;
 RECT 21.78 0.225 22.795 0.365 ;
 RECT 22.655 1.12 22.885 1.33 ;
 RECT 15.045 0.82 15.275 0.855 ;
 RECT 15.045 0.995 15.275 1.03 ;
 RECT 14.755 0.525 14.895 0.855 ;
 RECT 14.755 0.995 14.895 2.065 ;
 RECT 14.755 0.855 15.275 0.995 ;
 RECT 11.48 0.82 11.62 2.295 ;
 RECT 13.725 0.765 13.865 2.295 ;
 RECT 14.25 0.525 14.39 2.295 ;
 RECT 11.48 2.295 14.39 2.435 ;
 RECT 16.655 0.22 18.035 0.36 ;
 RECT 16.655 0.36 16.885 0.68 ;
 RECT 17.895 0.36 18.035 0.675 ;
 RECT 15.72 0.68 16.885 0.685 ;
 RECT 15.72 0.895 16.885 0.91 ;
 RECT 15.715 0.685 16.885 0.895 ;
 RECT 17.895 0.675 19.22 0.815 ;
 RECT 18.96 0.23 19.22 0.43 ;
 RECT 18.96 0.22 19.19 0.23 ;
 RECT 19.08 0.43 19.22 0.675 ;
 RECT 19.08 0.815 19.22 1.98 ;
 RECT 15.42 0.385 15.56 1.05 ;
 RECT 13.19 0.385 13.33 0.99 ;
 RECT 12.215 0.99 13.33 1.13 ;
 RECT 13.19 0.245 15.56 0.385 ;
 RECT 12.215 0.36 12.355 0.99 ;
 RECT 10.315 0.22 12.355 0.36 ;
 RECT 10.315 0.36 10.455 0.655 ;
 RECT 9.38 0.655 10.455 0.795 ;
 RECT 9.38 0.35 9.71 0.655 ;
 RECT 17.03 0.555 17.295 0.74 ;
 RECT 17.065 0.53 17.295 0.555 ;
 RECT 17.03 0.74 17.17 1.05 ;
 RECT 15.42 1.05 17.17 1.19 ;
 RECT 4.675 0.59 4.815 1.925 ;
 RECT 9.1 0.565 9.24 0.945 ;
 RECT 8.595 0.565 8.845 0.66 ;
 RECT 8.595 0.425 9.24 0.565 ;
 RECT 10.6 0.505 10.985 0.71 ;
 RECT 10.6 0.71 10.74 0.945 ;
 RECT 10.755 0.5 10.985 0.505 ;
 RECT 9.1 0.945 10.74 1.085 ;
 RECT 7.91 0.5 8.165 0.965 ;
 RECT 7.91 1.67 8.05 1.82 ;
 RECT 7.91 0.965 8.05 1.44 ;
 RECT 7.91 1.44 8.165 1.67 ;
 RECT 7.78 1.82 8.05 1.96 ;
 RECT 6.125 1.01 6.265 1.195 ;
 RECT 6.125 1.335 6.265 1.67 ;
 RECT 6.06 0.87 6.33 1.01 ;
 RECT 6.05 1.67 6.33 1.81 ;
 RECT 6.125 1.195 7.015 1.335 ;
 RECT 6.875 0.67 7.015 1.195 ;
 RECT 8.305 0.36 8.445 1.895 ;
 RECT 7.62 0.22 8.445 0.36 ;
 RECT 6.875 0.53 7.76 0.67 ;
 RECT 8.26 1.895 8.445 2.17 ;
 RECT 7.62 0.36 7.76 0.53 ;
 RECT 5.145 0.685 5.285 1.925 ;
 RECT 5.145 0.545 6.455 0.615 ;
 RECT 6.09 0.22 6.455 0.545 ;
 RECT 5.145 0.615 6.45 0.685 ;
 RECT 1.32 0.88 1.65 1.01 ;
 RECT 1.32 1.01 1.605 1.02 ;
 RECT 1.51 0.74 1.65 0.88 ;
 RECT 2.335 0.74 2.475 1.075 ;
 RECT 1.51 0.6 2.475 0.74 ;
 RECT 3.555 0.915 3.695 1.875 ;
 RECT 3.44 1.875 3.695 2.175 ;
 RECT 3.555 0.845 3.845 0.915 ;
 RECT 3.555 0.705 4.535 0.845 ;
 RECT 4.395 0.37 4.535 0.705 ;
 RECT 5.305 0.37 5.585 0.395 ;
 RECT 4.395 0.23 5.585 0.37 ;
 RECT 0.455 0.84 0.595 1.73 ;
 RECT 0.93 0.455 1.36 0.525 ;
 RECT 1.095 1.3 1.235 1.54 ;
 RECT 0.93 0.525 1.07 0.7 ;
 RECT 0.93 0.84 1.07 1.16 ;
 RECT 0.39 0.7 1.07 0.84 ;
 RECT 1.05 1.54 1.28 1.75 ;
 RECT 0.39 1.73 0.65 1.87 ;
 RECT 0.93 1.16 1.235 1.3 ;
 RECT 2.615 0.455 2.755 1.215 ;
 RECT 0.93 0.385 2.755 0.455 ;
 RECT 1.075 0.315 2.755 0.385 ;
 RECT 2.385 1.215 2.755 1.435 ;
 RECT 15.28 2.305 29.285 2.42 ;
 RECT 29.055 2.27 29.285 2.305 ;
 RECT 29.055 2.445 29.285 2.48 ;
 RECT 27.91 2.42 29.285 2.445 ;
 RECT 15.28 2.28 28.215 2.305 ;
 RECT 15.28 2.42 15.51 2.54 ;
 RECT 17.32 0.905 17.46 1.37 ;
 RECT 17.32 1.51 17.46 1.7 ;
 RECT 16.38 1.51 16.52 1.695 ;
 RECT 18.705 1.25 18.935 1.37 ;
 RECT 16.38 1.37 18.935 1.51 ;
 RECT 17.255 1.7 17.53 1.84 ;
 RECT 16.31 1.695 16.59 1.835 ;
 RECT 15.415 1.565 15.555 1.985 ;
 RECT 15.415 1.985 18.685 2.125 ;
 RECT 18.455 1.66 18.685 1.985 ;
 RECT 15.37 1.355 15.6 1.565 ;
 RECT 11.765 1.415 12.065 1.62 ;
 RECT 11.925 1.62 12.065 2.135 ;
 RECT 11.925 0.81 12.065 1.275 ;
 RECT 11.925 1.275 12.69 1.41 ;
 RECT 11.765 1.41 12.69 1.415 ;
 RECT 10.055 2.115 10.195 2.325 ;
 RECT 9.16 1.975 10.26 2.115 ;
 RECT 7.115 1.63 7.255 1.915 ;
 RECT 7.115 1.475 7.46 1.63 ;
 RECT 7.2 0.825 7.34 1.475 ;
 RECT 7.005 1.915 7.255 2.055 ;
 RECT 8.685 1.81 8.965 2.115 ;
 RECT 8.6 1.015 8.74 1.67 ;
 RECT 8.595 0.875 8.96 1.015 ;
 RECT 10.615 1.58 10.855 1.67 ;
 RECT 10.615 1.81 10.855 1.835 ;
 RECT 8.6 1.67 10.855 1.81 ;
 RECT 9 1.37 9.23 1.44 ;
 RECT 10.995 0.865 11.135 1.23 ;
 RECT 8.99 1.23 11.135 1.37 ;
 RECT 10.995 1.37 11.135 2.215 ;
 RECT 2.055 1.02 2.195 1.585 ;
 RECT 2.055 1.725 2.195 1.96 ;
 RECT 1.79 0.88 2.195 1.02 ;
 RECT 1.8 1.96 2.195 2.1 ;
 RECT 2.055 1.585 3.285 1.725 ;
 RECT 3.835 1.69 3.975 1.695 ;
 RECT 3.835 1.835 3.975 2.315 ;
 RECT 3.145 1.725 3.285 2.315 ;
 RECT 3.835 2.455 3.975 2.46 ;
 RECT 3.145 2.315 3.975 2.455 ;
 RECT 4.395 1.835 4.535 2.08 ;
 RECT 3.835 1.695 4.535 1.835 ;
 RECT 5.615 0.835 5.755 0.845 ;
 RECT 5.615 0.845 5.91 0.985 ;
 RECT 5.615 0.985 5.755 1.795 ;
 RECT 5.425 1.795 5.82 1.935 ;
 RECT 5.425 1.935 5.565 2.08 ;
 RECT 4.395 2.08 5.565 2.22 ;
 RECT 1.395 2.155 1.535 2.38 ;
 RECT 1.395 2.38 2.475 2.52 ;
 RECT 2.335 1.895 2.475 2.38 ;
 RECT 1.33 2.015 1.6 2.155 ;
 RECT 27.915 0.73 28.055 1.04 ;
 RECT 28.055 1.18 28.195 1.605 ;
 RECT 27.85 0.59 28.125 0.73 ;
 RECT 29.175 0.99 29.405 1.04 ;
 RECT 27.915 1.04 29.405 1.18 ;
 RECT 29.175 1.18 29.405 1.2 ;
 RECT 28.035 0.29 28.405 0.43 ;
 RECT 28.265 0.43 28.405 0.71 ;
 RECT 28.035 0.22 28.265 0.29 ;
 RECT 29.685 0.85 29.825 1.385 ;
 RECT 29.37 1.525 29.51 1.73 ;
 RECT 28.265 0.71 29.825 0.85 ;
 RECT 29.37 0.51 29.51 0.71 ;
 END
END RSDFFSRSSRX2

MACRO RSDFFSRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.52 BY 2.88 ;
 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 16.78 1.7 17.925 1.75 ;
 RECT 16.565 1.84 16.92 1.99 ;
 RECT 16.565 1.75 17.925 1.84 ;
 RECT 16.78 0.905 16.92 1.7 ;
 RECT 17.785 0.915 17.925 1.7 ;
 RECT 17.785 1.84 17.925 1.92 ;
 END
 ANTENNADIFFAREA 0.455 ;
 END QN

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.79 1.475 5.12 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.965 1.13 2.105 1.48 ;
 RECT 1.87 1.63 2.815 1.79 ;
 RECT 1.87 1.48 2.115 1.63 ;
 RECT 2.665 1.79 2.805 1.845 ;
 RECT 2.665 1.57 2.805 1.63 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.205 2.12 11.64 2.5 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 25.905 1.41 26.245 1.775 ;
 RECT 24.225 1.965 26.09 2.105 ;
 RECT 21.995 2.195 24.365 2.335 ;
 RECT 24.225 1.41 24.365 1.965 ;
 RECT 25.95 1.775 26.09 1.965 ;
 RECT 23.38 1.345 23.52 2.195 ;
 RECT 21.995 1.365 22.135 2.195 ;
 RECT 24.225 2.105 24.365 2.195 ;
 END
 END VDDG

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.565 0.57 21.045 0.78 ;
 RECT 20.565 0.78 20.935 0.865 ;
 RECT 20.565 0.565 20.935 0.57 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.33 1.155 2.75 1.415 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 27.52 2.96 ;
 RECT 5.415 2.34 5.665 2.8 ;
 RECT 1.36 2.005 1.5 2.8 ;
 RECT 3.27 2.03 3.41 2.8 ;
 RECT 18.78 2.57 18.92 2.8 ;
 RECT 15.205 2.57 15.345 2.8 ;
 RECT 0.385 1.74 0.525 2.8 ;
 RECT 10.77 2.375 10.91 2.8 ;
 RECT 17.265 2.57 17.405 2.8 ;
 RECT 8.67 2.07 8.81 2.8 ;
 RECT 4.74 1.98 4.88 2.8 ;
 RECT 14.36 2.57 14.5 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.08 1.16 18.445 1.4 ;
 RECT 18.305 0.695 18.445 1.16 ;
 RECT 19.365 1.905 19.505 1.91 ;
 RECT 18.305 1.765 19.505 1.905 ;
 RECT 19.365 0.71 19.505 1.765 ;
 RECT 18.305 1.4 18.445 1.765 ;
 END
 ANTENNADIFFAREA 0.717 ;
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 27.52 0.08 ;
 RECT 17.215 0.28 17.48 0.44 ;
 RECT 4.74 0.08 4.88 0.325 ;
 RECT 24.345 0.08 24.585 0.31 ;
 RECT 8.085 0.08 8.32 0.595 ;
 RECT 3.27 0.08 3.41 0.78 ;
 RECT 0.35 0.08 0.49 0.775 ;
 RECT 1.36 0.08 1.5 0.97 ;
 RECT 14.135 0.08 14.275 1.155 ;
 RECT 18.865 0.08 19.005 0.965 ;
 RECT 10.96 0.08 11.1 0.815 ;
 RECT 15.21 0.08 15.35 0.525 ;
 RECT 23.21 0.08 23.35 0.325 ;
 RECT 21.995 0.08 22.135 0.31 ;
 RECT 5.11 0.08 5.25 0.41 ;
 RECT 17.27 0.08 17.41 0.28 ;
 END
 END VSS

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.18 1.475 1.705 1.75 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 OBS
 LAYER PO ;
 RECT 15.735 1.3 16.525 1.4 ;
 RECT 16.41 0.63 16.64 0.84 ;
 RECT 13.85 0.19 13.95 1.795 ;
 RECT 13.85 0.09 15.565 0.19 ;
 RECT 13.155 1.71 13.255 1.795 ;
 RECT 8.945 0.47 9.13 0.5 ;
 RECT 15.465 0.19 15.565 1.18 ;
 RECT 13.155 1.795 13.95 1.895 ;
 RECT 12.685 1.71 12.785 2.445 ;
 RECT 12.135 0.47 12.235 1.61 ;
 RECT 12.135 1.61 13.255 1.71 ;
 RECT 8.945 0.37 12.235 0.47 ;
 RECT 8.9 0.5 9.13 0.71 ;
 RECT 21.02 1.175 21.305 1.305 ;
 RECT 25.655 0.19 25.755 2.64 ;
 RECT 24.645 0.09 25.755 0.19 ;
 RECT 24.645 0.19 24.745 0.94 ;
 RECT 21.02 1.305 21.12 2.64 ;
 RECT 21.02 2.64 25.755 2.74 ;
 RECT 21.02 1.075 21.35 1.175 ;
 RECT 24.955 2.245 25.24 2.455 ;
 RECT 24.955 1.22 25.055 2.245 ;
 RECT 24.955 0.37 25.055 1.01 ;
 RECT 24.955 1.01 25.205 1.22 ;
 RECT 8.76 1.61 9.025 1.82 ;
 RECT 8.925 1.82 9.025 2.49 ;
 RECT 8.555 0.66 8.655 1.51 ;
 RECT 8.555 1.51 9.025 1.61 ;
 RECT 5 0.57 5.1 1.495 ;
 RECT 4.805 1.495 5.1 1.745 ;
 RECT 5 1.745 5.1 2.37 ;
 RECT 1.145 1.475 1.715 1.75 ;
 RECT 1.615 0.555 1.715 1.475 ;
 RECT 1.615 1.75 1.715 2.735 ;
 RECT 1.145 0.555 1.245 1.475 ;
 RECT 1.145 1.75 1.245 2.685 ;
 RECT 5.34 1.52 5.94 1.62 ;
 RECT 6.705 0.47 6.99 0.705 ;
 RECT 6.705 0.705 6.805 1.17 ;
 RECT 5.775 1.62 5.875 2.69 ;
 RECT 8.455 1.79 8.555 2.69 ;
 RECT 5.84 0.685 5.94 1.17 ;
 RECT 5.84 1.17 6.805 1.27 ;
 RECT 5.84 1.27 5.94 1.52 ;
 RECT 5.34 1.44 5.585 1.52 ;
 RECT 5.34 1.62 5.585 1.69 ;
 RECT 5.775 2.69 8.555 2.79 ;
 RECT 4.525 0.52 4.625 2.465 ;
 RECT 4.285 0.27 4.625 0.52 ;
 RECT 11.22 0.655 11.32 1.24 ;
 RECT 10.785 1.205 11.035 1.24 ;
 RECT 10.785 1.34 11.035 1.44 ;
 RECT 10.785 1.24 11.32 1.34 ;
 RECT 19.145 0.365 19.245 1.285 ;
 RECT 18.55 1.285 19.245 1.385 ;
 RECT 19.145 1.385 19.245 2.645 ;
 RECT 19.815 0.365 20.045 0.435 ;
 RECT 19.815 0.2 20.045 0.265 ;
 RECT 19.145 0.265 20.045 0.365 ;
 RECT 18.55 1.2 18.76 1.285 ;
 RECT 18.55 1.385 18.76 1.435 ;
 RECT 18.565 0.47 18.665 1.2 ;
 RECT 18.565 1.435 18.665 2.645 ;
 RECT 17.045 0.39 17.145 1.4 ;
 RECT 16.04 0.29 17.145 0.39 ;
 RECT 16.04 0.225 16.27 0.29 ;
 RECT 16.04 0.39 16.27 0.435 ;
 RECT 17.045 1.5 17.145 2.275 ;
 RECT 17.535 0.505 17.635 1.4 ;
 RECT 17.535 1.5 17.635 2.275 ;
 RECT 17.045 1.4 17.635 1.5 ;
 RECT 2.615 1.59 2.855 1.82 ;
 RECT 2.755 1.82 2.855 2.735 ;
 RECT 11.615 2.69 13.265 2.695 ;
 RECT 13.09 2.54 13.265 2.69 ;
 RECT 12.405 2.695 13.265 2.79 ;
 RECT 11.615 0.655 11.715 2.595 ;
 RECT 11.615 2.595 12.505 2.69 ;
 RECT 13.09 2.33 13.32 2.54 ;
 RECT 7.195 1.295 7.455 1.3 ;
 RECT 7.195 0.65 7.295 1.295 ;
 RECT 7.09 1.55 7.19 2.405 ;
 RECT 7.09 1.3 7.455 1.55 ;
 RECT 10.325 0.655 10.425 1.13 ;
 RECT 10.325 1.23 10.425 1.655 ;
 RECT 9.41 0.66 9.51 1.13 ;
 RECT 10.325 1.655 11.285 1.755 ;
 RECT 11.185 1.755 11.285 2.285 ;
 RECT 10.325 1.755 10.425 2.57 ;
 RECT 11.185 2.285 11.435 2.495 ;
 RECT 9.41 1.13 10.425 1.23 ;
 RECT 12.65 0.19 12.75 1.29 ;
 RECT 12.65 1.29 13.67 1.39 ;
 RECT 7.895 0.19 7.995 2.25 ;
 RECT 13.44 1.285 13.67 1.29 ;
 RECT 13.44 1.39 13.67 1.615 ;
 RECT 7.895 2.46 7.995 2.475 ;
 RECT 7.895 0.09 12.75 0.19 ;
 RECT 7.765 2.25 7.995 2.46 ;
 RECT 6.615 1.67 6.715 2.405 ;
 RECT 6.12 1.46 6.35 1.57 ;
 RECT 6.12 1.57 6.715 1.67 ;
 RECT 22.12 1.01 22.355 1.22 ;
 RECT 22.255 1.22 22.355 1.995 ;
 RECT 21.78 0.87 21.88 2.175 ;
 RECT 20.815 0.77 22.35 0.78 ;
 RECT 21.78 0.73 22.35 0.77 ;
 RECT 24.48 1.125 24.58 2.175 ;
 RECT 20.82 0.78 22.35 0.83 ;
 RECT 20.82 0.83 21.88 0.87 ;
 RECT 22.25 0.19 22.35 0.73 ;
 RECT 21.78 0.185 21.88 0.73 ;
 RECT 20.815 0.57 21.045 0.77 ;
 RECT 21.78 2.175 24.58 2.275 ;
 RECT 14.615 0.64 14.715 1.26 ;
 RECT 14.41 1.26 14.715 1.47 ;
 RECT 14.615 1.47 14.715 2.21 ;
 RECT 22.56 0.19 22.66 0.97 ;
 RECT 22.56 0.97 22.8 1.18 ;
 RECT 22.56 1.18 22.66 1.975 ;
 RECT 15.46 1.635 15.56 1.66 ;
 RECT 15.46 1.66 15.715 1.87 ;
 RECT 15.46 1.87 15.56 2.565 ;
 RECT 3.525 0.335 3.625 1.155 ;
 RECT 3.525 1.365 3.625 2.745 ;
 RECT 3.335 1.155 3.625 1.365 ;
 RECT 1.95 0.555 2.05 1.145 ;
 RECT 1.91 1.145 2.155 1.385 ;
 RECT 2.565 0.555 2.665 1.18 ;
 RECT 2.335 1.41 2.435 1.645 ;
 RECT 2.335 1.18 2.665 1.41 ;
 RECT 2.285 1.645 2.435 1.745 ;
 RECT 2.285 1.745 2.385 2.735 ;
 RECT 23.47 0.355 23.57 0.985 ;
 RECT 23.47 0.255 24.205 0.355 ;
 RECT 23.975 0.355 24.205 0.465 ;
 RECT 23.64 1.215 23.74 1.815 ;
 RECT 23.08 1.115 23.74 1.215 ;
 RECT 23.08 0.985 23.57 1.115 ;
 RECT 2.85 0.175 3.155 0.405 ;
 RECT 3.055 0.405 3.155 2.735 ;
 RECT 9.4 1.575 9.5 2.485 ;
 RECT 9.91 1.41 10.14 1.475 ;
 RECT 9.91 1.575 10.14 1.62 ;
 RECT 9.4 1.475 10.14 1.575 ;
 RECT 15.735 1.25 15.995 1.3 ;
 RECT 15.895 0.61 15.995 1.25 ;
 RECT 16.425 0.84 16.525 1.3 ;
 RECT 15.895 1.46 15.995 2.56 ;
 RECT 15.735 1.4 15.995 1.46 ;
 LAYER CO ;
 RECT 2.31 0.775 2.44 0.905 ;
 RECT 1.37 1.55 1.5 1.68 ;
 RECT 10.775 2.445 10.905 2.575 ;
 RECT 22.78 1.46 22.91 1.59 ;
 RECT 5.485 2.345 5.615 2.475 ;
 RECT 14.14 0.955 14.27 1.085 ;
 RECT 18.31 0.77 18.44 0.9 ;
 RECT 22 0.11 22.13 0.24 ;
 RECT 2.505 2.115 2.635 2.245 ;
 RECT 0.39 2.345 0.52 2.475 ;
 RECT 18.59 1.25 18.72 1.38 ;
 RECT 25.175 0.59 25.305 0.72 ;
 RECT 23.215 0.11 23.345 0.24 ;
 RECT 14.365 2.64 14.495 2.77 ;
 RECT 8.135 0.455 8.265 0.585 ;
 RECT 3.745 2.05 3.875 2.18 ;
 RECT 15.21 2.64 15.34 2.77 ;
 RECT 5.115 0.21 5.245 0.34 ;
 RECT 11.875 0.875 12.005 1.005 ;
 RECT 8.205 2.03 8.335 2.16 ;
 RECT 17.27 2.64 17.4 2.77 ;
 RECT 9.63 2.07 9.76 2.2 ;
 RECT 5.995 1.825 6.125 1.955 ;
 RECT 4.345 0.325 4.475 0.455 ;
 RECT 1.365 2.315 1.495 2.445 ;
 RECT 4.745 0.13 4.875 0.26 ;
 RECT 8.675 2.135 8.805 2.265 ;
 RECT 16.785 1.72 16.915 1.85 ;
 RECT 16.115 1.78 16.245 1.91 ;
 RECT 23.86 1.38 23.99 1.51 ;
 RECT 2.67 1.64 2.8 1.77 ;
 RECT 18.31 1.725 18.44 1.855 ;
 RECT 5.4 1.495 5.53 1.625 ;
 RECT 6.455 0.88 6.585 1.01 ;
 RECT 4.275 0.79 4.405 0.92 ;
 RECT 0.39 1.825 0.52 1.955 ;
 RECT 17.79 1.72 17.92 1.85 ;
 RECT 12.4 0.595 12.53 0.725 ;
 RECT 8.815 1.63 8.945 1.76 ;
 RECT 3.275 2.09 3.405 2.22 ;
 RECT 23.695 0.59 23.825 0.72 ;
 RECT 24.23 1.465 24.36 1.595 ;
 RECT 4.865 1.55 4.995 1.68 ;
 RECT 0.39 2.085 0.52 2.215 ;
 RECT 4.745 2.05 4.875 2.18 ;
 RECT 12.905 1.87 13.035 2 ;
 RECT 9.63 0.88 9.76 1.01 ;
 RECT 24.395 0.115 24.525 0.245 ;
 RECT 21.53 1.4 21.66 1.53 ;
 RECT 10.835 1.245 10.965 1.375 ;
 RECT 6.06 0.905 6.19 1.035 ;
 RECT 9.96 1.45 10.09 1.58 ;
 RECT 16.46 0.67 16.59 0.8 ;
 RECT 8.95 0.54 9.08 0.67 ;
 RECT 21.125 1.135 21.255 1.265 ;
 RECT 25.025 1.05 25.155 1.18 ;
 RECT 15.215 0.33 15.345 0.46 ;
 RECT 6.81 0.525 6.94 0.655 ;
 RECT 18.785 2.64 18.915 2.77 ;
 RECT 10.965 0.62 11.095 0.75 ;
 RECT 12.4 1.9 12.53 2.03 ;
 RECT 7.275 1.345 7.405 1.475 ;
 RECT 23.385 1.42 23.515 1.55 ;
 RECT 19.37 1.71 19.5 1.84 ;
 RECT 17.275 0.305 17.405 0.435 ;
 RECT 1.97 1.195 2.1 1.325 ;
 RECT 0.355 0.59 0.485 0.72 ;
 RECT 25.175 1.44 25.305 1.57 ;
 RECT 14.835 0.96 14.965 1.09 ;
 RECT 5.22 1.995 5.35 2.125 ;
 RECT 6.925 0.88 7.055 1.01 ;
 RECT 2.9 0.225 3.03 0.355 ;
 RECT 11.875 1.945 12.005 2.075 ;
 RECT 10.075 1.885 10.205 2.015 ;
 RECT 2.49 1.23 2.62 1.36 ;
 RECT 22 1.45 22.13 1.58 ;
 RECT 11.255 2.325 11.385 2.455 ;
 RECT 7.815 2.29 7.945 2.42 ;
 RECT 6.17 1.5 6.3 1.63 ;
 RECT 25.06 2.285 25.19 2.415 ;
 RECT 22.17 1.05 22.3 1.18 ;
 RECT 20.865 0.61 20.995 0.74 ;
 RECT 14.46 1.3 14.59 1.43 ;
 RECT 22.62 1.01 22.75 1.14 ;
 RECT 24.025 0.295 24.155 0.425 ;
 RECT 23.13 1.025 23.26 1.155 ;
 RECT 15.785 1.29 15.915 1.42 ;
 RECT 15.535 1.7 15.665 1.83 ;
 RECT 13.49 1.445 13.62 1.575 ;
 RECT 19.865 0.265 19.995 0.395 ;
 RECT 4.275 2.115 4.405 2.245 ;
 RECT 12.905 0.595 13.035 0.725 ;
 RECT 10.075 0.88 10.205 1.01 ;
 RECT 18.87 0.77 19 0.9 ;
 RECT 6.835 2 6.965 2.13 ;
 RECT 3.745 0.775 3.875 0.905 ;
 RECT 0.895 2.055 1.025 2.185 ;
 RECT 16.115 0.83 16.245 0.96 ;
 RECT 9.145 2.015 9.275 2.145 ;
 RECT 7.31 2.04 7.44 2.17 ;
 RECT 1.365 2.055 1.495 2.185 ;
 RECT 0.355 0.33 0.485 0.46 ;
 RECT 13.14 2.37 13.27 2.5 ;
 RECT 16.09 0.265 16.22 0.395 ;
 RECT 3.275 0.585 3.405 0.715 ;
 RECT 3.745 1.79 3.875 1.92 ;
 RECT 21.28 0.505 21.41 0.635 ;
 RECT 3.275 2.35 3.405 2.48 ;
 RECT 1.365 0.775 1.495 0.905 ;
 RECT 19.37 0.78 19.5 0.91 ;
 RECT 9.145 0.93 9.275 1.06 ;
 RECT 22.78 0.41 22.91 0.54 ;
 RECT 25.955 1.45 26.085 1.58 ;
 RECT 0.895 0.775 1.025 0.905 ;
 RECT 5.35 0.97 5.48 1.1 ;
 RECT 14.835 1.705 14.965 1.835 ;
 RECT 3.385 1.195 3.515 1.325 ;
 RECT 16.785 0.975 16.915 1.105 ;
 RECT 17.79 0.975 17.92 1.105 ;
 RECT 6.365 2.035 6.495 2.165 ;
 LAYER M1 ;
 RECT 14.83 1.095 14.97 1.37 ;
 RECT 14.83 1.46 15.96 1.51 ;
 RECT 14.83 1.51 14.97 1.7 ;
 RECT 15.735 1.25 15.965 1.37 ;
 RECT 14.765 1.7 15.04 1.84 ;
 RECT 14.76 0.955 15.03 1.095 ;
 RECT 19.815 0.36 20.045 0.435 ;
 RECT 21.63 0.36 21.77 0.54 ;
 RECT 19.815 0.225 21.77 0.36 ;
 RECT 19.85 0.22 21.77 0.225 ;
 RECT 22.495 0.535 22.635 0.54 ;
 RECT 22.495 0.68 22.635 0.97 ;
 RECT 22.495 0.97 22.8 1.18 ;
 RECT 21.63 0.54 22.635 0.68 ;
 RECT 0.89 0.72 1.03 1.195 ;
 RECT 0.89 1.335 1.03 2.27 ;
 RECT 1.675 0.36 1.815 1.195 ;
 RECT 0.89 1.195 1.815 1.335 ;
 RECT 1.675 0.22 3.1 0.36 ;
 RECT 13.09 2.42 13.32 2.54 ;
 RECT 20.555 2.42 20.695 2.505 ;
 RECT 13.09 2.28 20.695 2.42 ;
 RECT 25.01 2.455 25.15 2.505 ;
 RECT 25.01 2.245 25.24 2.455 ;
 RECT 20.555 2.505 25.15 2.645 ;
 RECT 5.26 1.63 5.4 1.99 ;
 RECT 5.26 1.475 5.605 1.63 ;
 RECT 5.345 0.9 5.485 1.475 ;
 RECT 5.15 1.99 5.4 2.13 ;
 RECT 10.475 2.165 10.615 2.225 ;
 RECT 9.625 0.82 9.765 2.225 ;
 RECT 9.625 2.225 10.615 2.365 ;
 RECT 10.925 1.725 11.065 2.025 ;
 RECT 10.475 2.025 11.065 2.165 ;
 RECT 10.925 2.165 11.065 2.17 ;
 RECT 11.87 2.025 12.535 2.165 ;
 RECT 11.87 1.725 12.01 2.025 ;
 RECT 12.395 0.525 12.535 2.025 ;
 RECT 11.87 0.765 12.01 1.585 ;
 RECT 10.925 1.585 12.01 1.725 ;
 RECT 3.74 0.57 3.88 2.25 ;
 RECT 4.235 0.22 4.6 0.43 ;
 RECT 4.235 0.57 4.6 0.615 ;
 RECT 3.74 0.43 4.6 0.57 ;
 RECT 6.92 0.805 7.06 1.69 ;
 RECT 6.92 1.83 7.06 1.935 ;
 RECT 6.83 1.935 7.06 2.2 ;
 RECT 6.92 1.69 9 1.83 ;
 RECT 8.76 1.58 9 1.69 ;
 RECT 8.76 1.83 9 1.835 ;
 RECT 16.41 0.72 16.64 0.84 ;
 RECT 17.68 0.37 17.82 0.58 ;
 RECT 16.41 0.63 17.82 0.72 ;
 RECT 16.42 0.58 17.82 0.63 ;
 RECT 18.585 0.37 18.725 1.46 ;
 RECT 17.68 0.23 18.725 0.37 ;
 RECT 23.69 0.48 23.83 1.08 ;
 RECT 23.855 1.22 23.995 1.58 ;
 RECT 24.975 1.01 25.205 1.08 ;
 RECT 23.69 1.08 25.205 1.22 ;
 RECT 14.415 0.805 14.555 1.26 ;
 RECT 14.41 1.26 14.64 1.295 ;
 RECT 14.41 1.435 14.64 1.47 ;
 RECT 13.82 1.295 14.64 1.435 ;
 RECT 13.82 1.105 13.96 1.295 ;
 RECT 12.9 0.525 13.04 0.965 ;
 RECT 12.9 1.105 13.04 2.065 ;
 RECT 12.9 0.965 13.96 1.105 ;
 RECT 16.11 0.435 16.25 0.665 ;
 RECT 16.11 0.805 16.25 1.98 ;
 RECT 14.415 0.665 16.25 0.805 ;
 RECT 16.11 0.22 16.25 0.225 ;
 RECT 16.04 0.225 16.27 0.435 ;
 RECT 21.35 0.64 21.49 0.99 ;
 RECT 21.075 1.17 21.665 1.2 ;
 RECT 21.525 1.2 21.665 1.725 ;
 RECT 21.215 0.99 21.525 1.03 ;
 RECT 21.075 1.2 21.305 1.305 ;
 RECT 21.23 0.5 21.49 0.64 ;
 RECT 22.12 1.01 22.35 1.03 ;
 RECT 21.07 1.03 22.35 1.17 ;
 RECT 22.12 1.17 22.35 1.22 ;
 RECT 13.435 1.43 13.67 1.615 ;
 RECT 13.435 1.615 13.575 1.985 ;
 RECT 13.44 1.405 13.67 1.43 ;
 RECT 13.435 1.985 15.67 2.125 ;
 RECT 15.485 1.87 15.67 1.985 ;
 RECT 15.485 1.66 15.715 1.87 ;
 RECT 4.05 1.335 4.19 2.11 ;
 RECT 4.05 0.925 4.19 1.195 ;
 RECT 4.05 2.11 4.475 2.25 ;
 RECT 4.05 0.785 4.475 0.925 ;
 RECT 4.745 0.75 4.885 1.195 ;
 RECT 4.05 1.195 4.885 1.335 ;
 RECT 4.745 0.61 5.56 0.75 ;
 RECT 5.42 0.22 6.59 0.36 ;
 RECT 6.45 0.36 6.59 0.9 ;
 RECT 6.525 1.08 6.665 1.945 ;
 RECT 5.42 0.36 5.56 0.61 ;
 RECT 6.36 2.17 6.5 2.305 ;
 RECT 6.36 1.945 6.665 2.17 ;
 RECT 6.45 0.9 6.665 1.08 ;
 RECT 6.74 0.52 7.34 0.66 ;
 RECT 7.2 0.66 7.34 1.015 ;
 RECT 8.745 0.505 9.13 0.71 ;
 RECT 7.2 1.015 8.885 1.155 ;
 RECT 8.9 0.5 9.13 0.505 ;
 RECT 8.745 0.71 8.885 1.015 ;
 RECT 10.07 1.62 10.21 1.735 ;
 RECT 10.07 1.735 10.785 1.875 ;
 RECT 10.07 1.875 10.21 2.085 ;
 RECT 10.645 1.445 10.785 1.735 ;
 RECT 10.07 0.81 10.21 1.41 ;
 RECT 9.91 1.41 10.21 1.62 ;
 RECT 10.645 1.24 11.04 1.445 ;
 RECT 10.78 1.195 11.04 1.24 ;
 RECT 7.2 1.44 7.465 1.55 ;
 RECT 9.14 0.865 9.28 1.3 ;
 RECT 9.14 1.44 9.28 2.215 ;
 RECT 7.2 1.3 9.28 1.44 ;
 RECT 6.055 1.67 6.195 1.82 ;
 RECT 6.055 1.96 6.195 2.455 ;
 RECT 7.765 2.25 7.995 2.455 ;
 RECT 6.055 0.805 6.195 1.46 ;
 RECT 6.055 1.46 6.35 1.67 ;
 RECT 5.925 1.82 6.195 1.96 ;
 RECT 6.055 2.455 7.995 2.595 ;
 RECT 2.96 0.91 3.1 1.19 ;
 RECT 2.96 1.33 3.1 2.11 ;
 RECT 2.255 0.77 3.1 0.91 ;
 RECT 2.45 2.11 3.1 2.25 ;
 RECT 2.96 1.19 3.52 1.33 ;
 RECT 3.38 1.145 3.52 1.19 ;
 RECT 3.38 1.33 3.52 1.375 ;
 RECT 7.305 2.11 7.445 2.24 ;
 RECT 8.2 2.11 8.34 2.23 ;
 RECT 7.305 1.97 8.34 2.11 ;
 RECT 24.065 0.465 24.205 0.685 ;
 RECT 23.975 0.255 24.205 0.465 ;
 RECT 25.485 0.825 25.625 1.36 ;
 RECT 24.065 0.685 25.625 0.825 ;
 RECT 25.17 1.5 25.31 1.705 ;
 RECT 25.17 0.485 25.31 0.685 ;
 RECT 25.17 1.36 25.625 1.5 ;
 RECT 23.08 1.195 23.22 1.32 ;
 RECT 22.775 1.46 22.915 1.735 ;
 RECT 23.095 0.705 23.235 0.985 ;
 RECT 22.775 0.33 22.915 0.565 ;
 RECT 22.775 1.32 23.22 1.46 ;
 RECT 22.775 0.565 23.235 0.705 ;
 RECT 23.08 0.985 23.31 1.195 ;
 RECT 14.83 1.37 15.965 1.46 ;
 END
END RSDFFSRX1

MACRO RSDFFSRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.84 BY 2.88 ;
 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.265 1.41 26.605 1.775 ;
 RECT 24.72 1.41 24.86 1.965 ;
 RECT 23.875 2.105 24.015 2.11 ;
 RECT 23.875 1.345 24.015 1.965 ;
 RECT 22.49 1.365 22.63 1.965 ;
 RECT 22.49 1.965 26.45 2.105 ;
 RECT 26.31 1.775 26.45 1.965 ;
 END
 END VDDG

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.18 1.475 1.705 1.75 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.79 1.475 5.12 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 16.78 1.7 17.925 1.75 ;
 RECT 16.565 1.84 16.92 1.99 ;
 RECT 16.565 1.75 17.925 1.84 ;
 RECT 16.78 0.905 16.92 1.7 ;
 RECT 17.785 0.915 17.925 1.7 ;
 RECT 17.785 1.84 17.925 1.92 ;
 END
 ANTENNADIFFAREA 0.844 ;
 END QN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.33 1.155 2.75 1.415 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 21.06 0.78 21.43 0.865 ;
 RECT 21.06 0.57 21.54 0.78 ;
 RECT 21.06 0.565 21.43 0.57 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 27.84 0.08 ;
 RECT 17.215 0.28 17.48 0.44 ;
 RECT 8.085 0.08 8.32 0.595 ;
 RECT 24.84 0.08 25.08 0.31 ;
 RECT 4.74 0.08 4.88 0.325 ;
 RECT 3.27 0.08 3.41 0.78 ;
 RECT 5.11 0.08 5.25 0.41 ;
 RECT 0.35 0.08 0.49 0.775 ;
 RECT 10.96 0.08 11.1 0.815 ;
 RECT 15.21 0.08 15.35 0.525 ;
 RECT 1.36 0.08 1.5 0.97 ;
 RECT 14.135 0.08 14.275 1.155 ;
 RECT 18.865 0.08 19.005 0.965 ;
 RECT 19.865 0.08 20.005 0.98 ;
 RECT 23.705 0.08 23.845 0.325 ;
 RECT 22.49 0.08 22.63 0.31 ;
 RECT 17.27 0.08 17.41 0.28 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.305 1.765 20.485 1.905 ;
 RECT 18.08 1.16 18.445 1.4 ;
 RECT 18.305 0.695 18.445 1.16 ;
 RECT 19.365 0.71 19.505 1.765 ;
 RECT 20.345 0.71 20.485 1.765 ;
 RECT 18.305 1.4 18.445 1.765 ;
 END
 ANTENNADIFFAREA 1.137 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 27.84 2.96 ;
 RECT 5.415 2.34 5.665 2.8 ;
 RECT 1.36 2.005 1.5 2.8 ;
 RECT 14.36 2.57 14.5 2.8 ;
 RECT 17.265 2.57 17.405 2.8 ;
 RECT 4.74 1.98 4.88 2.8 ;
 RECT 0.385 1.74 0.525 2.8 ;
 RECT 10.77 2.375 10.91 2.8 ;
 RECT 3.27 2.03 3.41 2.8 ;
 RECT 15.205 2.57 15.345 2.8 ;
 RECT 18.78 2.57 18.92 2.8 ;
 RECT 8.67 2.07 8.81 2.8 ;
 RECT 19.845 2.57 19.985 2.8 ;
 END
 END VDD

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.965 1.13 2.105 1.48 ;
 RECT 1.87 1.63 2.815 1.79 ;
 RECT 1.87 1.48 2.115 1.63 ;
 RECT 2.665 1.79 2.805 1.845 ;
 RECT 2.665 1.57 2.805 1.63 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.08 2.12 11.32 2.475 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 OBS
 LAYER PO ;
 RECT 21.515 1.305 21.615 2.64 ;
 RECT 25.95 0.19 26.05 2.64 ;
 RECT 25.14 0.09 26.05 0.19 ;
 RECT 25.14 0.19 25.24 0.94 ;
 RECT 21.515 2.64 26.05 2.74 ;
 RECT 3.525 0.335 3.625 1.155 ;
 RECT 3.525 1.365 3.625 2.745 ;
 RECT 3.335 1.155 3.625 1.365 ;
 RECT 8.76 1.61 9.025 1.82 ;
 RECT 8.925 1.82 9.025 2.49 ;
 RECT 8.555 0.66 8.655 1.51 ;
 RECT 8.555 1.51 9.025 1.61 ;
 RECT 11.615 2.69 13.265 2.695 ;
 RECT 13.09 2.54 13.265 2.69 ;
 RECT 12.405 2.695 13.265 2.79 ;
 RECT 11.615 0.655 11.715 2.595 ;
 RECT 11.615 2.595 12.505 2.69 ;
 RECT 13.09 2.33 13.32 2.54 ;
 RECT 1.145 1.475 1.715 1.75 ;
 RECT 1.615 0.555 1.715 1.475 ;
 RECT 1.615 1.75 1.715 2.735 ;
 RECT 1.145 0.555 1.245 1.475 ;
 RECT 1.145 1.75 1.245 2.685 ;
 RECT 5 0.57 5.1 1.495 ;
 RECT 4.805 1.495 5.1 1.745 ;
 RECT 5 1.745 5.1 2.37 ;
 RECT 2.85 0.175 3.155 0.405 ;
 RECT 3.055 0.405 3.155 2.735 ;
 RECT 20.13 0.19 20.23 1.285 ;
 RECT 18.55 1.285 20.23 1.385 ;
 RECT 20.13 1.385 20.23 2.645 ;
 RECT 19.63 0.45 19.73 1.285 ;
 RECT 19.63 1.385 19.73 2.645 ;
 RECT 19.145 0.45 19.245 1.285 ;
 RECT 19.145 1.385 19.245 2.645 ;
 RECT 20.585 0.19 20.815 0.435 ;
 RECT 18.55 1.2 18.76 1.285 ;
 RECT 18.55 1.385 18.76 1.435 ;
 RECT 18.565 0.47 18.665 1.2 ;
 RECT 18.565 1.435 18.665 2.645 ;
 RECT 20.13 0.09 20.815 0.19 ;
 RECT 13.85 0.19 13.95 1.795 ;
 RECT 13.85 0.09 15.565 0.19 ;
 RECT 13.155 1.71 13.255 1.795 ;
 RECT 15.465 0.19 15.565 1.18 ;
 RECT 13.155 1.795 13.95 1.895 ;
 RECT 12.685 1.71 12.785 2.445 ;
 RECT 8.945 0.47 9.13 0.5 ;
 RECT 12.135 0.47 12.235 1.61 ;
 RECT 12.135 1.61 13.255 1.71 ;
 RECT 8.945 0.37 12.235 0.47 ;
 RECT 8.9 0.5 9.13 0.71 ;
 RECT 5.775 1.62 5.875 2.69 ;
 RECT 6.705 0.47 6.99 0.705 ;
 RECT 6.705 0.705 6.805 1.17 ;
 RECT 5.84 0.685 5.94 1.17 ;
 RECT 5.84 1.17 6.805 1.27 ;
 RECT 5.84 1.27 5.94 1.52 ;
 RECT 5.34 1.44 5.585 1.52 ;
 RECT 5.34 1.62 5.585 1.69 ;
 RECT 5.34 1.52 5.94 1.62 ;
 RECT 8.455 1.79 8.555 2.69 ;
 RECT 5.775 2.69 8.555 2.79 ;
 RECT 1.95 0.555 2.05 1.145 ;
 RECT 1.91 1.145 2.155 1.385 ;
 RECT 2.565 0.555 2.665 1.18 ;
 RECT 2.335 1.41 2.435 1.645 ;
 RECT 2.335 1.18 2.665 1.41 ;
 RECT 2.285 1.645 2.435 1.745 ;
 RECT 2.285 1.745 2.385 2.735 ;
 RECT 17.045 0.39 17.145 1.4 ;
 RECT 16.04 0.225 16.27 0.29 ;
 RECT 16.04 0.29 17.145 0.39 ;
 RECT 16.04 0.39 16.27 0.435 ;
 RECT 17.045 1.5 17.145 2.65 ;
 RECT 17.535 0.43 17.635 1.4 ;
 RECT 17.535 1.5 17.635 2.65 ;
 RECT 17.045 1.4 17.635 1.5 ;
 RECT 2.755 1.82 2.855 2.735 ;
 RECT 2.615 1.59 2.855 1.82 ;
 RECT 23.965 0.355 24.065 0.985 ;
 RECT 23.965 0.255 24.7 0.355 ;
 RECT 24.47 0.355 24.7 0.465 ;
 RECT 24.135 1.215 24.235 1.815 ;
 RECT 23.575 1.115 24.235 1.215 ;
 RECT 23.575 0.985 24.065 1.115 ;
 RECT 4.285 0.27 4.625 0.52 ;
 RECT 4.525 0.52 4.625 2.465 ;
 RECT 7.195 1.295 7.455 1.3 ;
 RECT 7.195 0.65 7.295 1.295 ;
 RECT 7.09 1.55 7.19 2.405 ;
 RECT 7.09 1.3 7.455 1.55 ;
 RECT 10.325 0.655 10.425 1.13 ;
 RECT 10.325 1.23 10.425 1.655 ;
 RECT 9.41 0.66 9.51 1.13 ;
 RECT 10.325 1.655 11.285 1.755 ;
 RECT 11.185 1.755 11.285 2.255 ;
 RECT 10.325 1.755 10.425 2.57 ;
 RECT 9.41 1.13 10.425 1.23 ;
 RECT 11.085 2.255 11.315 2.465 ;
 RECT 12.65 0.19 12.75 1.29 ;
 RECT 12.65 1.29 13.67 1.39 ;
 RECT 7.895 0.19 7.995 2.25 ;
 RECT 13.44 1.285 13.67 1.29 ;
 RECT 13.44 1.39 13.67 1.615 ;
 RECT 7.895 0.09 12.75 0.19 ;
 RECT 7.765 2.25 7.995 2.46 ;
 RECT 6.615 1.67 6.715 2.405 ;
 RECT 6.12 1.46 6.35 1.57 ;
 RECT 6.12 1.57 6.715 1.67 ;
 RECT 11.22 0.655 11.32 1.24 ;
 RECT 11.09 1.24 11.32 1.475 ;
 RECT 22.275 0.87 22.375 2 ;
 RECT 21.31 0.77 22.845 0.78 ;
 RECT 22.275 0.73 22.845 0.77 ;
 RECT 24.975 1.125 25.075 2 ;
 RECT 21.315 0.78 22.845 0.83 ;
 RECT 21.315 0.83 22.375 0.87 ;
 RECT 22.745 0.19 22.845 0.73 ;
 RECT 22.275 0.185 22.375 0.73 ;
 RECT 21.31 0.57 21.54 0.77 ;
 RECT 22.275 2 25.075 2.1 ;
 RECT 14.615 0.64 14.715 1.26 ;
 RECT 14.41 1.26 14.715 1.47 ;
 RECT 14.615 1.47 14.715 2.21 ;
 RECT 9.4 1.575 9.5 2.485 ;
 RECT 9.91 1.41 10.14 1.475 ;
 RECT 9.91 1.575 10.14 1.62 ;
 RECT 9.4 1.475 10.14 1.575 ;
 RECT 23.055 0.19 23.155 0.97 ;
 RECT 23.055 0.97 23.295 1.18 ;
 RECT 23.055 1.18 23.155 1.81 ;
 RECT 15.735 1.25 15.995 1.3 ;
 RECT 15.895 0.61 15.995 1.25 ;
 RECT 16.425 0.84 16.525 1.3 ;
 RECT 15.895 1.46 15.995 2.56 ;
 RECT 15.735 1.4 15.995 1.46 ;
 RECT 15.735 1.3 16.525 1.4 ;
 RECT 16.41 0.63 16.64 0.84 ;
 RECT 25.45 0.37 25.55 1.01 ;
 RECT 25.45 1.01 25.7 1.22 ;
 RECT 25.45 1.22 25.55 2.245 ;
 RECT 25.45 2.245 25.735 2.455 ;
 RECT 22.615 1.01 22.85 1.22 ;
 RECT 22.75 1.22 22.85 1.81 ;
 RECT 15.46 1.635 15.56 1.66 ;
 RECT 15.46 1.66 15.715 1.87 ;
 RECT 15.46 1.87 15.56 2.565 ;
 RECT 21.515 1.075 21.8 1.305 ;
 LAYER CO ;
 RECT 22.025 1.4 22.155 1.53 ;
 RECT 17.79 0.975 17.92 1.105 ;
 RECT 4.275 2.115 4.405 2.245 ;
 RECT 5.4 1.495 5.53 1.625 ;
 RECT 0.39 2.345 0.52 2.475 ;
 RECT 3.745 2.05 3.875 2.18 ;
 RECT 12.905 0.595 13.035 0.725 ;
 RECT 12.4 1.9 12.53 2.03 ;
 RECT 16.115 0.83 16.245 0.96 ;
 RECT 6.835 2 6.965 2.13 ;
 RECT 5.35 0.97 5.48 1.1 ;
 RECT 3.745 0.775 3.875 0.905 ;
 RECT 14.835 1.705 14.965 1.835 ;
 RECT 14.835 0.96 14.965 1.09 ;
 RECT 0.895 0.775 1.025 0.905 ;
 RECT 9.145 2.015 9.275 2.145 ;
 RECT 3.745 1.79 3.875 1.92 ;
 RECT 9.63 0.88 9.76 1.01 ;
 RECT 17.275 0.305 17.405 0.435 ;
 RECT 6.81 0.525 6.94 0.655 ;
 RECT 7.275 1.345 7.405 1.475 ;
 RECT 8.135 0.455 8.265 0.585 ;
 RECT 5.115 0.21 5.245 0.34 ;
 RECT 25.67 0.59 25.8 0.72 ;
 RECT 12.905 1.87 13.035 2 ;
 RECT 1.37 1.55 1.5 1.68 ;
 RECT 2.505 2.115 2.635 2.245 ;
 RECT 6.925 0.88 7.055 1.01 ;
 RECT 10.075 1.885 10.205 2.015 ;
 RECT 2.49 1.23 2.62 1.36 ;
 RECT 5.485 2.345 5.615 2.475 ;
 RECT 11.14 1.28 11.27 1.41 ;
 RECT 16.115 1.78 16.245 1.91 ;
 RECT 11.875 0.875 12.005 1.005 ;
 RECT 2.9 0.225 3.03 0.355 ;
 RECT 15.215 0.33 15.345 0.46 ;
 RECT 25.67 1.44 25.8 1.57 ;
 RECT 18.785 2.64 18.915 2.77 ;
 RECT 5.22 1.995 5.35 2.125 ;
 RECT 0.39 1.825 0.52 1.955 ;
 RECT 17.27 2.64 17.4 2.77 ;
 RECT 0.895 2.055 1.025 2.185 ;
 RECT 4.345 0.325 4.475 0.455 ;
 RECT 9.63 2.07 9.76 2.2 ;
 RECT 7.31 2.04 7.44 2.17 ;
 RECT 16.785 0.975 16.915 1.105 ;
 RECT 15.21 2.64 15.34 2.77 ;
 RECT 1.97 1.195 2.1 1.325 ;
 RECT 10.965 0.62 11.095 0.75 ;
 RECT 24.725 1.465 24.855 1.595 ;
 RECT 4.865 1.55 4.995 1.68 ;
 RECT 14.365 2.64 14.495 2.77 ;
 RECT 1.365 2.315 1.495 2.445 ;
 RECT 11.875 1.945 12.005 2.075 ;
 RECT 0.355 0.59 0.485 0.72 ;
 RECT 24.89 0.115 25.02 0.245 ;
 RECT 9.145 0.93 9.275 1.06 ;
 RECT 8.675 2.135 8.805 2.265 ;
 RECT 19.37 1.71 19.5 1.84 ;
 RECT 8.205 2.03 8.335 2.16 ;
 RECT 1.365 0.775 1.495 0.905 ;
 RECT 12.4 0.595 12.53 0.725 ;
 RECT 4.745 2.05 4.875 2.18 ;
 RECT 24.355 1.38 24.485 1.51 ;
 RECT 5.995 1.825 6.125 1.955 ;
 RECT 4.745 0.13 4.875 0.26 ;
 RECT 6.365 2.035 6.495 2.165 ;
 RECT 4.275 0.79 4.405 0.92 ;
 RECT 6.455 0.88 6.585 1.01 ;
 RECT 2.67 1.64 2.8 1.77 ;
 RECT 19.37 0.78 19.5 0.91 ;
 RECT 18.31 0.77 18.44 0.9 ;
 RECT 18.31 1.725 18.44 1.855 ;
 RECT 6.06 0.905 6.19 1.035 ;
 RECT 21.775 0.505 21.905 0.635 ;
 RECT 8.815 1.63 8.945 1.76 ;
 RECT 3.385 1.195 3.515 1.325 ;
 RECT 0.39 2.085 0.52 2.215 ;
 RECT 18.59 1.25 18.72 1.38 ;
 RECT 16.785 1.72 16.915 1.85 ;
 RECT 17.79 1.72 17.92 1.85 ;
 RECT 3.275 2.09 3.405 2.22 ;
 RECT 26.315 1.45 26.445 1.58 ;
 RECT 23.275 0.41 23.405 0.54 ;
 RECT 3.275 0.585 3.405 0.715 ;
 RECT 11.135 2.295 11.265 2.425 ;
 RECT 7.815 2.29 7.945 2.42 ;
 RECT 6.17 1.5 6.3 1.63 ;
 RECT 23.71 0.11 23.84 0.24 ;
 RECT 21.36 0.61 21.49 0.74 ;
 RECT 13.49 1.445 13.62 1.575 ;
 RECT 8.95 0.54 9.08 0.67 ;
 RECT 16.09 0.265 16.22 0.395 ;
 RECT 14.46 1.3 14.59 1.43 ;
 RECT 13.14 2.37 13.27 2.5 ;
 RECT 21.62 1.135 21.75 1.265 ;
 RECT 15.785 1.29 15.915 1.42 ;
 RECT 25.52 1.05 25.65 1.18 ;
 RECT 9.96 1.45 10.09 1.58 ;
 RECT 23.115 1.01 23.245 1.14 ;
 RECT 23.625 1.025 23.755 1.155 ;
 RECT 16.46 0.67 16.59 0.8 ;
 RECT 25.555 2.285 25.685 2.415 ;
 RECT 24.52 0.295 24.65 0.425 ;
 RECT 22.665 1.05 22.795 1.18 ;
 RECT 15.535 1.7 15.665 1.83 ;
 RECT 20.635 0.265 20.765 0.395 ;
 RECT 19.85 2.64 19.98 2.77 ;
 RECT 20.35 0.78 20.48 0.91 ;
 RECT 20.35 1.71 20.48 1.84 ;
 RECT 19.87 0.78 20 0.91 ;
 RECT 0.355 0.33 0.485 0.46 ;
 RECT 24.19 0.59 24.32 0.72 ;
 RECT 22.495 0.11 22.625 0.24 ;
 RECT 1.365 2.055 1.495 2.185 ;
 RECT 18.87 0.77 19 0.9 ;
 RECT 14.14 0.955 14.27 1.085 ;
 RECT 23.88 1.42 24.01 1.55 ;
 RECT 22.495 1.45 22.625 1.58 ;
 RECT 10.775 2.445 10.905 2.575 ;
 RECT 23.275 1.46 23.405 1.59 ;
 RECT 3.275 2.35 3.405 2.48 ;
 RECT 10.075 0.88 10.205 1.01 ;
 RECT 2.31 0.775 2.44 0.905 ;
 LAYER M1 ;
 RECT 12.9 0.965 13.96 1.105 ;
 RECT 14.415 0.665 16.25 0.805 ;
 RECT 16.11 0.22 16.25 0.225 ;
 RECT 16.11 0.435 16.25 0.665 ;
 RECT 16.11 0.805 16.25 1.98 ;
 RECT 16.04 0.225 16.27 0.435 ;
 RECT 14.83 1.37 15.965 1.46 ;
 RECT 14.83 1.095 14.97 1.37 ;
 RECT 14.83 1.46 15.96 1.51 ;
 RECT 14.83 1.51 14.97 1.7 ;
 RECT 15.735 1.25 15.965 1.37 ;
 RECT 14.765 1.7 15.04 1.84 ;
 RECT 14.76 0.955 15.03 1.095 ;
 RECT 9.91 1.41 10.21 1.46 ;
 RECT 9.91 1.6 10.21 1.62 ;
 RECT 10.07 0.81 10.21 1.41 ;
 RECT 10.07 1.62 10.21 2.085 ;
 RECT 10.82 1.415 10.96 1.46 ;
 RECT 9.91 1.46 10.96 1.6 ;
 RECT 10.82 1.275 11.34 1.415 ;
 RECT 23.575 1.195 23.715 1.32 ;
 RECT 23.27 1.46 23.41 1.735 ;
 RECT 23.59 0.705 23.73 0.985 ;
 RECT 23.27 0.33 23.41 0.565 ;
 RECT 23.27 1.32 23.715 1.46 ;
 RECT 23.27 0.565 23.73 0.705 ;
 RECT 23.575 0.985 23.805 1.195 ;
 RECT 16.41 0.72 16.64 0.84 ;
 RECT 17.68 0.37 17.82 0.58 ;
 RECT 16.41 0.63 17.82 0.72 ;
 RECT 16.42 0.58 17.82 0.63 ;
 RECT 18.585 0.37 18.725 1.46 ;
 RECT 17.68 0.23 18.725 0.37 ;
 RECT 13.09 2.42 13.32 2.54 ;
 RECT 25.505 2.245 25.735 2.28 ;
 RECT 25.505 2.42 25.735 2.455 ;
 RECT 13.09 2.28 25.735 2.42 ;
 RECT 24.56 0.465 24.7 0.685 ;
 RECT 24.47 0.255 24.7 0.465 ;
 RECT 24.56 0.685 25.985 0.825 ;
 RECT 25.845 0.825 25.985 1.36 ;
 RECT 25.665 1.5 25.805 1.705 ;
 RECT 25.665 0.485 25.805 0.685 ;
 RECT 25.665 1.36 25.985 1.5 ;
 RECT 21.845 0.64 21.985 1.03 ;
 RECT 22.02 1.17 22.16 1.6 ;
 RECT 21.57 1.17 21.8 1.305 ;
 RECT 21.725 0.5 21.985 0.64 ;
 RECT 22.615 1.01 22.845 1.03 ;
 RECT 22.615 1.17 22.845 1.22 ;
 RECT 21.565 1.03 22.845 1.17 ;
 RECT 20.585 0.36 20.815 0.435 ;
 RECT 22.125 0.36 22.265 0.54 ;
 RECT 20.585 0.22 22.265 0.36 ;
 RECT 22.99 0.97 23.295 1.18 ;
 RECT 22.99 0.68 23.13 0.97 ;
 RECT 22.125 0.54 23.13 0.68 ;
 RECT 22.99 0.535 23.13 0.54 ;
 RECT 0.89 0.72 1.03 1.195 ;
 RECT 0.89 1.335 1.03 2.27 ;
 RECT 1.675 0.36 1.815 1.195 ;
 RECT 0.89 1.195 1.815 1.335 ;
 RECT 1.675 0.22 3.1 0.36 ;
 RECT 5.26 1.63 5.4 1.99 ;
 RECT 5.26 1.475 5.605 1.63 ;
 RECT 5.345 0.9 5.485 1.475 ;
 RECT 5.15 1.99 5.4 2.13 ;
 RECT 13.435 1.43 13.67 1.615 ;
 RECT 13.435 1.615 13.575 1.985 ;
 RECT 13.44 1.405 13.67 1.43 ;
 RECT 13.435 1.985 15.67 2.125 ;
 RECT 15.485 1.87 15.67 1.985 ;
 RECT 15.485 1.66 15.715 1.87 ;
 RECT 24.185 0.48 24.325 1.08 ;
 RECT 24.35 1.22 24.49 1.58 ;
 RECT 25.47 1.01 25.7 1.08 ;
 RECT 24.185 1.08 25.7 1.22 ;
 RECT 6.92 0.805 7.06 1.69 ;
 RECT 6.92 1.83 7.06 1.935 ;
 RECT 6.83 1.935 7.06 2.2 ;
 RECT 6.92 1.69 9 1.83 ;
 RECT 8.76 1.58 9 1.69 ;
 RECT 8.76 1.83 9 1.835 ;
 RECT 4.05 0.925 4.19 1.195 ;
 RECT 4.05 1.335 4.19 2.11 ;
 RECT 4.05 0.785 4.475 0.925 ;
 RECT 4.05 2.11 4.475 2.25 ;
 RECT 4.745 0.75 4.885 1.195 ;
 RECT 4.05 1.195 4.885 1.335 ;
 RECT 4.745 0.61 5.56 0.75 ;
 RECT 5.42 0.22 6.59 0.36 ;
 RECT 6.45 0.36 6.59 0.9 ;
 RECT 6.525 1.08 6.665 1.945 ;
 RECT 5.42 0.36 5.56 0.61 ;
 RECT 6.36 2.17 6.5 2.305 ;
 RECT 6.36 1.945 6.665 2.17 ;
 RECT 6.45 0.9 6.665 1.08 ;
 RECT 6.74 0.52 7.34 0.66 ;
 RECT 7.2 0.66 7.34 1.015 ;
 RECT 8.745 0.505 9.13 0.71 ;
 RECT 7.2 1.015 8.885 1.155 ;
 RECT 8.9 0.5 9.13 0.505 ;
 RECT 8.745 0.71 8.885 1.015 ;
 RECT 3.74 0.57 3.88 2.25 ;
 RECT 4.235 0.22 4.6 0.43 ;
 RECT 4.235 0.57 4.6 0.615 ;
 RECT 3.74 0.43 4.6 0.57 ;
 RECT 10.475 1.88 10.615 2.225 ;
 RECT 9.625 0.82 9.765 2.225 ;
 RECT 9.625 2.225 10.615 2.365 ;
 RECT 10.475 1.755 12.545 1.88 ;
 RECT 10.485 1.74 12.545 1.755 ;
 RECT 11.87 0.765 12.01 1.74 ;
 RECT 11.87 1.88 12.01 2.165 ;
 RECT 12.395 0.525 12.535 1.74 ;
 RECT 12.395 1.88 12.535 2.155 ;
 RECT 7.2 1.44 7.465 1.55 ;
 RECT 9.14 0.865 9.28 1.3 ;
 RECT 9.14 1.44 9.28 2.215 ;
 RECT 7.2 1.3 9.28 1.44 ;
 RECT 6.055 1.67 6.195 1.82 ;
 RECT 6.055 1.96 6.195 2.455 ;
 RECT 7.765 2.25 7.995 2.455 ;
 RECT 6.055 0.805 6.195 1.46 ;
 RECT 6.055 1.46 6.35 1.67 ;
 RECT 5.925 1.82 6.195 1.96 ;
 RECT 6.055 2.455 7.995 2.595 ;
 RECT 2.96 0.91 3.1 1.19 ;
 RECT 2.96 1.33 3.1 2.11 ;
 RECT 2.255 0.77 3.1 0.91 ;
 RECT 2.45 2.11 3.1 2.25 ;
 RECT 3.38 1.145 3.52 1.19 ;
 RECT 3.38 1.33 3.52 1.375 ;
 RECT 2.96 1.19 3.52 1.33 ;
 RECT 8.2 2.11 8.34 2.23 ;
 RECT 7.305 2.11 7.445 2.24 ;
 RECT 7.305 1.97 8.34 2.11 ;
 RECT 14.415 0.805 14.555 1.26 ;
 RECT 14.41 1.26 14.64 1.295 ;
 RECT 14.41 1.435 14.64 1.47 ;
 RECT 13.82 1.295 14.64 1.435 ;
 RECT 13.82 1.105 13.96 1.295 ;
 RECT 12.9 0.525 13.04 0.965 ;
 RECT 12.9 1.105 13.04 2.065 ;
 END
END RSDFFSRX2

MACRO MUX21X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN S
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.95 1.475 1.475 1.75 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END S

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 1.13 1.985 1.27 2.8 ;
 RECT 3.04 2.04 3.18 2.8 ;
 RECT 0.24 1.545 0.38 2.8 ;
 RECT 3.98 1.545 4.12 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.735 1.14 1.875 1.475 ;
 RECT 1.64 1.63 2.585 1.79 ;
 RECT 1.64 1.475 1.88 1.63 ;
 RECT 2.435 1.79 2.575 1.845 ;
 RECT 2.435 1.57 2.575 1.63 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 3.04 0.08 3.18 0.78 ;
 RECT 3.98 0.08 4.12 0.78 ;
 RECT 0.24 0.08 0.38 0.88 ;
 RECT 1.13 0.08 1.27 0.97 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.51 1.415 3.65 2.25 ;
 RECT 3.51 1.15 3.8 1.415 ;
 RECT 3.51 0.715 3.65 1.15 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END Q

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.1 1.155 2.485 1.415 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 2.105 1.41 2.205 1.645 ;
 RECT 2.335 0.555 2.435 1.18 ;
 RECT 2.055 1.745 2.155 2.735 ;
 RECT 2.055 1.645 2.205 1.745 ;
 RECT 2.105 1.18 2.435 1.41 ;
 RECT 3.15 1.08 3.395 1.15 ;
 RECT 3.15 1.15 3.865 1.25 ;
 RECT 3.15 1.25 3.395 1.29 ;
 RECT 3.765 0.335 3.865 1.15 ;
 RECT 3.765 1.25 3.865 2.745 ;
 RECT 3.295 0.335 3.395 1.08 ;
 RECT 3.295 1.29 3.395 2.745 ;
 RECT 2.525 1.82 2.625 2.735 ;
 RECT 2.385 1.59 2.625 1.82 ;
 RECT 2.825 0.515 2.925 2.735 ;
 RECT 2.62 0.285 2.925 0.515 ;
 RECT 1.72 0.555 1.82 1.145 ;
 RECT 1.68 1.145 1.925 1.385 ;
 RECT 0.915 1.475 1.485 1.75 ;
 RECT 0.915 0.555 1.015 1.475 ;
 RECT 0.915 1.75 1.015 2.685 ;
 RECT 1.385 0.555 1.485 1.475 ;
 RECT 1.385 1.75 1.485 2.735 ;
 LAYER CO ;
 RECT 1.135 2.315 1.265 2.445 ;
 RECT 3.985 1.595 4.115 1.725 ;
 RECT 3.985 1.855 4.115 1.985 ;
 RECT 3.985 2.115 4.115 2.245 ;
 RECT 3.515 1.53 3.645 1.66 ;
 RECT 3.045 2.09 3.175 2.22 ;
 RECT 3.985 0.585 4.115 0.715 ;
 RECT 3.985 2.375 4.115 2.505 ;
 RECT 0.665 2.055 0.795 2.185 ;
 RECT 1.135 0.775 1.265 0.905 ;
 RECT 0.245 0.43 0.375 0.56 ;
 RECT 0.245 0.69 0.375 0.82 ;
 RECT 3.515 2.05 3.645 2.18 ;
 RECT 0.665 0.775 0.795 0.905 ;
 RECT 2.26 1.23 2.39 1.36 ;
 RECT 2.08 0.775 2.21 0.905 ;
 RECT 3.045 0.585 3.175 0.715 ;
 RECT 2.44 1.64 2.57 1.77 ;
 RECT 1.14 1.55 1.27 1.68 ;
 RECT 3.045 2.35 3.175 2.48 ;
 RECT 0.245 2.12 0.375 2.25 ;
 RECT 1.74 1.195 1.87 1.325 ;
 RECT 3.2 1.12 3.33 1.25 ;
 RECT 1.135 2.055 1.265 2.185 ;
 RECT 3.515 1.79 3.645 1.92 ;
 RECT 2.275 2.115 2.405 2.245 ;
 RECT 2.67 0.335 2.8 0.465 ;
 RECT 3.515 0.775 3.645 0.905 ;
 RECT 0.245 1.6 0.375 1.73 ;
 RECT 0.245 1.86 0.375 1.99 ;
 LAYER M1 ;
 RECT 2.73 0.91 2.87 1.115 ;
 RECT 2.73 1.255 2.87 2.11 ;
 RECT 2.025 0.77 2.87 0.91 ;
 RECT 2.22 2.11 2.87 2.25 ;
 RECT 2.73 1.115 3.35 1.255 ;
 RECT 3.195 1.07 3.335 1.115 ;
 RECT 3.195 1.255 3.335 1.3 ;
 RECT 0.66 0.72 0.8 1.195 ;
 RECT 0.66 1.335 0.8 2.305 ;
 RECT 1.445 0.47 1.585 1.195 ;
 RECT 0.66 1.195 1.585 1.335 ;
 RECT 1.445 0.33 2.87 0.47 ;
 END
END MUX21X2

MACRO MUX41X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8 2.96 ;
 RECT 3.57 2.335 3.71 2.8 ;
 RECT 7.275 1.71 7.415 2.8 ;
 RECT 0.195 1.545 0.335 2.8 ;
 RECT 5.51 1.71 5.65 2.8 ;
 RECT 1.065 1.795 1.205 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.8 2.25 6.08 2.55 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.745 2.245 7.135 2.515 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END IN1

 PIN S1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.555 2.115 7.82 2.43 ;
 END
 ANTENNAGATEAREA 0.233 ;
 END S1

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.755 1.205 4.13 1.6 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END IN4

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8 0.08 ;
 RECT 5.51 0.08 5.65 0.805 ;
 RECT 7.275 0.08 7.415 0.805 ;
 RECT 1.065 0.08 1.205 0.775 ;
 RECT 3.58 0.08 3.72 0.785 ;
 RECT 0.195 0.08 0.335 0.88 ;
 END
 END VSS

 PIN S0
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.98 1.155 1.43 1.295 ;
 RECT 0.98 1.295 1.33 1.4 ;
 END
 ANTENNAGATEAREA 0.118 ;
 END S0

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.36 1.14 0.735 1.4 ;
 RECT 0.595 1.4 0.735 2.225 ;
 RECT 0.595 0.735 0.735 1.14 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END Q

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.985 2.255 5.365 2.54 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END IN3

 OBS
 LAYER PO ;
 RECT 7.53 2.21 7.785 2.43 ;
 RECT 4.605 1.25 4.705 2.395 ;
 RECT 4.145 0.22 4.245 1.15 ;
 RECT 6.645 1.43 6.745 2.69 ;
 RECT 6.175 0.22 6.275 0.97 ;
 RECT 4.145 0.12 7.63 0.22 ;
 RECT 7.53 2.43 7.63 2.69 ;
 RECT 7.53 0.22 7.63 2.21 ;
 RECT 4.145 1.15 4.705 1.25 ;
 RECT 6.645 2.69 7.63 2.79 ;
 RECT 5.765 0.4 5.865 2.295 ;
 RECT 5.765 2.295 5.995 2.505 ;
 RECT 4.615 0.9 5.105 0.97 ;
 RECT 4.615 0.4 4.715 0.87 ;
 RECT 4.615 0.87 5.095 0.9 ;
 RECT 4.895 0.97 5.105 1.13 ;
 RECT 0.85 0.35 0.95 2.645 ;
 RECT 1.855 2.34 1.955 2.645 ;
 RECT 0.85 2.645 1.955 2.745 ;
 RECT 1.79 2.13 2.02 2.34 ;
 RECT 6.645 0.4 6.745 1.035 ;
 RECT 4.135 1.43 4.235 2.685 ;
 RECT 6.175 1.25 6.275 2.685 ;
 RECT 6.175 1.15 6.875 1.245 ;
 RECT 6.645 1.035 6.875 1.15 ;
 RECT 6.175 1.245 6.745 1.25 ;
 RECT 4.135 2.685 6.275 2.785 ;
 RECT 6.95 1.53 7.05 2.28 ;
 RECT 7.06 0.4 7.16 1.43 ;
 RECT 6.95 1.43 7.16 1.53 ;
 RECT 6.93 2.28 7.19 2.51 ;
 RECT 1.32 0.57 1.42 1.11 ;
 RECT 1.32 1.34 1.42 1.835 ;
 RECT 1.21 1.15 2.96 1.25 ;
 RECT 1.21 1.11 1.42 1.15 ;
 RECT 1.21 1.25 1.42 1.34 ;
 RECT 2.86 0.4 2.96 1.15 ;
 RECT 2.39 1.25 2.49 2.395 ;
 RECT 5.295 0.4 5.395 2.295 ;
 RECT 5.17 2.295 5.4 2.505 ;
 RECT 3.835 0.385 3.935 1.26 ;
 RECT 3.835 1.47 3.935 2.395 ;
 RECT 3.71 1.26 3.94 1.47 ;
 RECT 2.39 0.43 2.49 0.97 ;
 RECT 2.39 0.22 2.6 0.43 ;
 RECT 2.86 1.435 2.96 2.295 ;
 RECT 2.86 2.295 3.455 2.395 ;
 RECT 3.355 0.22 3.455 2.295 ;
 RECT 2.39 0.12 3.455 0.22 ;
 LAYER CO ;
 RECT 0.6 1.515 0.73 1.645 ;
 RECT 0.2 2.12 0.33 2.25 ;
 RECT 3.575 2.385 3.705 2.515 ;
 RECT 3.08 1.715 3.21 1.845 ;
 RECT 7.28 2.03 7.41 2.16 ;
 RECT 3.76 1.3 3.89 1.43 ;
 RECT 3.585 0.605 3.715 0.735 ;
 RECT 2.43 0.25 2.56 0.38 ;
 RECT 5.515 2.03 5.645 2.16 ;
 RECT 1.54 1.485 1.67 1.615 ;
 RECT 1.635 0.79 1.765 0.92 ;
 RECT 7.28 0.62 7.41 0.75 ;
 RECT 7.6 2.25 7.73 2.38 ;
 RECT 5.815 2.335 5.945 2.465 ;
 RECT 6.395 0.62 6.525 0.75 ;
 RECT 2.14 0.62 2.27 0.75 ;
 RECT 6.395 1.715 6.525 1.845 ;
 RECT 4.365 0.62 4.495 0.75 ;
 RECT 4.355 1.715 4.485 1.845 ;
 RECT 7.75 0.62 7.88 0.75 ;
 RECT 4.935 0.95 5.065 1.08 ;
 RECT 2.14 1.705 2.27 1.835 ;
 RECT 2.61 0.62 2.74 0.75 ;
 RECT 7.75 1.695 7.88 1.825 ;
 RECT 0.6 0.79 0.73 0.92 ;
 RECT 3.08 0.62 3.21 0.75 ;
 RECT 0.6 2.035 0.73 2.165 ;
 RECT 4.355 1.975 4.485 2.105 ;
 RECT 7.28 1.77 7.41 1.9 ;
 RECT 6.395 1.975 6.525 2.105 ;
 RECT 5.515 1.77 5.645 1.9 ;
 RECT 1.07 1.85 1.2 1.98 ;
 RECT 1.07 2.11 1.2 2.24 ;
 RECT 0.6 1.775 0.73 1.905 ;
 RECT 2.61 1.715 2.74 1.845 ;
 RECT 1.07 2.37 1.2 2.5 ;
 RECT 1.84 2.17 1.97 2.3 ;
 RECT 0.2 1.6 0.33 1.73 ;
 RECT 0.2 0.43 0.33 0.56 ;
 RECT 6.695 1.075 6.825 1.205 ;
 RECT 6.975 2.33 7.105 2.46 ;
 RECT 0.2 1.86 0.33 1.99 ;
 RECT 1.07 0.59 1.2 0.72 ;
 RECT 1.25 1.16 1.38 1.29 ;
 RECT 0.2 0.69 0.33 0.82 ;
 RECT 5.515 0.62 5.645 0.75 ;
 RECT 5.22 2.335 5.35 2.465 ;
 LAYER M1 ;
 RECT 3.075 0.56 3.215 0.925 ;
 RECT 3.075 1.065 3.215 1.895 ;
 RECT 3.075 0.925 4.5 1.065 ;
 RECT 4.36 0.57 4.5 0.925 ;
 RECT 4.35 1.065 4.49 2.16 ;
 RECT 1.63 0.385 1.77 1.48 ;
 RECT 1.63 0.245 2.61 0.385 ;
 RECT 1.48 1.48 1.77 1.62 ;
 RECT 4.705 1.365 4.845 2.35 ;
 RECT 3.965 2.35 4.845 2.49 ;
 RECT 3.355 1.905 4.105 2.035 ;
 RECT 3.965 2.045 4.105 2.35 ;
 RECT 2.925 2.035 4.105 2.045 ;
 RECT 2.925 2.175 3.065 2.5 ;
 RECT 1.485 2.5 3.065 2.64 ;
 RECT 2.135 0.56 2.275 1.76 ;
 RECT 2.925 2.045 3.495 2.175 ;
 RECT 1.485 1.9 1.625 2.5 ;
 RECT 1.485 1.76 2.275 1.9 ;
 RECT 6.39 0.56 6.53 1.225 ;
 RECT 6.39 1.365 6.53 2.17 ;
 RECT 4.705 1.225 6.53 1.365 ;
 RECT 2.605 0.56 2.745 2.05 ;
 RECT 1.835 2.19 1.975 2.35 ;
 RECT 1.835 2.05 2.745 2.19 ;
 RECT 5.79 0.41 5.93 0.945 ;
 RECT 6.69 1.205 6.83 1.255 ;
 RECT 4.885 0.945 5.93 1.085 ;
 RECT 5.79 0.27 6.83 0.41 ;
 RECT 6.69 0.41 6.83 1.065 ;
 RECT 7.745 0.565 7.885 1.065 ;
 RECT 7.745 1.205 7.885 1.895 ;
 RECT 6.69 1.065 7.885 1.205 ;
 END
END MUX41X1

MACRO SHFILL1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 0.32 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 0.32 2.96 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 0.32 0.08 ;
 END
 END VSS

END SHFILL1

MACRO SHFILL128
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 40.96 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 40.96 0.08 ;
 RECT 0.41 0.08 0.55 0.79 ;
 RECT 40.405 0.08 40.545 0.785 ;
 RECT 30.485 0.08 30.625 0.785 ;
 RECT 20.565 0.08 20.705 0.785 ;
 RECT 10.645 0.08 10.785 0.785 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 40.96 2.96 ;
 RECT 0.41 2.095 0.55 2.8 ;
 RECT 40.405 2.09 40.545 2.8 ;
 RECT 30.485 2.09 30.625 2.8 ;
 RECT 20.565 2.09 20.705 2.8 ;
 RECT 10.645 2.09 10.785 2.8 ;
 END
 END VDD

 OBS
 LAYER CO ;
 RECT 10.65 2.16 10.78 2.29 ;
 RECT 10.65 0.325 10.78 0.455 ;
 RECT 10.65 2.44 10.78 2.57 ;
 RECT 10.65 0.605 10.78 0.735 ;
 RECT 20.57 2.44 20.7 2.57 ;
 RECT 20.57 2.16 20.7 2.29 ;
 RECT 20.57 0.325 20.7 0.455 ;
 RECT 20.57 0.605 20.7 0.735 ;
 RECT 30.49 2.44 30.62 2.57 ;
 RECT 30.49 2.16 30.62 2.29 ;
 RECT 30.49 0.325 30.62 0.455 ;
 RECT 30.49 0.605 30.62 0.735 ;
 RECT 40.41 0.325 40.54 0.455 ;
 RECT 40.41 0.605 40.54 0.735 ;
 RECT 40.41 2.44 40.54 2.57 ;
 RECT 40.41 2.16 40.54 2.29 ;
 RECT 0.415 2.165 0.545 2.295 ;
 RECT 0.415 0.325 0.545 0.455 ;
 RECT 0.415 2.445 0.545 2.575 ;
 RECT 0.415 0.605 0.545 0.735 ;
 END
END SHFILL128

MACRO SHFILL2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 0.64 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 0.64 2.96 ;
 RECT 0.265 2.095 0.405 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 0.64 0.08 ;
 RECT 0.265 0.08 0.405 0.79 ;
 END
 END VSS

 OBS
 LAYER CO ;
 RECT 0.27 0.305 0.4 0.435 ;
 RECT 0.27 0.585 0.4 0.715 ;
 RECT 0.27 2.165 0.4 2.295 ;
 RECT 0.27 2.445 0.4 2.575 ;
 END
END SHFILL2

MACRO SHFILL3
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 0.96 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 0.96 2.96 ;
 RECT 0.41 2.095 0.55 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 0.96 0.08 ;
 RECT 0.41 0.08 0.55 0.79 ;
 END
 END VSS

 OBS
 LAYER CO ;
 RECT 0.415 2.165 0.545 2.295 ;
 RECT 0.415 0.305 0.545 0.435 ;
 RECT 0.415 2.445 0.545 2.575 ;
 RECT 0.415 0.585 0.545 0.715 ;
 END
END SHFILL3

MACRO SHFILL64
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 20.48 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 20.48 0.08 ;
 RECT 10.645 0.08 10.785 0.785 ;
 RECT 19.935 0.08 20.075 0.785 ;
 RECT 0.41 0.08 0.55 0.79 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 20.48 2.96 ;
 RECT 10.645 2.09 10.785 2.8 ;
 RECT 19.935 2.09 20.075 2.8 ;
 RECT 0.41 2.095 0.55 2.8 ;
 END
 END VDD

 OBS
 LAYER CO ;
 RECT 0.415 0.605 0.545 0.735 ;
 RECT 0.415 2.445 0.545 2.575 ;
 RECT 0.415 0.325 0.545 0.455 ;
 RECT 0.415 2.165 0.545 2.295 ;
 RECT 19.94 0.6 20.07 0.73 ;
 RECT 19.94 0.32 20.07 0.45 ;
 RECT 19.94 2.16 20.07 2.29 ;
 RECT 19.94 2.44 20.07 2.57 ;
 RECT 10.65 0.6 10.78 0.73 ;
 RECT 10.65 2.44 10.78 2.57 ;
 RECT 10.65 0.32 10.78 0.45 ;
 RECT 10.65 2.16 10.78 2.29 ;
 END
END SHFILL64

MACRO TIEH
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 1.6 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 1.6 0.08 ;
 RECT 0.73 0.08 0.87 0.92 ;
 RECT 0.27 0.08 0.41 0.76 ;
 END
 END VSS

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.13 2.095 1.43 2.39 ;
 RECT 1.2 2.39 1.34 2.535 ;
 RECT 1.2 1.475 1.34 2.095 ;
 END
 ANTENNADIFFAREA 0.325 ;
 END Z

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0.65 2.25 0.95 2.545 ;
 RECT 0.73 1.475 0.87 2.25 ;
 RECT 0 2.8 1.6 2.96 ;
 RECT 0.73 2.545 0.87 2.8 ;
 RECT 0.315 1.5 0.455 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.985 0.22 1.085 2.74 ;
 RECT 0.935 1.08 1.165 1.29 ;
 LAYER CO ;
 RECT 0.32 1.55 0.45 1.68 ;
 RECT 0.32 1.81 0.45 1.94 ;
 RECT 0.275 0.58 0.405 0.71 ;
 RECT 0.275 0.32 0.405 0.45 ;
 RECT 0.32 2.07 0.45 2.2 ;
 RECT 1.205 2.355 1.335 2.485 ;
 RECT 1.205 1.525 1.335 1.655 ;
 RECT 1.205 2.095 1.335 2.225 ;
 RECT 1.205 1.785 1.335 1.915 ;
 RECT 1.205 0.515 1.335 0.645 ;
 RECT 1.205 0.775 1.335 0.905 ;
 RECT 0.735 0.48 0.865 0.61 ;
 RECT 0.735 0.74 0.865 0.87 ;
 RECT 0.735 2.355 0.865 2.485 ;
 RECT 0.735 1.525 0.865 1.655 ;
 RECT 0.735 1.785 0.865 1.915 ;
 RECT 0.735 2.095 0.865 2.225 ;
 RECT 0.985 1.12 1.115 1.25 ;
 LAYER M1 ;
 RECT 1.2 0.44 1.34 1.255 ;
 RECT 0.98 1.115 1.34 1.255 ;
 RECT 0.935 1.08 1.34 1.255 ;
 RECT 0.935 1.08 1.165 1.29 ;
 END
END TIEH

MACRO TIEL
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 1.6 BY 2.88 ;
 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.13 0.47 1.43 0.79 ;
 RECT 1.2 0.79 1.34 0.92 ;
 END
 ANTENNADIFFAREA 0.162 ;
 END ZN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0.65 0.645 0.95 0.94 ;
 RECT 0 -0.08 1.6 0.08 ;
 RECT 0.73 0.08 0.87 0.645 ;
 RECT 0.27 0.08 0.41 0.76 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 1.6 2.96 ;
 RECT 0.73 1.475 0.87 2.8 ;
 RECT 0.315 1.5 0.455 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.985 0.22 1.085 2.74 ;
 RECT 0.935 1.08 1.165 1.29 ;
 LAYER CO ;
 RECT 1.205 0.74 1.335 0.87 ;
 RECT 1.205 0.48 1.335 0.61 ;
 RECT 0.735 0.74 0.865 0.87 ;
 RECT 1.205 2.355 1.335 2.485 ;
 RECT 0.735 0.48 0.865 0.61 ;
 RECT 0.735 2.355 0.865 2.485 ;
 RECT 0.32 1.55 0.45 1.68 ;
 RECT 0.275 0.32 0.405 0.45 ;
 RECT 0.275 0.58 0.405 0.71 ;
 RECT 0.32 1.81 0.45 1.94 ;
 RECT 0.735 1.525 0.865 1.655 ;
 RECT 1.205 2.095 1.335 2.225 ;
 RECT 0.735 2.095 0.865 2.225 ;
 RECT 1.205 1.525 1.335 1.655 ;
 RECT 0.32 2.07 0.45 2.2 ;
 RECT 1.205 1.785 1.335 1.915 ;
 RECT 0.735 1.785 0.865 1.915 ;
 RECT 0.985 1.12 1.115 1.25 ;
 LAYER M1 ;
 RECT 1.2 1.11 1.34 2.535 ;
 RECT 0.98 1.115 1.34 1.255 ;
 RECT 0.935 1.08 1.34 1.29 ;
 RECT 0.935 1.115 1.34 1.29 ;
 RECT 0.935 1.08 1.165 1.29 ;
 END
END TIEL

MACRO DEC24X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.24 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.27 2.11 5.56 2.365 ;
 END
 ANTENNAGATEAREA 0.174 ;
 END IN2

 PIN Q2
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.03 1.48 4.34 1.795 ;
 RECT 4.145 0.71 4.285 1.48 ;
 END
 ANTENNADIFFAREA 0.502 ;
 END Q2

 PIN Q3
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.105 1.8 1.4 2.05 ;
 RECT 1.105 0.775 1.5 0.915 ;
 RECT 1.105 2.05 1.245 2.62 ;
 RECT 1.105 0.915 1.245 1.8 ;
 END
 ANTENNADIFFAREA 0.441 ;
 END Q3

 PIN Q1
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.545 0.775 10.04 0.915 ;
 RECT 9.77 0.52 10.04 0.775 ;
 RECT 9.62 0.915 9.76 1.575 ;
 RECT 9.615 1.73 9.755 2.62 ;
 RECT 9.615 1.575 9.76 1.73 ;
 END
 ANTENNADIFFAREA 0.502 ;
 END Q1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.24 2.96 ;
 RECT 6.985 2.435 7.255 2.575 ;
 RECT 9.125 1.865 9.265 2.8 ;
 RECT 8.01 1.865 8.15 2.8 ;
 RECT 1.575 1.865 1.715 2.8 ;
 RECT 3.65 2.555 3.79 2.8 ;
 RECT 2.535 1.865 2.675 2.8 ;
 RECT 0.61 1.74 0.75 2.8 ;
 RECT 4.95 2.635 5.22 2.8 ;
 RECT 7.035 2.575 7.175 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.24 0.08 ;
 RECT 9.15 0.08 9.29 0.965 ;
 RECT 0.62 0.08 0.76 0.775 ;
 RECT 1.765 0.08 1.905 0.965 ;
 RECT 7.175 0.08 7.445 0.245 ;
 RECT 4.92 0.08 5.19 0.245 ;
 RECT 3.61 0.08 3.88 0.245 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.825 1.155 5.245 1.43 ;
 END
 ANTENNAGATEAREA 0.174 ;
 END IN1

 PIN Q0
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.58 1.08 6.72 1.735 ;
 RECT 6.58 0.77 6.975 0.91 ;
 RECT 6.58 0.91 6.845 1.08 ;
 END
 ANTENNADIFFAREA 0.458 ;
 END Q0

 OBS
 LAYER PO ;
 RECT 7.165 1.47 7.595 1.57 ;
 RECT 7.165 1.57 7.405 1.69 ;
 RECT 8.735 1.38 8.835 2.6 ;
 RECT 7.305 1.69 7.405 2.6 ;
 RECT 7.495 0.51 7.595 1.47 ;
 RECT 8.935 0.53 9.035 1.28 ;
 RECT 8.735 1.28 9.035 1.38 ;
 RECT 7.305 2.6 8.835 2.7 ;
 RECT 4.765 1.215 5.055 1.425 ;
 RECT 4.8 1.43 4.9 2.21 ;
 RECT 4.765 0.38 4.865 1.215 ;
 RECT 4.765 1.425 4.9 1.43 ;
 RECT 4.655 2.21 4.9 2.42 ;
 RECT 1.83 1.325 1.93 2.6 ;
 RECT 3.26 1.38 3.36 2.41 ;
 RECT 1.83 2.6 3.48 2.62 ;
 RECT 3.25 2.41 3.48 2.6 ;
 RECT 1.83 2.62 3.36 2.7 ;
 RECT 2.02 0.53 2.12 1.225 ;
 RECT 3.46 0.53 3.56 1.28 ;
 RECT 1.83 1.225 2.12 1.325 ;
 RECT 3.26 1.28 3.56 1.38 ;
 RECT 7.795 0.53 7.895 2.21 ;
 RECT 7.67 2.21 7.9 2.42 ;
 RECT 2.79 1.1 2.89 2.21 ;
 RECT 3.16 0.53 3.26 1 ;
 RECT 2.79 2.21 3.07 2.42 ;
 RECT 2.79 1 3.26 1.1 ;
 RECT 8.635 0.56 8.735 1 ;
 RECT 8.265 1.1 8.365 2.305 ;
 RECT 8.49 0.35 8.735 0.56 ;
 RECT 8.265 1 8.735 1.1 ;
 RECT 2.32 0.56 2.42 2.305 ;
 RECT 2.32 0.35 2.55 0.56 ;
 RECT 9.39 1.375 9.49 2.79 ;
 RECT 9.405 0.38 9.505 1.135 ;
 RECT 9.39 1.345 9.505 1.375 ;
 RECT 9.275 1.135 9.505 1.345 ;
 RECT 1.36 1.375 1.46 2.79 ;
 RECT 1.55 0.38 1.65 1.135 ;
 RECT 1.42 1.135 1.65 1.275 ;
 RECT 1.36 1.275 1.65 1.375 ;
 RECT 3.915 1.375 4.015 2.79 ;
 RECT 3.93 0.38 4.03 1.065 ;
 RECT 3.915 1.275 4.03 1.375 ;
 RECT 3.8 1.065 4.03 1.275 ;
 RECT 5.245 0.395 5.345 1.33 ;
 RECT 5.275 1.43 5.375 2.125 ;
 RECT 5.275 2.125 5.54 2.335 ;
 RECT 5.245 0.185 5.58 0.395 ;
 RECT 5.245 1.33 5.375 1.43 ;
 RECT 6.835 1.155 7.24 1.275 ;
 RECT 6.835 1.275 6.935 2.79 ;
 RECT 7.025 0.26 7.125 1.065 ;
 RECT 6.885 1.11 7.24 1.155 ;
 RECT 7.01 1.065 7.24 1.11 ;
 LAYER CO ;
 RECT 1.11 1.645 1.24 1.775 ;
 RECT 3.68 0.11 3.81 0.24 ;
 RECT 3.01 1.605 3.14 1.735 ;
 RECT 2.05 1.925 2.18 2.055 ;
 RECT 1.11 1.905 1.24 2.035 ;
 RECT 4.15 0.78 4.28 0.91 ;
 RECT 2.91 0.75 3.04 0.88 ;
 RECT 1.58 1.935 1.71 2.065 ;
 RECT 1.11 2.165 1.24 2.295 ;
 RECT 1.3 0.78 1.43 0.91 ;
 RECT 1.11 2.425 1.24 2.555 ;
 RECT 1.77 0.75 1.9 0.88 ;
 RECT 5.36 2.165 5.49 2.295 ;
 RECT 7.06 1.105 7.19 1.235 ;
 RECT 2.54 1.925 2.67 2.055 ;
 RECT 4.15 1.645 4.28 1.775 ;
 RECT 3.655 2.625 3.785 2.755 ;
 RECT 2.54 0.75 2.67 0.88 ;
 RECT 4.875 1.255 5.005 1.385 ;
 RECT 4.99 0.11 5.12 0.24 ;
 RECT 5.02 2.64 5.15 2.77 ;
 RECT 4.515 0.79 4.645 0.92 ;
 RECT 4.55 1.665 4.68 1.795 ;
 RECT 0.625 0.59 0.755 0.72 ;
 RECT 0.625 0.33 0.755 0.46 ;
 RECT 0.615 2.345 0.745 2.475 ;
 RECT 0.615 2.085 0.745 2.215 ;
 RECT 0.615 1.825 0.745 1.955 ;
 RECT 7.215 1.515 7.345 1.645 ;
 RECT 4.705 2.25 4.835 2.38 ;
 RECT 3.3 2.45 3.43 2.58 ;
 RECT 7.72 2.25 7.85 2.38 ;
 RECT 5.96 0.79 6.09 0.92 ;
 RECT 5.5 1.545 5.63 1.675 ;
 RECT 2.89 2.25 3.02 2.38 ;
 RECT 5.4 0.225 5.53 0.355 ;
 RECT 8.54 0.39 8.67 0.52 ;
 RECT 2.37 0.39 2.5 0.52 ;
 RECT 9.325 1.175 9.455 1.305 ;
 RECT 9.62 1.905 9.75 2.035 ;
 RECT 9.62 2.165 9.75 2.295 ;
 RECT 9.62 1.645 9.75 1.775 ;
 RECT 9.62 2.425 9.75 2.555 ;
 RECT 6.585 1.535 6.715 1.665 ;
 RECT 9.155 0.75 9.285 0.88 ;
 RECT 8.385 0.75 8.515 0.88 ;
 RECT 7.245 0.11 7.375 0.24 ;
 RECT 9.13 1.935 9.26 2.065 ;
 RECT 8.485 1.925 8.615 2.055 ;
 RECT 7.055 2.44 7.185 2.57 ;
 RECT 6.775 0.775 6.905 0.905 ;
 RECT 9.625 0.78 9.755 0.91 ;
 RECT 7.525 1.815 7.655 1.945 ;
 RECT 8.015 1.925 8.145 2.055 ;
 RECT 8.015 0.75 8.145 0.88 ;
 RECT 1.47 1.175 1.6 1.305 ;
 RECT 3.85 1.105 3.98 1.235 ;
 LAYER M1 ;
 RECT 2.045 1.085 2.185 1.17 ;
 RECT 2.045 1.31 2.185 2.13 ;
 RECT 1.4 1.17 2.185 1.31 ;
 RECT 2.535 0.7 2.675 0.945 ;
 RECT 2.045 0.945 2.675 1.085 ;
 RECT 6.58 0.36 6.72 0.385 ;
 RECT 5.33 0.36 5.47 0.385 ;
 RECT 5.33 0.22 6.72 0.36 ;
 RECT 2.3 0.385 5.47 0.525 ;
 RECT 6.58 0.385 8.74 0.525 ;
 RECT 3.295 2.385 3.435 2.66 ;
 RECT 3.295 2.245 4.905 2.385 ;
 RECT 4.545 0.925 4.685 1.66 ;
 RECT 4.48 1.66 4.75 1.8 ;
 RECT 4.445 0.785 5.75 0.925 ;
 RECT 5.61 0.64 5.75 0.785 ;
 RECT 6.3 0.64 6.44 1.875 ;
 RECT 5.61 0.5 6.44 0.64 ;
 RECT 7.21 1.445 7.35 1.875 ;
 RECT 6.3 1.875 7.35 2.015 ;
 RECT 2.885 2.08 3.025 2.465 ;
 RECT 2.885 1.965 5.04 2.08 ;
 RECT 4.9 1.82 5.04 1.825 ;
 RECT 5.495 1.68 5.635 1.825 ;
 RECT 2.885 1.94 6.155 1.965 ;
 RECT 6.015 1.965 6.155 2.155 ;
 RECT 4.9 1.825 6.155 1.94 ;
 RECT 5.955 0.925 6.095 1.065 ;
 RECT 5.495 1.205 5.635 1.54 ;
 RECT 5.89 0.785 6.16 0.925 ;
 RECT 5.495 1.065 6.095 1.205 ;
 RECT 5.43 1.54 5.7 1.68 ;
 RECT 7.715 2.295 7.855 2.45 ;
 RECT 6.015 2.155 7.86 2.29 ;
 RECT 6.02 2.29 7.86 2.295 ;
 RECT 8.48 1.085 8.62 1.17 ;
 RECT 8.48 1.31 8.62 2.13 ;
 RECT 8.38 0.7 8.52 0.945 ;
 RECT 8.38 0.945 8.62 1.085 ;
 RECT 8.48 1.17 9.46 1.31 ;
 RECT 9.32 1.105 9.46 1.17 ;
 RECT 9.32 1.31 9.46 1.38 ;
 RECT 3.005 1.21 3.145 1.6 ;
 RECT 2.905 0.945 3.145 1.07 ;
 RECT 2.905 1.07 3.985 1.085 ;
 RECT 3.005 1.085 3.985 1.21 ;
 RECT 3.845 1.055 3.985 1.07 ;
 RECT 3.845 1.21 3.985 1.335 ;
 RECT 2.905 0.7 3.045 0.945 ;
 RECT 2.94 1.6 3.21 1.74 ;
 RECT 7.52 1.085 7.66 1.13 ;
 RECT 7.52 1.27 7.66 2.015 ;
 RECT 7.01 1.065 7.24 1.13 ;
 RECT 7.01 1.27 7.24 1.275 ;
 RECT 6.985 1.13 7.66 1.27 ;
 RECT 8.01 0.7 8.15 0.945 ;
 RECT 7.52 0.945 8.15 1.085 ;
 END
END DEC24X1

MACRO DEC24X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 12.8 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.6 2.265 6.915 2.645 ;
 END
 ANTENNAGATEAREA 0.188 ;
 END IN2

 PIN Q2
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.75 1.52 5.1 1.795 ;
 RECT 4.87 1.455 5.1 1.52 ;
 RECT 4.87 0.71 5.01 1.455 ;
 END
 ANTENNADIFFAREA 0.678 ;
 END Q2

 PIN Q3
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.83 0.775 2.225 0.915 ;
 RECT 1.83 2.555 1.97 2.62 ;
 RECT 1.61 2.23 1.97 2.555 ;
 RECT 1.83 0.915 1.97 2.23 ;
 END
 ANTENNADIFFAREA 0.7 ;
 END Q3

 PIN Q1
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.485 1.69 11.815 2.05 ;
 RECT 11.585 0.71 11.725 1.69 ;
 END
 ANTENNADIFFAREA 0.642 ;
 END Q1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 12.8 2.96 ;
 RECT 8.9 2.435 9.17 2.575 ;
 RECT 7.96 2.435 8.23 2.575 ;
 RECT 11.065 2.335 11.205 2.8 ;
 RECT 9.925 1.865 10.065 2.8 ;
 RECT 6.295 2.51 6.435 2.8 ;
 RECT 1.31 1.565 1.45 2.8 ;
 RECT 2.3 1.865 2.44 2.8 ;
 RECT 4.375 2.555 4.515 2.8 ;
 RECT 3.26 1.865 3.4 2.8 ;
 RECT 5.435 2.555 5.575 2.8 ;
 RECT 12.095 2.335 12.235 2.8 ;
 RECT 0.585 1.74 0.725 2.8 ;
 RECT 8.965 2.575 9.105 2.8 ;
 RECT 8.025 2.575 8.165 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 12.8 0.08 ;
 RECT 11.02 0.595 11.29 0.735 ;
 RECT 12.015 0.595 12.285 0.735 ;
 RECT 5.35 0.08 5.62 0.245 ;
 RECT 1.315 0.08 1.455 0.99 ;
 RECT 0.595 0.08 0.735 0.775 ;
 RECT 2.49 0.08 2.63 0.965 ;
 RECT 9.09 0.08 9.36 0.245 ;
 RECT 6.195 0.08 6.465 0.245 ;
 RECT 4.335 0.08 4.605 0.245 ;
 RECT 8.17 0.08 8.44 0.245 ;
 RECT 11.085 0.08 11.225 0.595 ;
 RECT 12.08 0.08 12.22 0.595 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.1 1.155 6.395 1.48 ;
 END
 ANTENNAGATEAREA 0.188 ;
 END IN1

 PIN Q0
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.495 0.67 8.955 0.96 ;
 RECT 8.495 0.96 8.635 1.735 ;
 END
 ANTENNADIFFAREA 0.562 ;
 END Q0

 OBS
 LAYER PO ;
 RECT 10.65 1.38 10.75 2.6 ;
 RECT 9.22 1.695 9.32 2.6 ;
 RECT 9.22 1.305 9.32 1.485 ;
 RECT 9.08 1.485 9.32 1.695 ;
 RECT 10.85 0.53 10.95 1.28 ;
 RECT 10.65 1.28 10.95 1.38 ;
 RECT 9.41 0.51 9.51 1.205 ;
 RECT 9.22 2.6 10.75 2.7 ;
 RECT 9.22 1.205 9.51 1.305 ;
 RECT 2.555 1.325 2.655 2.6 ;
 RECT 3.985 1.38 4.085 2.41 ;
 RECT 2.555 2.6 4.205 2.62 ;
 RECT 3.975 2.41 4.205 2.6 ;
 RECT 2.555 2.62 4.085 2.7 ;
 RECT 2.745 0.53 2.845 1.225 ;
 RECT 4.185 0.53 4.285 1.28 ;
 RECT 2.555 1.225 2.845 1.325 ;
 RECT 3.985 1.28 4.285 1.38 ;
 RECT 9.71 0.53 9.81 2.21 ;
 RECT 9.585 2.21 9.815 2.42 ;
 RECT 3.515 1.1 3.615 2.21 ;
 RECT 3.885 0.53 3.985 1 ;
 RECT 3.515 2.21 3.795 2.42 ;
 RECT 3.515 1 3.985 1.1 ;
 RECT 10.55 0.565 10.65 1 ;
 RECT 10.18 1.1 10.28 2.305 ;
 RECT 10.18 1 10.65 1.1 ;
 RECT 10.405 0.35 10.65 0.565 ;
 RECT 3.045 0.56 3.145 2.305 ;
 RECT 3.045 0.35 3.275 0.56 ;
 RECT 11.85 1.375 11.95 2.79 ;
 RECT 11.325 1.41 11.425 2.79 ;
 RECT 11.195 1.275 11.965 1.375 ;
 RECT 11.35 0.38 11.45 1.2 ;
 RECT 11.195 1.2 11.45 1.275 ;
 RECT 11.195 1.375 11.425 1.41 ;
 RECT 11.865 0.38 11.965 1.275 ;
 RECT 8.28 1.205 9.04 1.305 ;
 RECT 8.47 0.35 8.57 1.205 ;
 RECT 8.81 1.095 9.04 1.155 ;
 RECT 8.28 1.305 8.38 2.79 ;
 RECT 8.75 1.305 8.85 2.79 ;
 RECT 8.94 0.26 9.04 1.095 ;
 RECT 8.75 1.155 9.04 1.205 ;
 RECT 1.575 1.275 2.375 1.375 ;
 RECT 1.575 1.375 1.675 2.79 ;
 RECT 1.575 0.35 1.675 1.275 ;
 RECT 2.085 1.375 2.185 2.79 ;
 RECT 2.275 0.38 2.375 1.135 ;
 RECT 2.145 1.135 2.375 1.275 ;
 RECT 5.19 1.375 5.29 2.79 ;
 RECT 5.19 0.38 5.29 1.275 ;
 RECT 4.64 1.375 4.74 2.79 ;
 RECT 4.655 0.38 4.755 1.135 ;
 RECT 4.64 1.345 5.29 1.375 ;
 RECT 4.525 1.275 5.29 1.345 ;
 RECT 4.525 1.135 4.755 1.275 ;
 RECT 6.55 2.435 6.915 2.645 ;
 RECT 6.55 1.43 6.65 2.435 ;
 RECT 6.52 0.395 6.62 1.33 ;
 RECT 6.52 0.185 6.855 0.395 ;
 RECT 6.52 1.33 6.65 1.43 ;
 RECT 6.04 1.22 6.29 1.43 ;
 RECT 6.075 1.43 6.175 2.275 ;
 RECT 5.93 2.275 6.175 2.485 ;
 RECT 6.04 0.38 6.14 1.22 ;
 LAYER CO ;
 RECT 4.38 2.625 4.51 2.755 ;
 RECT 3.265 0.75 3.395 0.88 ;
 RECT 6.72 2.475 6.85 2.605 ;
 RECT 6.11 1.26 6.24 1.39 ;
 RECT 6.265 0.11 6.395 0.24 ;
 RECT 6.3 2.64 6.43 2.77 ;
 RECT 5.79 0.79 5.92 0.92 ;
 RECT 5.825 1.665 5.955 1.795 ;
 RECT 0.6 0.59 0.73 0.72 ;
 RECT 0.6 0.33 0.73 0.46 ;
 RECT 0.59 2.345 0.72 2.475 ;
 RECT 0.59 2.085 0.72 2.215 ;
 RECT 0.59 1.825 0.72 1.955 ;
 RECT 9.13 1.525 9.26 1.655 ;
 RECT 5.98 2.315 6.11 2.445 ;
 RECT 4.025 2.45 4.155 2.58 ;
 RECT 9.635 2.25 9.765 2.38 ;
 RECT 7.235 0.79 7.365 0.92 ;
 RECT 6.775 1.83 6.905 1.96 ;
 RECT 12.1 2.41 12.23 2.54 ;
 RECT 12.085 0.6 12.215 0.73 ;
 RECT 11.59 1.785 11.72 1.915 ;
 RECT 11.59 0.78 11.72 0.91 ;
 RECT 8.24 0.11 8.37 0.24 ;
 RECT 8.03 2.44 8.16 2.57 ;
 RECT 5.42 0.11 5.55 0.24 ;
 RECT 1.315 1.645 1.445 1.775 ;
 RECT 1.315 2.17 1.445 2.3 ;
 RECT 1.315 1.91 1.445 2.04 ;
 RECT 1.32 0.78 1.45 0.91 ;
 RECT 5.44 2.625 5.57 2.755 ;
 RECT 3.615 2.25 3.745 2.38 ;
 RECT 6.675 0.225 6.805 0.355 ;
 RECT 10.455 0.39 10.585 0.52 ;
 RECT 3.095 0.39 3.225 0.52 ;
 RECT 11.245 1.24 11.375 1.37 ;
 RECT 8.5 1.535 8.63 1.665 ;
 RECT 11.09 0.6 11.22 0.73 ;
 RECT 10.3 0.75 10.43 0.88 ;
 RECT 9.16 0.11 9.29 0.24 ;
 RECT 11.07 2.41 11.2 2.54 ;
 RECT 10.4 1.925 10.53 2.055 ;
 RECT 8.86 1.135 8.99 1.265 ;
 RECT 8.97 2.44 9.1 2.57 ;
 RECT 8.69 0.775 8.82 0.905 ;
 RECT 9.44 1.815 9.57 1.945 ;
 RECT 9.93 1.925 10.06 2.055 ;
 RECT 9.93 0.75 10.06 0.88 ;
 RECT 2.195 1.175 2.325 1.305 ;
 RECT 4.575 1.175 4.705 1.305 ;
 RECT 1.835 1.645 1.965 1.775 ;
 RECT 4.405 0.11 4.535 0.24 ;
 RECT 3.735 1.605 3.865 1.735 ;
 RECT 2.775 1.925 2.905 2.055 ;
 RECT 1.835 1.905 1.965 2.035 ;
 RECT 4.875 0.78 5.005 0.91 ;
 RECT 3.635 0.75 3.765 0.88 ;
 RECT 2.305 1.935 2.435 2.065 ;
 RECT 1.835 2.165 1.965 2.295 ;
 RECT 2.025 0.78 2.155 0.91 ;
 RECT 1.835 2.425 1.965 2.555 ;
 RECT 2.495 0.75 2.625 0.88 ;
 RECT 3.265 1.925 3.395 2.055 ;
 RECT 4.86 1.645 4.99 1.775 ;
 LAYER M1 ;
 RECT 2.77 1.085 2.91 1.17 ;
 RECT 2.77 1.31 2.91 2.13 ;
 RECT 2.125 1.17 2.91 1.31 ;
 RECT 3.26 0.7 3.4 0.945 ;
 RECT 2.77 0.945 3.4 1.085 ;
 RECT 3.73 1.085 3.87 1.17 ;
 RECT 3.73 1.17 4.71 1.31 ;
 RECT 3.73 1.31 3.87 1.6 ;
 RECT 4.57 1.105 4.71 1.17 ;
 RECT 4.57 1.31 4.71 1.38 ;
 RECT 3.63 0.7 3.77 0.945 ;
 RECT 3.63 0.945 3.87 1.085 ;
 RECT 3.665 1.6 3.935 1.74 ;
 RECT 7.855 0.36 7.995 0.385 ;
 RECT 6.605 0.22 7.995 0.36 ;
 RECT 6.605 0.36 6.745 0.385 ;
 RECT 3.03 0.385 6.745 0.525 ;
 RECT 7.855 0.385 10.65 0.525 ;
 RECT 4.02 2.385 4.16 2.66 ;
 RECT 5.975 2.385 6.115 2.515 ;
 RECT 4.02 2.245 6.115 2.385 ;
 RECT 3.61 2.08 3.75 2.465 ;
 RECT 7.23 0.925 7.37 1.065 ;
 RECT 6.77 1.205 6.91 1.94 ;
 RECT 7.075 2.08 7.215 2.155 ;
 RECT 7.165 0.785 7.435 0.925 ;
 RECT 6.77 1.065 7.37 1.205 ;
 RECT 3.61 1.94 7.215 2.08 ;
 RECT 9.63 2.295 9.77 2.45 ;
 RECT 7.075 2.155 9.775 2.295 ;
 RECT 5.82 0.925 5.96 1.66 ;
 RECT 5.755 1.66 6.025 1.8 ;
 RECT 5.72 0.785 7.025 0.925 ;
 RECT 6.885 0.64 7.025 0.785 ;
 RECT 7.575 0.64 7.715 1.875 ;
 RECT 6.885 0.5 7.715 0.64 ;
 RECT 7.575 1.875 9.265 2.015 ;
 RECT 9.125 1.455 9.265 1.875 ;
 RECT 10.395 1.085 10.535 1.235 ;
 RECT 10.395 1.375 10.535 2.13 ;
 RECT 10.295 0.7 10.435 0.945 ;
 RECT 10.295 0.945 10.535 1.085 ;
 RECT 10.395 1.235 11.445 1.375 ;
 RECT 9.435 1.085 9.575 1.13 ;
 RECT 9.435 1.27 9.575 2.015 ;
 RECT 8.79 1.13 9.575 1.27 ;
 RECT 9.925 0.7 10.065 0.945 ;
 RECT 9.435 0.945 10.065 1.085 ;
 END
END DEC24X2

MACRO DFFARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.2 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.2 2.96 ;
 RECT 1.945 2.34 2.195 2.8 ;
 RECT 5.355 2.635 5.615 2.8 ;
 RECT 8.005 1.955 8.145 2.8 ;
 RECT 9.185 2.06 9.325 2.8 ;
 RECT 10.71 1.73 10.85 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.27 1.98 1.41 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.2 0.08 ;
 RECT 4.615 0.08 4.85 0.595 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 9.205 0.08 9.345 0.67 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 8.1 0.08 8.24 0.6 ;
 RECT 2.015 0.08 2.155 0.39 ;
 RECT 10.795 0.08 10.935 0.88 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.475 1.65 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.96 0.36 6.2 0.6 ;
 RECT 4.055 0.735 5.13 0.875 ;
 RECT 7.66 0.36 7.8 0.785 ;
 RECT 7.66 0.785 8.635 0.925 ;
 RECT 8.495 0.225 8.635 0.785 ;
 RECT 4.99 0.36 5.13 0.735 ;
 RECT 4.055 0.445 4.195 0.735 ;
 RECT 4.99 0.22 7.8 0.36 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.85 0.55 9.99 2.07 ;
 RECT 9.64 2.07 9.99 2.57 ;
 END
 ANTENNADIFFAREA 0.505 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.235 2.015 10.545 2.38 ;
 RECT 10.235 2.38 10.375 2.61 ;
 RECT 10.235 0.7 10.375 2.015 ;
 END
 ANTENNADIFFAREA 0.483 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.765 0.22 1.13 0.615 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 6.53 0.69 6.63 1.35 ;
 RECT 5.52 0.46 5.75 0.575 ;
 RECT 5.52 0.575 6.63 0.69 ;
 RECT 6.72 1.45 7.075 1.545 ;
 RECT 6.53 0.165 7.965 0.265 ;
 RECT 6.53 1.35 6.82 1.445 ;
 RECT 6.53 1.445 7.075 1.45 ;
 RECT 0.815 0.27 1.155 0.52 ;
 RECT 1.055 0.52 1.155 2.465 ;
 RECT 1.53 0.655 1.63 1.495 ;
 RECT 1.335 1.495 1.63 1.745 ;
 RECT 1.53 1.745 1.63 2.37 ;
 RECT 4.425 0.285 4.525 1.24 ;
 RECT 2.69 0.185 4.525 0.285 ;
 RECT 2.69 0.285 2.79 0.51 ;
 RECT 2.65 0.51 2.895 0.755 ;
 RECT 3.685 1.33 3.825 1.475 ;
 RECT 3.685 1.71 3.785 2.475 ;
 RECT 3.725 0.65 3.825 1.33 ;
 RECT 3.685 1.475 3.915 1.71 ;
 RECT 3.19 1.595 3.29 2.48 ;
 RECT 2.65 1.445 2.895 1.495 ;
 RECT 2.65 1.495 3.29 1.595 ;
 RECT 2.65 1.595 2.895 1.69 ;
 RECT 7.79 1.575 7.89 2.585 ;
 RECT 6.57 2.47 6.79 2.585 ;
 RECT 6.57 2.685 6.79 2.71 ;
 RECT 6.57 2.585 7.89 2.685 ;
 RECT 10.495 0.315 10.595 1.19 ;
 RECT 10.495 1.425 10.595 2.79 ;
 RECT 10.48 1.19 10.69 1.425 ;
 RECT 9.635 0.135 9.735 1.05 ;
 RECT 9.635 1.28 9.735 2.79 ;
 RECT 9.27 1.05 9.735 1.28 ;
 RECT 6.095 1.64 6.48 1.87 ;
 RECT 6.095 1.105 6.35 1.64 ;
 RECT 5.95 0.875 6.35 1.105 ;
 RECT 1.87 1.52 2.47 1.62 ;
 RECT 3.235 0.47 3.52 0.705 ;
 RECT 3.235 0.705 3.335 1.165 ;
 RECT 2.305 1.62 2.405 2.68 ;
 RECT 4.985 1.79 5.085 2.68 ;
 RECT 2.37 0.585 2.47 1.165 ;
 RECT 2.37 1.265 2.47 1.52 ;
 RECT 1.87 1.44 2.115 1.52 ;
 RECT 1.87 1.62 2.115 1.69 ;
 RECT 2.305 2.68 5.085 2.78 ;
 RECT 2.37 1.165 3.335 1.265 ;
 RECT 8.88 1.32 8.98 2.7 ;
 RECT 8.58 0.47 8.68 1.22 ;
 RECT 8.58 1.22 8.98 1.32 ;
 RECT 8.45 0.23 8.68 0.47 ;
 RECT 4.125 0.695 4.225 1.61 ;
 RECT 4.16 1.71 4.26 2.48 ;
 RECT 4.125 1.61 4.26 1.71 ;
 RECT 4.005 0.465 4.245 0.695 ;
 RECT 7.47 0.645 7.57 1.18 ;
 RECT 7.47 1.39 7.57 2.295 ;
 RECT 7.45 1.18 7.685 1.39 ;
 RECT 7 0.685 7.1 1.255 ;
 RECT 6.925 0.455 7.155 0.685 ;
 RECT 8.28 0.65 8.38 1.71 ;
 RECT 8.28 1.71 8.525 1.95 ;
 RECT 8.28 1.95 8.38 2.7 ;
 RECT 5.29 1.61 5.555 1.82 ;
 RECT 5.455 1.82 5.555 2.49 ;
 RECT 5.085 0.635 5.185 1.51 ;
 RECT 5.085 1.51 5.555 1.61 ;
 RECT 6.975 1.545 7.075 2.405 ;
 RECT 7.865 0.265 7.965 1.32 ;
 RECT 6.53 0.265 6.63 0.575 ;
 LAYER CO ;
 RECT 6.02 0.915 6.15 1.045 ;
 RECT 8.5 0.285 8.63 0.415 ;
 RECT 8.105 0.4 8.235 0.53 ;
 RECT 4.06 0.515 4.19 0.645 ;
 RECT 4.665 0.455 4.795 0.585 ;
 RECT 7.22 1.875 7.35 2.005 ;
 RECT 7.22 0.87 7.35 1 ;
 RECT 6.75 0.87 6.88 1 ;
 RECT 6.975 0.505 7.105 0.635 ;
 RECT 8.8 0.87 8.93 1 ;
 RECT 8.01 2.01 8.14 2.14 ;
 RECT 9.19 2.19 9.32 2.32 ;
 RECT 8.63 2.17 8.76 2.3 ;
 RECT 5.345 1.63 5.475 1.76 ;
 RECT 3.735 1.525 3.865 1.655 ;
 RECT 0.875 0.325 1.005 0.455 ;
 RECT 5.68 0.88 5.81 1.01 ;
 RECT 5.675 2.015 5.805 2.145 ;
 RECT 2.02 0.21 2.15 0.34 ;
 RECT 5.405 2.64 5.535 2.77 ;
 RECT 4.735 2.125 4.865 2.255 ;
 RECT 4.385 1.825 4.515 1.955 ;
 RECT 10.715 1.8 10.845 1.93 ;
 RECT 10.715 2.06 10.845 2.19 ;
 RECT 2.94 2.105 3.07 2.235 ;
 RECT 2.985 0.88 3.115 1.01 ;
 RECT 2.705 1.49 2.835 1.62 ;
 RECT 2.59 0.905 2.72 1.035 ;
 RECT 1.75 1.995 1.88 2.125 ;
 RECT 1.88 0.875 2.01 1.005 ;
 RECT 7.5 1.22 7.63 1.35 ;
 RECT 1.275 2.05 1.405 2.18 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 0.805 2.115 0.935 2.245 ;
 RECT 1.395 1.55 1.525 1.68 ;
 RECT 10.24 1.565 10.37 1.695 ;
 RECT 10.24 1.83 10.37 1.96 ;
 RECT 10.24 2.09 10.37 2.22 ;
 RECT 10.24 2.39 10.37 2.52 ;
 RECT 9.855 2.085 9.985 2.215 ;
 RECT 2.705 0.555 2.835 0.685 ;
 RECT 5.56 0.51 5.69 0.64 ;
 RECT 8.35 1.765 8.48 1.895 ;
 RECT 2.525 1.825 2.655 1.955 ;
 RECT 3.34 0.525 3.47 0.655 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 6.62 2.525 6.75 2.655 ;
 RECT 6.725 1.815 6.855 1.945 ;
 RECT 10.52 1.24 10.65 1.37 ;
 RECT 10.8 0.68 10.93 0.81 ;
 RECT 9.855 2.35 9.985 2.48 ;
 RECT 10.715 2.32 10.845 2.45 ;
 RECT 10.24 0.75 10.37 0.88 ;
 RECT 9.32 1.1 9.45 1.23 ;
 RECT 9.855 0.615 9.985 0.745 ;
 RECT 9.855 1.535 9.985 1.665 ;
 RECT 9.855 1.795 9.985 1.925 ;
 RECT 9.21 0.485 9.34 0.615 ;
 RECT 6.3 1.69 6.43 1.82 ;
 RECT 3.905 2.125 4.035 2.255 ;
 RECT 1.93 1.495 2.06 1.625 ;
 RECT 2.015 2.345 2.145 2.475 ;
 RECT 3.435 2.07 3.565 2.2 ;
 RECT 3.455 0.88 3.585 1.01 ;
 LAYER M1 ;
 RECT 3.835 2.12 4.935 2.26 ;
 RECT 5.67 1.05 5.81 1.3 ;
 RECT 4.395 1.3 5.81 1.44 ;
 RECT 5.67 1.44 5.81 2.215 ;
 RECT 5.61 0.91 6.22 1.015 ;
 RECT 5.61 0.875 5.88 0.91 ;
 RECT 5.67 1.015 6.22 1.05 ;
 RECT 3.665 1.52 4.535 1.66 ;
 RECT 4.395 1.44 4.535 1.52 ;
 RECT 3.27 0.52 3.915 0.66 ;
 RECT 3.775 0.66 3.915 1.015 ;
 RECT 3.775 1.015 5.41 1.155 ;
 RECT 5.27 0.505 5.75 0.645 ;
 RECT 5.27 0.645 5.41 1.015 ;
 RECT 7.495 1.395 8.935 1.535 ;
 RECT 8.795 0.955 8.935 1.395 ;
 RECT 8.625 1.535 8.765 2.36 ;
 RECT 7.495 1.17 7.635 1.395 ;
 RECT 9.485 0.36 9.625 0.815 ;
 RECT 8.795 0.815 9.625 0.955 ;
 RECT 10.515 0.36 10.655 1.45 ;
 RECT 9.485 0.22 10.655 0.36 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.11 ;
 RECT 0.58 2.25 0.72 2.255 ;
 RECT 0.58 2.11 1.005 2.25 ;
 RECT 0.58 0.87 1.005 1.01 ;
 RECT 1.55 0.67 1.69 1.195 ;
 RECT 0.58 1.195 1.69 1.335 ;
 RECT 2.98 0.36 3.12 2.035 ;
 RECT 1.55 0.53 2.435 0.67 ;
 RECT 2.295 0.22 3.12 0.36 ;
 RECT 2.295 0.36 2.435 0.53 ;
 RECT 2.935 2.035 3.12 2.17 ;
 RECT 2.935 2.17 3.075 2.305 ;
 RECT 3.275 1.22 3.59 1.36 ;
 RECT 3.45 0.805 3.59 1.22 ;
 RECT 3.36 1.96 3.64 2.215 ;
 RECT 3.275 1.36 3.415 1.82 ;
 RECT 3.275 1.82 5.48 1.96 ;
 RECT 5.34 1.58 5.48 1.82 ;
 RECT 7.215 1.815 7.425 1.87 ;
 RECT 7.215 0.805 7.355 1.675 ;
 RECT 7.145 1.87 7.425 2.01 ;
 RECT 8.905 1.92 9.045 2.505 ;
 RECT 7.215 1.675 8.485 1.815 ;
 RECT 8.345 2.505 9.045 2.645 ;
 RECT 8.345 1.815 8.485 2.505 ;
 RECT 9.14 1.235 9.28 1.78 ;
 RECT 9.14 1.095 9.52 1.235 ;
 RECT 8.905 1.78 9.28 1.92 ;
 RECT 6.23 1.685 6.885 1.81 ;
 RECT 6.745 1.005 6.885 1.685 ;
 RECT 6.23 1.81 6.925 1.825 ;
 RECT 6.655 1.825 6.925 1.95 ;
 RECT 6.675 0.865 6.955 1.005 ;
 RECT 2.585 0.5 2.84 0.965 ;
 RECT 2.585 1.96 2.725 2.51 ;
 RECT 2.585 1.67 2.725 1.82 ;
 RECT 2.585 0.965 2.725 1.44 ;
 RECT 2.585 1.44 2.84 1.67 ;
 RECT 2.455 1.82 2.725 1.96 ;
 RECT 2.585 2.51 5.215 2.65 ;
 RECT 5.075 2.495 5.215 2.51 ;
 RECT 5.95 1.21 6.53 1.35 ;
 RECT 6.55 2.24 6.69 2.52 ;
 RECT 5.95 1.35 6.09 2.1 ;
 RECT 5.95 2.24 6.09 2.355 ;
 RECT 5.95 2.1 6.69 2.24 ;
 RECT 5.075 2.355 6.09 2.495 ;
 RECT 6.67 0.5 7.18 0.58 ;
 RECT 6.39 0.58 7.18 0.64 ;
 RECT 6.39 0.64 6.85 0.72 ;
 RECT 6.39 0.72 6.53 1.21 ;
 RECT 6.55 2.52 6.82 2.66 ;
 RECT 1.79 1.63 1.93 1.99 ;
 RECT 1.79 1.475 2.135 1.63 ;
 RECT 1.875 0.825 2.015 1.475 ;
 RECT 1.68 1.99 1.93 2.13 ;
 END
END DFFARX1

MACRO DFFARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.84 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.84 2.96 ;
 RECT 5.355 2.635 5.615 2.8 ;
 RECT 1.945 2.34 2.195 2.8 ;
 RECT 1.27 1.98 1.41 2.8 ;
 RECT 8.005 1.955 8.145 2.8 ;
 RECT 9.185 2.06 9.325 2.8 ;
 RECT 11.285 1.73 11.425 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 10.32 1.485 10.46 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.84 0.08 ;
 RECT 4.615 0.08 4.85 0.595 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 11.595 0.08 11.735 0.88 ;
 RECT 9.205 0.08 9.345 0.67 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 8.1 0.08 8.24 0.6 ;
 RECT 2.015 0.08 2.155 0.39 ;
 RECT 10.475 0.08 10.615 0.3 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.475 1.645 1.76 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.925 0.36 6.26 0.46 ;
 RECT 7.66 0.36 7.8 0.785 ;
 RECT 4.055 0.735 5.13 0.875 ;
 RECT 7.66 0.785 8.635 0.925 ;
 RECT 8.495 0.225 8.635 0.785 ;
 RECT 4.99 0.36 5.13 0.735 ;
 RECT 4.99 0.22 7.8 0.36 ;
 RECT 4.055 0.445 4.195 0.735 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.85 0.72 9.99 2.07 ;
 RECT 9.64 2.07 9.99 2.57 ;
 END
 ANTENNADIFFAREA 0.616 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.6 2.015 10.95 2.38 ;
 RECT 10.81 0.845 11.11 0.985 ;
 RECT 10.81 2.38 10.95 2.61 ;
 RECT 10.97 0.72 11.11 0.845 ;
 RECT 10.81 0.985 10.95 2.015 ;
 END
 ANTENNADIFFAREA 0.642 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 0.36 1.13 0.61 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 8.28 0.65 8.38 1.71 ;
 RECT 8.28 1.71 8.525 1.95 ;
 RECT 8.28 1.95 8.38 2.7 ;
 RECT 5.29 1.61 5.555 1.82 ;
 RECT 5.455 1.82 5.555 2.49 ;
 RECT 5.085 0.635 5.185 1.51 ;
 RECT 5.085 1.51 5.555 1.61 ;
 RECT 11.07 1.265 11.48 1.425 ;
 RECT 10.575 1.265 10.675 2.79 ;
 RECT 10.575 1.165 11.48 1.265 ;
 RECT 10.755 0.38 10.855 1.165 ;
 RECT 11.38 0.38 11.48 1.165 ;
 RECT 11.07 1.425 11.17 2.79 ;
 RECT 1.87 1.52 2.47 1.62 ;
 RECT 3.235 0.47 3.52 0.705 ;
 RECT 3.235 0.705 3.335 1.165 ;
 RECT 2.37 0.585 2.47 1.165 ;
 RECT 2.37 1.265 2.47 1.52 ;
 RECT 2.305 1.62 2.405 2.68 ;
 RECT 4.985 1.79 5.085 2.68 ;
 RECT 1.87 1.44 2.115 1.52 ;
 RECT 1.87 1.62 2.115 1.69 ;
 RECT 2.37 1.165 3.335 1.265 ;
 RECT 2.305 2.68 5.085 2.78 ;
 RECT 5.555 0.59 6.63 0.69 ;
 RECT 6.53 0.69 6.63 1.35 ;
 RECT 6.975 1.545 7.075 2.405 ;
 RECT 7.865 0.265 7.965 1.22 ;
 RECT 5.555 0.46 5.785 0.59 ;
 RECT 6.53 0.265 6.63 0.59 ;
 RECT 6.53 0.165 7.965 0.265 ;
 RECT 6.72 1.45 7.075 1.545 ;
 RECT 6.53 1.35 6.82 1.445 ;
 RECT 6.53 1.445 7.075 1.45 ;
 RECT 3.685 1.33 3.825 1.475 ;
 RECT 3.685 1.71 3.785 2.475 ;
 RECT 3.725 0.65 3.825 1.33 ;
 RECT 3.685 1.475 3.915 1.71 ;
 RECT 9.27 1.05 9.735 1.09 ;
 RECT 9.27 1.09 10.205 1.19 ;
 RECT 9.635 0.135 9.735 1.05 ;
 RECT 9.635 1.28 9.735 2.79 ;
 RECT 9.27 1.19 9.735 1.28 ;
 RECT 10.105 0.135 10.205 1.09 ;
 RECT 10.105 1.19 10.205 2.79 ;
 RECT 0.84 0.36 1.155 0.61 ;
 RECT 1.055 0.61 1.155 2.465 ;
 RECT 1.53 0.655 1.63 1.495 ;
 RECT 1.335 1.495 1.63 1.745 ;
 RECT 1.53 1.745 1.63 2.37 ;
 RECT 7.47 0.645 7.57 1.18 ;
 RECT 7.47 1.39 7.57 2.295 ;
 RECT 7.45 1.18 7.685 1.39 ;
 RECT 7 0.685 7.1 1.255 ;
 RECT 6.925 0.455 7.155 0.685 ;
 RECT 2.69 0.285 2.79 0.51 ;
 RECT 2.69 0.185 4.525 0.285 ;
 RECT 4.425 0.285 4.525 1.24 ;
 RECT 2.65 0.51 2.895 0.755 ;
 RECT 7.79 1.575 7.89 2.585 ;
 RECT 6.57 2.47 6.79 2.585 ;
 RECT 6.57 2.685 6.79 2.71 ;
 RECT 6.57 2.585 7.89 2.685 ;
 RECT 6.09 1.64 6.48 1.87 ;
 RECT 6.09 1.105 6.35 1.64 ;
 RECT 5.95 0.875 6.35 1.105 ;
 RECT 8.88 1.32 8.98 2.7 ;
 RECT 8.58 0.47 8.68 1.22 ;
 RECT 8.58 1.22 8.98 1.32 ;
 RECT 8.45 0.23 8.68 0.47 ;
 RECT 4.125 0.695 4.225 1.61 ;
 RECT 4.16 1.71 4.26 2.48 ;
 RECT 4.125 1.61 4.26 1.71 ;
 RECT 4.005 0.465 4.245 0.695 ;
 RECT 3.19 1.595 3.29 2.48 ;
 RECT 2.65 1.445 2.895 1.495 ;
 RECT 2.65 1.595 2.895 1.69 ;
 RECT 2.65 1.495 3.29 1.595 ;
 LAYER CO ;
 RECT 9.855 1.535 9.985 1.665 ;
 RECT 9.855 1.795 9.985 1.925 ;
 RECT 9.21 0.485 9.34 0.615 ;
 RECT 6.3 1.69 6.43 1.82 ;
 RECT 4.385 1.825 4.515 1.955 ;
 RECT 3.905 2.125 4.035 2.255 ;
 RECT 1.93 1.495 2.06 1.625 ;
 RECT 2.015 2.345 2.145 2.475 ;
 RECT 3.435 2.07 3.565 2.2 ;
 RECT 3.455 0.88 3.585 1.01 ;
 RECT 2.94 2.105 3.07 2.235 ;
 RECT 1.88 0.875 2.01 1.005 ;
 RECT 1.275 2.05 1.405 2.18 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 0.805 2.115 0.935 2.245 ;
 RECT 10.48 0.12 10.61 0.25 ;
 RECT 5.68 0.88 5.81 1.01 ;
 RECT 10.325 1.535 10.455 1.665 ;
 RECT 5.405 2.64 5.535 2.77 ;
 RECT 4.735 2.125 4.865 2.255 ;
 RECT 0.9 0.415 1.03 0.545 ;
 RECT 1.395 1.55 1.525 1.68 ;
 RECT 10.815 1.565 10.945 1.695 ;
 RECT 10.815 1.83 10.945 1.96 ;
 RECT 10.815 2.09 10.945 2.22 ;
 RECT 2.705 0.555 2.835 0.685 ;
 RECT 5.595 0.51 5.725 0.64 ;
 RECT 6.975 0.505 7.105 0.635 ;
 RECT 7.5 1.22 7.63 1.35 ;
 RECT 3.34 0.525 3.47 0.655 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 6.62 2.525 6.75 2.655 ;
 RECT 6.725 1.815 6.855 1.945 ;
 RECT 11.13 1.24 11.26 1.37 ;
 RECT 11.6 0.68 11.73 0.81 ;
 RECT 9.855 2.35 9.985 2.48 ;
 RECT 11.29 2.32 11.42 2.45 ;
 RECT 10.975 0.77 11.105 0.9 ;
 RECT 9.32 1.1 9.45 1.23 ;
 RECT 11.29 1.8 11.42 1.93 ;
 RECT 11.29 2.06 11.42 2.19 ;
 RECT 9.855 0.77 9.985 0.9 ;
 RECT 10.325 2.085 10.455 2.215 ;
 RECT 10.325 1.795 10.455 1.925 ;
 RECT 10.325 2.35 10.455 2.48 ;
 RECT 6.02 0.915 6.15 1.045 ;
 RECT 8.5 0.285 8.63 0.415 ;
 RECT 8.105 0.4 8.235 0.53 ;
 RECT 4.06 0.515 4.19 0.645 ;
 RECT 4.665 0.455 4.795 0.585 ;
 RECT 7.22 1.875 7.35 2.005 ;
 RECT 7.22 0.87 7.35 1 ;
 RECT 6.75 0.87 6.88 1 ;
 RECT 2.985 0.88 3.115 1.01 ;
 RECT 2.705 1.49 2.835 1.62 ;
 RECT 2.59 0.905 2.72 1.035 ;
 RECT 1.75 1.995 1.88 2.125 ;
 RECT 8.8 0.87 8.93 1 ;
 RECT 8.01 2.01 8.14 2.14 ;
 RECT 9.19 2.19 9.32 2.32 ;
 RECT 8.63 2.17 8.76 2.3 ;
 RECT 5.345 1.63 5.475 1.76 ;
 RECT 3.735 1.525 3.865 1.655 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 5.675 2.015 5.805 2.145 ;
 RECT 2.02 0.21 2.15 0.34 ;
 RECT 10.815 2.39 10.945 2.52 ;
 RECT 9.855 2.085 9.985 2.215 ;
 RECT 8.35 1.765 8.48 1.895 ;
 RECT 2.525 1.825 2.655 1.955 ;
 LAYER M1 ;
 RECT 3.835 2.12 4.935 2.26 ;
 RECT 3.27 0.52 3.915 0.66 ;
 RECT 3.775 0.66 3.915 1.015 ;
 RECT 3.775 1.015 5.41 1.155 ;
 RECT 5.27 0.505 5.785 0.645 ;
 RECT 5.27 0.645 5.41 1.015 ;
 RECT 5.67 1.015 6.22 1.05 ;
 RECT 5.67 1.05 5.81 1.3 ;
 RECT 5.61 0.91 6.22 1.015 ;
 RECT 5.61 0.875 5.88 0.91 ;
 RECT 4.395 1.3 5.81 1.44 ;
 RECT 5.67 1.44 5.81 2.215 ;
 RECT 4.395 1.44 4.535 1.52 ;
 RECT 3.665 1.52 4.535 1.66 ;
 RECT 1.79 1.63 1.93 1.99 ;
 RECT 1.79 1.475 2.135 1.63 ;
 RECT 1.875 0.825 2.015 1.475 ;
 RECT 1.68 1.99 1.93 2.13 ;
 RECT 7.495 1.395 8.935 1.535 ;
 RECT 8.795 0.955 8.935 1.395 ;
 RECT 8.625 1.535 8.765 2.36 ;
 RECT 7.495 1.17 7.635 1.395 ;
 RECT 9.485 0.58 9.625 0.815 ;
 RECT 8.795 0.815 9.625 0.955 ;
 RECT 11.25 0.58 11.39 1.17 ;
 RECT 11.125 1.17 11.39 1.235 ;
 RECT 9.485 0.44 11.39 0.58 ;
 RECT 11.125 1.375 11.39 1.44 ;
 RECT 11.09 1.235 11.39 1.375 ;
 RECT 7.215 1.815 7.425 1.87 ;
 RECT 7.215 0.805 7.355 1.675 ;
 RECT 7.145 1.87 7.425 2.01 ;
 RECT 8.905 1.92 9.045 2.505 ;
 RECT 7.215 1.675 8.485 1.815 ;
 RECT 8.345 2.505 9.045 2.645 ;
 RECT 8.345 1.815 8.485 2.505 ;
 RECT 9.14 1.235 9.28 1.78 ;
 RECT 9.14 1.095 9.52 1.235 ;
 RECT 8.905 1.78 9.28 1.92 ;
 RECT 6.23 1.685 6.885 1.81 ;
 RECT 6.745 1.005 6.885 1.685 ;
 RECT 6.23 1.81 6.925 1.825 ;
 RECT 6.655 1.825 6.925 1.95 ;
 RECT 6.675 0.865 6.955 1.005 ;
 RECT 3.36 1.96 3.64 2.215 ;
 RECT 3.275 1.22 3.59 1.36 ;
 RECT 3.45 0.805 3.59 1.22 ;
 RECT 3.275 1.36 3.415 1.82 ;
 RECT 3.275 1.82 5.48 1.96 ;
 RECT 5.34 1.58 5.48 1.82 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.11 ;
 RECT 0.58 2.25 0.72 2.255 ;
 RECT 0.58 2.11 1.005 2.25 ;
 RECT 0.58 0.87 1.005 1.01 ;
 RECT 1.55 0.67 1.69 1.195 ;
 RECT 0.58 1.195 1.69 1.335 ;
 RECT 2.98 0.36 3.12 2.035 ;
 RECT 1.55 0.53 2.435 0.67 ;
 RECT 2.295 0.22 3.12 0.36 ;
 RECT 2.295 0.36 2.435 0.53 ;
 RECT 2.935 2.035 3.12 2.17 ;
 RECT 2.935 2.17 3.075 2.305 ;
 RECT 2.585 0.5 2.84 0.965 ;
 RECT 2.585 1.96 2.725 2.51 ;
 RECT 2.585 0.965 2.725 1.44 ;
 RECT 2.585 1.67 2.725 1.82 ;
 RECT 2.585 1.44 2.84 1.67 ;
 RECT 2.455 1.82 2.725 1.96 ;
 RECT 2.585 2.51 5.215 2.65 ;
 RECT 5.075 2.495 5.215 2.51 ;
 RECT 5.075 2.355 6.09 2.495 ;
 RECT 5.95 1.35 6.09 2.1 ;
 RECT 5.95 2.1 6.69 2.24 ;
 RECT 5.95 2.24 6.09 2.355 ;
 RECT 6.55 2.24 6.69 2.52 ;
 RECT 5.95 1.21 6.53 1.35 ;
 RECT 6.55 2.52 6.82 2.66 ;
 RECT 6.67 0.5 7.18 0.58 ;
 RECT 6.39 0.58 7.18 0.64 ;
 RECT 6.39 0.64 6.85 0.72 ;
 RECT 6.39 0.72 6.53 1.21 ;
 END
END DFFARX2

MACRO DFFASRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 12.16 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 12.16 2.96 ;
 RECT 5.345 2.635 5.605 2.8 ;
 RECT 2.095 1.95 2.265 2.8 ;
 RECT 1.26 1.93 1.4 2.8 ;
 RECT 6.365 2.38 6.505 2.8 ;
 RECT 9.155 2.15 9.295 2.8 ;
 RECT 10.275 2.06 10.415 2.8 ;
 RECT 11.8 1.52 11.94 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 12.16 0.08 ;
 RECT 8.63 0.08 8.885 1.01 ;
 RECT 4.605 0.08 4.84 0.37 ;
 RECT 1.26 0.08 1.4 1.055 ;
 RECT 1.96 0.08 2.19 0.39 ;
 RECT 11.915 0.08 12.055 0.87 ;
 RECT 10.295 0.08 10.435 0.725 ;
 RECT 0.28 0.08 0.42 0.775 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.275 1.475 1.575 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4 0.51 5.155 0.65 ;
 RECT 5.885 0.36 6.21 0.46 ;
 RECT 5.015 0.36 5.155 0.51 ;
 RECT 9.175 1.325 9.315 1.33 ;
 RECT 8.345 1.185 9.58 1.325 ;
 RECT 8.345 0.36 8.485 1.185 ;
 RECT 5.015 0.22 8.485 0.36 ;
 RECT 9.175 1.105 9.58 1.185 ;
 RECT 9.175 0.285 9.315 1.105 ;
 END
 ANTENNAGATEAREA 0.117 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.815 0.5 8.18 0.84 ;
 END
 ANTENNAGATEAREA 0.098 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.86 1.425 11 2.62 ;
 RECT 10.86 1.105 11.17 1.425 ;
 RECT 10.86 0.69 11 1.105 ;
 END
 ANTENNADIFFAREA 0.64 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.15 2.015 11.48 2.38 ;
 RECT 11.325 2.38 11.465 2.61 ;
 RECT 11.18 0.745 11.465 0.885 ;
 RECT 11.325 0.885 11.465 2.015 ;
 END
 ANTENNADIFFAREA 0.469 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.31 1.16 0.805 1.49 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 9.285 1.63 9.51 1.94 ;
 RECT 8.95 0.65 9.05 1.53 ;
 RECT 9.41 1.94 9.51 2.695 ;
 RECT 6.225 1.64 6.655 1.87 ;
 RECT 6.225 1.095 6.44 1.64 ;
 RECT 6.125 0.865 6.44 1.095 ;
 RECT 9.97 1.345 10.07 2.69 ;
 RECT 9.39 0.635 9.49 1.105 ;
 RECT 9.32 1.105 9.55 1.245 ;
 RECT 9.32 1.245 10.07 1.345 ;
 RECT 4.115 0.695 4.215 1.61 ;
 RECT 4.15 1.71 4.25 2.48 ;
 RECT 4.115 1.61 4.25 1.71 ;
 RECT 3.995 0.465 4.235 0.695 ;
 RECT 1.52 0.655 1.62 1.48 ;
 RECT 1.335 1.48 1.62 1.72 ;
 RECT 1.52 1.72 1.62 2.37 ;
 RECT 2.36 1.31 2.46 1.52 ;
 RECT 1.86 1.52 2.46 1.62 ;
 RECT 2.36 1.62 2.46 2.685 ;
 RECT 3.225 0.47 3.51 0.705 ;
 RECT 3.225 0.705 3.325 1.21 ;
 RECT 4.975 1.79 5.075 2.685 ;
 RECT 2.36 0.585 2.46 1.21 ;
 RECT 2.36 2.685 5.075 2.785 ;
 RECT 1.86 1.44 2.105 1.52 ;
 RECT 1.86 1.62 2.105 1.69 ;
 RECT 2.36 1.21 3.325 1.31 ;
 RECT 6.7 0.56 6.8 1.35 ;
 RECT 8.455 0.265 8.555 1.32 ;
 RECT 5.51 0.56 5.74 0.69 ;
 RECT 5.51 0.46 6.8 0.56 ;
 RECT 6.7 0.265 6.8 0.46 ;
 RECT 7.145 1.545 7.245 2.38 ;
 RECT 6.7 0.165 8.555 0.265 ;
 RECT 6.7 1.35 6.99 1.445 ;
 RECT 6.7 1.445 7.245 1.45 ;
 RECT 6.89 1.45 7.245 1.545 ;
 RECT 0.6 1.185 1.145 1.425 ;
 RECT 1.045 0.655 1.145 1.185 ;
 RECT 1.045 1.425 1.145 2.465 ;
 RECT 5.28 1.61 5.545 1.82 ;
 RECT 5.445 1.82 5.545 2.49 ;
 RECT 4.875 0.625 4.975 1.51 ;
 RECT 4.875 1.51 5.545 1.61 ;
 RECT 4.415 0.285 4.515 1.24 ;
 RECT 2.68 0.185 4.515 0.285 ;
 RECT 2.68 0.285 2.78 0.525 ;
 RECT 2.64 0.525 2.87 0.76 ;
 RECT 8.725 2.47 9.04 2.71 ;
 RECT 8.94 1.95 9.04 2.47 ;
 RECT 10.61 0.21 10.71 1.125 ;
 RECT 10.61 1.355 10.71 2.79 ;
 RECT 10.36 1.125 10.71 1.355 ;
 RECT 3.18 1.675 3.28 2.495 ;
 RECT 2.655 1.555 2.9 1.575 ;
 RECT 2.655 1.575 3.28 1.675 ;
 RECT 2.655 1.675 2.9 1.79 ;
 RECT 5.75 1.33 5.85 1.565 ;
 RECT 5.945 1.665 6.045 2.69 ;
 RECT 8.115 0.76 8.215 2.69 ;
 RECT 7.925 0.54 8.215 0.76 ;
 RECT 5.23 0.635 5.33 1.23 ;
 RECT 5.23 1.23 5.85 1.33 ;
 RECT 5.75 1.565 6.045 1.665 ;
 RECT 5.945 2.69 8.215 2.79 ;
 RECT 7.64 0.645 7.74 1.24 ;
 RECT 7.64 1.24 7.885 1.45 ;
 RECT 7.64 1.45 7.74 2.37 ;
 RECT 7.17 0.685 7.27 1.255 ;
 RECT 7.095 0.455 7.325 0.685 ;
 RECT 11.585 1.425 11.685 2.79 ;
 RECT 11.48 0.36 11.58 1.19 ;
 RECT 11.48 1.19 11.97 1.425 ;
 RECT 3.675 1.33 3.815 1.475 ;
 RECT 3.675 1.71 3.775 2.475 ;
 RECT 3.715 0.65 3.815 1.33 ;
 RECT 3.675 1.475 3.905 1.71 ;
 RECT 8.95 1.53 9.51 1.63 ;
 LAYER CO ;
 RECT 9.785 0.87 9.915 1 ;
 RECT 9.16 2.2 9.29 2.33 ;
 RECT 8.69 2.19 8.82 2.32 ;
 RECT 10.28 2.13 10.41 2.26 ;
 RECT 9.72 2.13 9.85 2.26 ;
 RECT 9.335 1.76 9.465 1.89 ;
 RECT 3.725 1.525 3.855 1.655 ;
 RECT 5.67 0.88 5.8 1.01 ;
 RECT 5.665 2.015 5.795 2.145 ;
 RECT 2.01 0.255 2.14 0.385 ;
 RECT 5.395 2.64 5.525 2.77 ;
 RECT 4.725 2.125 4.855 2.255 ;
 RECT 3.895 2.105 4.025 2.235 ;
 RECT 1.92 1.495 2.05 1.625 ;
 RECT 2.11 2.015 2.24 2.145 ;
 RECT 2.69 0.58 2.82 0.71 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 11.33 2.41 11.46 2.54 ;
 RECT 8.79 2.525 8.92 2.655 ;
 RECT 6.895 1.815 7.025 1.945 ;
 RECT 6.37 2.44 6.5 2.57 ;
 RECT 0.645 1.245 0.775 1.375 ;
 RECT 2.58 2.015 2.71 2.145 ;
 RECT 3.33 0.525 3.46 0.655 ;
 RECT 0.285 0.59 0.415 0.72 ;
 RECT 0.285 0.33 0.415 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 7.985 0.58 8.115 0.71 ;
 RECT 8.34 1.925 8.47 2.055 ;
 RECT 7.86 2.04 7.99 2.17 ;
 RECT 6.92 0.87 7.05 1 ;
 RECT 7.145 0.505 7.275 0.635 ;
 RECT 7.7 1.28 7.83 1.41 ;
 RECT 11.8 1.24 11.93 1.37 ;
 RECT 11.92 0.67 12.05 0.8 ;
 RECT 11.23 0.75 11.36 0.88 ;
 RECT 10.41 1.175 10.54 1.305 ;
 RECT 5.335 1.63 5.465 1.76 ;
 RECT 10.865 0.765 10.995 0.895 ;
 RECT 10.865 2.15 10.995 2.28 ;
 RECT 10.865 2.41 10.995 2.54 ;
 RECT 10.3 0.525 10.43 0.655 ;
 RECT 6.475 1.69 6.605 1.82 ;
 RECT 6.195 0.915 6.325 1.045 ;
 RECT 9.37 1.16 9.5 1.29 ;
 RECT 8.69 0.87 8.82 1 ;
 RECT 4.375 1.825 4.505 1.955 ;
 RECT 4.05 0.515 4.18 0.645 ;
 RECT 4.655 0.235 4.785 0.365 ;
 RECT 5.56 0.51 5.69 0.64 ;
 RECT 7.39 1.825 7.52 1.955 ;
 RECT 7.39 0.87 7.52 1 ;
 RECT 3.425 2.07 3.555 2.2 ;
 RECT 3.445 0.88 3.575 1.01 ;
 RECT 2.93 2.105 3.06 2.235 ;
 RECT 2.975 0.88 3.105 1.01 ;
 RECT 2.71 1.6 2.84 1.73 ;
 RECT 2.58 0.905 2.71 1.035 ;
 RECT 1.385 1.535 1.515 1.665 ;
 RECT 1.74 1.995 1.87 2.125 ;
 RECT 1.87 0.875 2 1.005 ;
 RECT 1.265 1.995 1.395 2.125 ;
 RECT 1.265 0.875 1.395 1.005 ;
 RECT 0.795 2.095 0.925 2.225 ;
 RECT 11.805 1.605 11.935 1.735 ;
 RECT 11.805 1.865 11.935 1.995 ;
 RECT 11.805 2.15 11.935 2.28 ;
 RECT 11.805 2.41 11.935 2.54 ;
 RECT 11.33 1.605 11.46 1.735 ;
 RECT 11.33 1.865 11.46 1.995 ;
 RECT 11.33 2.15 11.46 2.28 ;
 RECT 10.865 1.605 10.995 1.735 ;
 RECT 10.865 1.865 10.995 1.995 ;
 RECT 0.785 0.875 0.915 1.005 ;
 LAYER M1 ;
 RECT 3.26 0.52 3.86 0.66 ;
 RECT 3.72 0.66 3.86 0.79 ;
 RECT 5.295 0.505 5.74 0.645 ;
 RECT 3.72 0.79 5.435 0.93 ;
 RECT 5.295 0.645 5.435 0.79 ;
 RECT 5.66 1.015 6.395 1.05 ;
 RECT 5.66 1.05 5.8 1.185 ;
 RECT 5.66 1.325 5.8 2.01 ;
 RECT 5.05 1.185 5.8 1.325 ;
 RECT 5.6 0.875 6.395 1.015 ;
 RECT 5.61 2.01 5.865 2.15 ;
 RECT 5.05 1.325 5.19 1.52 ;
 RECT 3.655 1.52 5.19 1.66 ;
 RECT 3.825 2.12 4.925 2.24 ;
 RECT 3.825 2.1 4.095 2.12 ;
 RECT 3.89 2.24 4.925 2.26 ;
 RECT 10.575 0.36 10.715 0.885 ;
 RECT 9.78 0.885 10.715 1.025 ;
 RECT 11.605 0.56 11.745 1.235 ;
 RECT 10.575 0.22 11.41 0.36 ;
 RECT 11.27 0.42 11.745 0.56 ;
 RECT 11.27 0.36 11.41 0.42 ;
 RECT 9.78 1.025 9.92 1.475 ;
 RECT 7.695 1.475 9.92 1.615 ;
 RECT 9.715 1.615 9.855 2.325 ;
 RECT 9.78 0.8 9.92 0.885 ;
 RECT 7.695 1.21 7.835 1.475 ;
 RECT 11.605 1.235 11.995 1.375 ;
 RECT 2.575 2.43 6.145 2.435 ;
 RECT 6.005 1.35 6.145 2.1 ;
 RECT 6.005 2.24 6.145 2.295 ;
 RECT 5.065 2.295 6.145 2.43 ;
 RECT 2.575 2.435 5.205 2.57 ;
 RECT 2.575 0.84 2.825 1.035 ;
 RECT 2.575 1.78 2.715 2.43 ;
 RECT 2.685 0.51 2.825 0.84 ;
 RECT 2.575 1.035 2.715 1.55 ;
 RECT 2.575 1.55 2.845 1.78 ;
 RECT 7.505 2.24 7.645 2.52 ;
 RECT 6.56 0.5 7.35 0.64 ;
 RECT 6.005 2.1 7.645 2.24 ;
 RECT 6.56 0.64 6.7 1.21 ;
 RECT 6.005 1.21 6.7 1.35 ;
 RECT 7.505 2.52 9 2.66 ;
 RECT 1.54 0.67 1.68 1.195 ;
 RECT 0.98 1.195 1.68 1.335 ;
 RECT 0.98 1.01 1.12 1.195 ;
 RECT 0.98 1.335 1.12 1.945 ;
 RECT 0.79 2.085 0.93 2.305 ;
 RECT 0.715 0.87 1.12 1.01 ;
 RECT 0.79 1.945 1.12 2.085 ;
 RECT 1.54 0.53 2.49 0.67 ;
 RECT 2.97 0.36 3.11 1.175 ;
 RECT 2.35 0.22 3.11 0.36 ;
 RECT 2.985 1.27 3.125 2.1 ;
 RECT 2.35 0.36 2.49 0.53 ;
 RECT 2.86 2.1 3.125 2.24 ;
 RECT 2.97 1.175 3.125 1.27 ;
 RECT 7.81 2.22 8.825 2.36 ;
 RECT 7.81 2.035 8.04 2.22 ;
 RECT 8.685 2.14 8.825 2.22 ;
 RECT 8.685 2.36 8.825 2.375 ;
 RECT 3.265 1.82 5.47 1.96 ;
 RECT 3.265 1.22 3.58 1.36 ;
 RECT 3.44 0.805 3.58 1.22 ;
 RECT 3.35 1.96 3.63 2.215 ;
 RECT 5.33 1.56 5.47 1.82 ;
 RECT 3.265 1.36 3.405 1.82 ;
 RECT 1.865 0.825 2.005 1.475 ;
 RECT 1.735 1.63 1.875 2.2 ;
 RECT 1.735 1.475 2.125 1.63 ;
 RECT 7.315 1.82 9.575 1.895 ;
 RECT 7.385 1.755 9.575 1.82 ;
 RECT 9.995 1.92 10.135 2.505 ;
 RECT 9.435 2.505 10.135 2.645 ;
 RECT 9.435 1.895 9.575 2.505 ;
 RECT 7.315 1.895 7.595 1.96 ;
 RECT 7.385 0.805 7.525 1.755 ;
 RECT 8.29 1.895 8.52 2.06 ;
 RECT 10.23 1.31 10.37 1.78 ;
 RECT 10.23 1.17 10.61 1.31 ;
 RECT 9.995 1.78 10.37 1.92 ;
 RECT 6.405 1.685 7.125 1.825 ;
 RECT 6.825 1.825 7.125 1.95 ;
 RECT 6.915 1.005 7.125 1.685 ;
 RECT 6.845 0.865 7.125 1.005 ;
 END
END DFFASRX1

MACRO DFFASRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 12.8 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 12.8 2.96 ;
 RECT 5.345 2.635 5.605 2.8 ;
 RECT 2.095 1.95 2.265 2.8 ;
 RECT 11.33 1.56 11.47 2.8 ;
 RECT 9.155 2.15 9.295 2.8 ;
 RECT 10.275 2.06 10.415 2.8 ;
 RECT 12.28 1.52 12.42 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.26 1.93 1.4 2.8 ;
 RECT 6.365 2.38 6.505 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 12.8 0.08 ;
 RECT 8.625 0.08 8.88 1.005 ;
 RECT 4.605 0.08 4.84 0.37 ;
 RECT 1.26 0.08 1.4 1.055 ;
 RECT 1.96 0.08 2.19 0.39 ;
 RECT 12.555 0.08 12.695 0.87 ;
 RECT 11.535 0.08 11.675 0.885 ;
 RECT 10.295 0.08 10.435 0.725 ;
 RECT 0.28 0.08 0.42 0.775 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.275 1.475 1.575 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4 0.51 5.155 0.65 ;
 RECT 6.085 0.36 6.41 0.6 ;
 RECT 5.015 0.36 5.155 0.51 ;
 RECT 8.325 1.295 9.26 1.325 ;
 RECT 9.12 1.155 9.575 1.185 ;
 RECT 8.325 1.185 9.575 1.295 ;
 RECT 8.325 0.36 8.465 1.185 ;
 RECT 5.015 0.22 8.465 0.36 ;
 END
 ANTENNAGATEAREA 0.117 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.855 0.5 8.185 0.885 ;
 END
 ANTENNAGATEAREA 0.098 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.585 2.085 11 2.405 ;
 RECT 10.86 2.405 11 2.62 ;
 RECT 10.86 0.69 11 2.085 ;
 END
 ANTENNADIFFAREA 0.676 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.805 2.015 12.135 2.38 ;
 RECT 11.805 1.025 12.225 1.165 ;
 RECT 11.805 2.38 11.945 2.61 ;
 RECT 12.085 0.675 12.225 1.025 ;
 RECT 11.805 1.165 11.945 2.015 ;
 END
 ANTENNADIFFAREA 0.568 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.31 1.16 0.805 1.49 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 8.455 0.265 8.555 1.32 ;
 RECT 5.715 0.56 5.945 0.69 ;
 RECT 5.715 0.46 6.8 0.56 ;
 RECT 6.7 0.265 6.8 0.46 ;
 RECT 7.145 1.545 7.245 2.38 ;
 RECT 6.7 0.165 8.555 0.265 ;
 RECT 6.7 1.35 6.99 1.445 ;
 RECT 6.7 1.445 7.245 1.45 ;
 RECT 6.89 1.45 7.245 1.545 ;
 RECT 0.6 1.185 1.145 1.425 ;
 RECT 1.045 0.655 1.145 1.185 ;
 RECT 1.045 1.425 1.145 2.465 ;
 RECT 8.725 2.47 9.04 2.71 ;
 RECT 8.94 1.95 9.04 2.47 ;
 RECT 11.48 1.19 12.44 1.29 ;
 RECT 11.87 0.345 11.97 1.19 ;
 RECT 12.065 1.29 12.165 2.79 ;
 RECT 11.48 1.29 11.69 1.425 ;
 RECT 11.59 1.425 11.69 2.79 ;
 RECT 12.34 0.36 12.44 1.19 ;
 RECT 10.61 0.21 10.71 1.125 ;
 RECT 10.36 1.125 10.71 1.19 ;
 RECT 10.61 1.355 10.71 2.79 ;
 RECT 10.36 1.29 10.71 1.355 ;
 RECT 10.36 1.19 11.215 1.29 ;
 RECT 11.115 0.21 11.215 1.19 ;
 RECT 11.115 1.29 11.215 2.79 ;
 RECT 8.95 1.53 9.51 1.63 ;
 RECT 9.285 1.63 9.51 1.94 ;
 RECT 8.95 0.65 9.05 1.53 ;
 RECT 9.41 1.94 9.51 2.695 ;
 RECT 6.235 1.64 6.655 1.87 ;
 RECT 6.235 1.095 6.44 1.64 ;
 RECT 6.125 0.865 6.44 1.095 ;
 RECT 9.97 1.345 10.07 2.69 ;
 RECT 9.39 0.635 9.49 1.105 ;
 RECT 9.32 1.105 9.55 1.245 ;
 RECT 9.32 1.245 10.07 1.345 ;
 RECT 4.115 0.695 4.215 1.61 ;
 RECT 4.15 1.71 4.25 2.48 ;
 RECT 4.115 1.61 4.25 1.71 ;
 RECT 3.995 0.465 4.235 0.695 ;
 RECT 5.75 1.33 5.85 1.565 ;
 RECT 5.955 1.665 6.055 2.69 ;
 RECT 8.115 0.745 8.215 2.69 ;
 RECT 5.23 0.635 5.33 1.23 ;
 RECT 5.23 1.23 5.85 1.33 ;
 RECT 5.75 1.565 6.055 1.665 ;
 RECT 5.955 2.69 8.215 2.79 ;
 RECT 7.92 0.525 8.215 0.745 ;
 RECT 7.64 0.645 7.74 1.24 ;
 RECT 7.64 1.24 7.885 1.45 ;
 RECT 7.64 1.45 7.74 2.37 ;
 RECT 7.17 0.685 7.27 1.255 ;
 RECT 7.095 0.455 7.325 0.685 ;
 RECT 5.28 1.61 5.545 1.82 ;
 RECT 5.445 1.82 5.545 2.49 ;
 RECT 4.875 0.625 4.975 1.51 ;
 RECT 4.875 1.51 5.545 1.61 ;
 RECT 3.675 1.33 3.815 1.475 ;
 RECT 3.675 1.71 3.775 2.475 ;
 RECT 3.715 0.65 3.815 1.33 ;
 RECT 3.675 1.475 3.905 1.71 ;
 RECT 4.415 0.285 4.515 1.24 ;
 RECT 2.68 0.185 4.515 0.285 ;
 RECT 2.68 0.285 2.78 0.525 ;
 RECT 2.64 0.525 2.87 0.76 ;
 RECT 3.18 1.675 3.28 2.495 ;
 RECT 2.655 1.555 2.9 1.575 ;
 RECT 2.655 1.675 2.9 1.79 ;
 RECT 2.655 1.575 3.28 1.675 ;
 RECT 1.52 0.655 1.62 1.48 ;
 RECT 1.335 1.48 1.62 1.72 ;
 RECT 1.52 1.72 1.62 2.37 ;
 RECT 2.36 1.31 2.46 1.52 ;
 RECT 1.86 1.52 2.46 1.62 ;
 RECT 2.36 1.62 2.46 2.685 ;
 RECT 3.225 0.47 3.51 0.705 ;
 RECT 3.225 0.705 3.325 1.21 ;
 RECT 4.975 1.79 5.075 2.685 ;
 RECT 2.36 2.685 5.075 2.785 ;
 RECT 2.36 0.585 2.46 1.21 ;
 RECT 1.86 1.44 2.105 1.52 ;
 RECT 1.86 1.62 2.105 1.69 ;
 RECT 2.36 1.21 3.325 1.31 ;
 RECT 6.7 0.56 6.8 1.35 ;
 LAYER CO ;
 RECT 0.645 1.245 0.775 1.375 ;
 RECT 2.58 2.015 2.71 2.145 ;
 RECT 3.33 0.525 3.46 0.655 ;
 RECT 0.285 0.59 0.415 0.72 ;
 RECT 0.285 0.33 0.415 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 4.05 0.515 4.18 0.645 ;
 RECT 7.98 0.575 8.11 0.705 ;
 RECT 7.39 1.825 7.52 1.955 ;
 RECT 8.34 1.925 8.47 2.055 ;
 RECT 7.86 2.04 7.99 2.17 ;
 RECT 6.92 0.87 7.05 1 ;
 RECT 7.145 0.505 7.275 0.635 ;
 RECT 7.7 1.28 7.83 1.41 ;
 RECT 9.785 0.87 9.915 1 ;
 RECT 9.16 2.2 9.29 2.33 ;
 RECT 8.69 2.19 8.82 2.32 ;
 RECT 10.28 2.13 10.41 2.26 ;
 RECT 9.72 2.13 9.85 2.26 ;
 RECT 9.335 1.76 9.465 1.89 ;
 RECT 5.335 1.63 5.465 1.76 ;
 RECT 3.725 1.525 3.855 1.655 ;
 RECT 5.67 0.88 5.8 1.01 ;
 RECT 5.665 2.015 5.795 2.145 ;
 RECT 2.01 0.255 2.14 0.385 ;
 RECT 5.395 2.64 5.525 2.77 ;
 RECT 4.725 2.125 4.855 2.255 ;
 RECT 11.54 0.665 11.67 0.795 ;
 RECT 11.335 1.61 11.465 1.74 ;
 RECT 11.335 1.87 11.465 2 ;
 RECT 11.335 2.155 11.465 2.285 ;
 RECT 7.39 0.87 7.52 1 ;
 RECT 11.335 2.415 11.465 2.545 ;
 RECT 4.375 1.825 4.505 1.955 ;
 RECT 3.895 2.105 4.025 2.235 ;
 RECT 1.92 1.495 2.05 1.625 ;
 RECT 2.11 2.015 2.24 2.145 ;
 RECT 2.69 0.58 2.82 0.71 ;
 RECT 3.425 2.07 3.555 2.2 ;
 RECT 3.445 0.88 3.575 1.01 ;
 RECT 2.93 2.105 3.06 2.235 ;
 RECT 2.975 0.88 3.105 1.01 ;
 RECT 2.71 1.6 2.84 1.73 ;
 RECT 2.58 0.905 2.71 1.035 ;
 RECT 1.385 1.535 1.515 1.665 ;
 RECT 1.74 1.995 1.87 2.125 ;
 RECT 1.87 0.875 2 1.005 ;
 RECT 1.265 1.995 1.395 2.125 ;
 RECT 1.265 0.875 1.395 1.005 ;
 RECT 0.795 2.095 0.925 2.225 ;
 RECT 12.285 1.605 12.415 1.735 ;
 RECT 12.285 1.865 12.415 1.995 ;
 RECT 12.285 2.15 12.415 2.28 ;
 RECT 12.285 2.41 12.415 2.54 ;
 RECT 11.81 1.605 11.94 1.735 ;
 RECT 11.81 1.865 11.94 1.995 ;
 RECT 11.81 2.15 11.94 2.28 ;
 RECT 10.865 1.605 10.995 1.735 ;
 RECT 0.785 0.875 0.915 1.005 ;
 RECT 11.81 2.41 11.94 2.54 ;
 RECT 10.865 1.865 10.995 1.995 ;
 RECT 8.79 2.525 8.92 2.655 ;
 RECT 6.895 1.815 7.025 1.945 ;
 RECT 6.37 2.44 6.5 2.57 ;
 RECT 11.52 1.24 11.65 1.37 ;
 RECT 12.56 0.67 12.69 0.8 ;
 RECT 12.09 0.75 12.22 0.88 ;
 RECT 10.41 1.175 10.54 1.305 ;
 RECT 10.865 0.765 10.995 0.895 ;
 RECT 10.865 2.15 10.995 2.28 ;
 RECT 10.865 2.41 10.995 2.54 ;
 RECT 10.3 0.525 10.43 0.655 ;
 RECT 6.475 1.69 6.605 1.82 ;
 RECT 6.195 0.915 6.325 1.045 ;
 RECT 9.37 1.16 9.5 1.29 ;
 RECT 8.7 0.87 8.83 1 ;
 RECT 4.655 0.235 4.785 0.365 ;
 RECT 5.765 0.51 5.895 0.64 ;
 LAYER M1 ;
 RECT 3.825 2.12 4.925 2.24 ;
 RECT 3.825 2.1 4.095 2.12 ;
 RECT 3.89 2.24 4.925 2.26 ;
 RECT 5.66 1.325 5.8 2.01 ;
 RECT 5.66 1.05 5.8 1.185 ;
 RECT 5.05 1.185 5.8 1.325 ;
 RECT 5.66 1.015 6.395 1.05 ;
 RECT 3.655 1.52 5.19 1.66 ;
 RECT 5.05 1.325 5.19 1.52 ;
 RECT 5.61 2.01 5.865 2.15 ;
 RECT 5.6 0.875 6.395 1.015 ;
 RECT 3.26 0.52 3.86 0.66 ;
 RECT 3.72 0.66 3.86 0.79 ;
 RECT 3.72 0.79 5.435 0.93 ;
 RECT 5.295 0.505 5.945 0.645 ;
 RECT 5.295 0.645 5.435 0.79 ;
 RECT 7.695 1.21 7.835 1.475 ;
 RECT 9.78 0.865 10.715 1.005 ;
 RECT 10.575 0.525 10.715 0.865 ;
 RECT 11.165 0.525 11.305 1.1 ;
 RECT 10.575 0.385 11.305 0.525 ;
 RECT 7.695 1.475 9.92 1.615 ;
 RECT 9.78 1.005 9.92 1.475 ;
 RECT 9.78 0.8 9.92 0.865 ;
 RECT 9.715 1.615 9.855 2.325 ;
 RECT 11.515 1.24 11.655 1.42 ;
 RECT 11.165 1.1 11.655 1.24 ;
 RECT 7.81 2.22 8.825 2.36 ;
 RECT 7.81 2.035 8.04 2.22 ;
 RECT 8.685 2.14 8.825 2.22 ;
 RECT 8.685 2.36 8.825 2.375 ;
 RECT 2.575 2.43 6.145 2.435 ;
 RECT 6.005 1.35 6.145 2.1 ;
 RECT 6.005 2.24 6.145 2.295 ;
 RECT 5.065 2.295 6.145 2.43 ;
 RECT 2.575 2.435 5.205 2.57 ;
 RECT 2.575 0.84 2.825 1.035 ;
 RECT 2.575 1.78 2.715 2.43 ;
 RECT 2.685 0.51 2.825 0.84 ;
 RECT 2.575 1.035 2.715 1.55 ;
 RECT 2.575 1.55 2.845 1.78 ;
 RECT 7.505 2.24 7.645 2.52 ;
 RECT 6.56 0.5 7.35 0.64 ;
 RECT 6.56 0.64 6.7 1.21 ;
 RECT 6.005 1.21 6.7 1.35 ;
 RECT 6.005 2.1 7.645 2.24 ;
 RECT 7.505 2.52 9 2.66 ;
 RECT 1.735 1.63 1.875 2.2 ;
 RECT 1.865 0.825 2.005 1.475 ;
 RECT 1.735 1.475 2.125 1.63 ;
 RECT 0.98 1.01 1.12 1.195 ;
 RECT 0.98 1.335 1.12 1.945 ;
 RECT 0.79 2.085 0.93 2.305 ;
 RECT 0.715 0.87 1.12 1.01 ;
 RECT 0.79 1.945 1.12 2.085 ;
 RECT 1.54 0.67 1.68 1.195 ;
 RECT 0.98 1.195 1.68 1.335 ;
 RECT 1.54 0.53 2.49 0.67 ;
 RECT 2.97 0.36 3.11 1.175 ;
 RECT 2.35 0.22 3.11 0.36 ;
 RECT 2.985 1.27 3.125 2.1 ;
 RECT 2.35 0.36 2.49 0.53 ;
 RECT 2.86 2.1 3.125 2.24 ;
 RECT 2.97 1.175 3.125 1.27 ;
 RECT 3.265 1.82 5.47 1.96 ;
 RECT 3.265 1.22 3.58 1.36 ;
 RECT 3.44 0.805 3.58 1.22 ;
 RECT 3.35 1.96 3.63 2.215 ;
 RECT 5.33 1.56 5.47 1.82 ;
 RECT 3.265 1.36 3.405 1.82 ;
 RECT 6.405 1.685 7.125 1.825 ;
 RECT 6.825 1.825 7.125 1.95 ;
 RECT 6.915 1.005 7.125 1.685 ;
 RECT 6.845 0.865 7.125 1.005 ;
 RECT 7.315 1.895 7.595 1.96 ;
 RECT 7.385 0.805 7.525 1.755 ;
 RECT 7.315 1.82 9.575 1.895 ;
 RECT 7.385 1.755 9.575 1.82 ;
 RECT 9.995 1.92 10.135 2.505 ;
 RECT 9.435 2.505 10.135 2.645 ;
 RECT 9.435 1.895 9.575 2.505 ;
 RECT 8.29 1.895 8.52 2.06 ;
 RECT 10.23 1.31 10.37 1.78 ;
 RECT 9.995 1.78 10.37 1.92 ;
 RECT 10.23 1.17 10.61 1.31 ;
 END
END DFFASRX2

MACRO DFFASX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.88 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.88 2.96 ;
 RECT 4.495 2.635 4.755 2.8 ;
 RECT 2.155 2.36 2.405 2.8 ;
 RECT 0.54 1.76 0.68 2.8 ;
 RECT 8.26 2.055 8.4 2.8 ;
 RECT 9.935 1.48 10.075 2.8 ;
 RECT 5.485 2.38 5.625 2.8 ;
 RECT 1.5 2.06 1.64 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.88 0.08 ;
 RECT 1.455 0.84 1.685 0.98 ;
 RECT 2.075 0.08 2.305 0.385 ;
 RECT 10.03 0.08 10.17 0.76 ;
 RECT 4.465 0.08 4.605 0.38 ;
 RECT 0.54 0.08 0.68 0.795 ;
 RECT 7.775 0.08 7.915 1.07 ;
 RECT 1.5 0.08 1.64 0.84 ;
 END
 END VSS

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.025 0.435 7.375 0.8 ;
 END
 ANTENNAGATEAREA 0.088 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.27 0.52 9.605 0.77 ;
 RECT 9.38 0.77 9.52 2.51 ;
 END
 ANTENNADIFFAREA 0.611 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.28 2.065 10.555 2.385 ;
 RECT 10.415 0.77 10.64 0.91 ;
 RECT 10.5 0.555 10.64 0.77 ;
 RECT 10.415 2.385 10.555 2.52 ;
 RECT 10.415 0.91 10.555 2.065 ;
 END
 ANTENNADIFFAREA 0.469 ;
 END Q

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.845 1.48 2.21 1.805 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 1.495 1.49 1.88 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 3.42 1.77 3.52 2.495 ;
 RECT 2.815 1.77 3.06 1.92 ;
 RECT 2.815 1.67 3.52 1.77 ;
 RECT 1.76 0.625 1.86 1.5 ;
 RECT 1.76 1.5 2.03 1.74 ;
 RECT 1.76 1.74 1.86 2.39 ;
 RECT 4.575 0.625 4.675 1.58 ;
 RECT 4.705 1.82 4.805 2.39 ;
 RECT 4.575 1.58 4.815 1.82 ;
 RECT 5.46 1.64 5.84 1.87 ;
 RECT 5.46 1.095 5.625 1.64 ;
 RECT 5.355 0.865 5.625 1.095 ;
 RECT 5.805 0.265 5.905 0.575 ;
 RECT 5.155 0.575 5.905 0.675 ;
 RECT 5.805 0.675 5.905 1.35 ;
 RECT 6.25 1.545 6.35 2.415 ;
 RECT 7.56 0.265 7.66 1.32 ;
 RECT 5.155 0.455 5.385 0.575 ;
 RECT 5.155 0.675 5.385 0.685 ;
 RECT 5.995 1.45 6.35 1.545 ;
 RECT 5.805 0.165 7.66 0.265 ;
 RECT 5.805 1.35 6.095 1.445 ;
 RECT 5.805 1.445 6.35 1.45 ;
 RECT 2.535 1.69 2.635 2.685 ;
 RECT 2.535 1.355 2.635 1.44 ;
 RECT 3.465 0.705 3.565 1.255 ;
 RECT 4.22 1.795 4.32 2.685 ;
 RECT 3.465 0.47 3.75 0.705 ;
 RECT 2.535 2.685 4.32 2.785 ;
 RECT 2.535 1.255 3.565 1.355 ;
 RECT 2.285 1.44 2.635 1.69 ;
 RECT 2.6 0.515 2.7 1.255 ;
 RECT 8.39 1.63 8.615 1.94 ;
 RECT 8.515 1.94 8.615 2.66 ;
 RECT 8.03 0.65 8.13 1.53 ;
 RECT 8.03 1.53 8.615 1.63 ;
 RECT 10.285 0.215 10.385 1.035 ;
 RECT 10.195 1.27 10.295 2.79 ;
 RECT 10.035 1.035 10.385 1.27 ;
 RECT 9.645 0.145 9.745 1.18 ;
 RECT 9.645 1.28 9.745 2.79 ;
 RECT 9.065 1.18 9.745 1.28 ;
 RECT 9.065 1.28 9.275 1.415 ;
 RECT 7.83 2.47 8.145 2.71 ;
 RECT 8.045 1.88 8.145 2.47 ;
 RECT 6.745 0.645 6.845 1.24 ;
 RECT 6.745 1.24 6.99 1.45 ;
 RECT 6.745 1.45 6.845 2.37 ;
 RECT 6.275 0.685 6.375 1.23 ;
 RECT 6.2 0.455 6.43 0.685 ;
 RECT 2.92 0.285 3.02 0.5 ;
 RECT 2.92 0.185 4.35 0.285 ;
 RECT 4.25 0.285 4.35 1.24 ;
 RECT 2.88 0.5 3.11 0.735 ;
 RECT 3.915 1.43 4.015 1.475 ;
 RECT 3.915 1.71 4.015 2.505 ;
 RECT 3.935 0.65 4.035 1.33 ;
 RECT 3.915 1.33 4.035 1.43 ;
 RECT 3.785 1.475 4.015 1.71 ;
 RECT 1.285 0.195 1.385 1.5 ;
 RECT 1.285 1.74 1.385 2.485 ;
 RECT 1.27 1.5 1.49 1.74 ;
 RECT 7.22 0.715 7.32 2.69 ;
 RECT 5.18 2.69 7.32 2.79 ;
 RECT 5.18 1.375 5.28 2.69 ;
 RECT 4.875 1.275 5.28 1.375 ;
 RECT 7.1 0.475 7.32 0.715 ;
 RECT 4.875 0.635 4.975 1.275 ;
 LAYER CO ;
 RECT 1.505 0.845 1.635 0.975 ;
 RECT 1.035 2.11 1.165 2.24 ;
 RECT 0.545 2.365 0.675 2.495 ;
 RECT 1.98 2.015 2.11 2.145 ;
 RECT 0.545 2.105 0.675 2.235 ;
 RECT 2.11 0.855 2.24 0.985 ;
 RECT 7.895 2.525 8.025 2.655 ;
 RECT 10.42 2.05 10.55 2.18 ;
 RECT 10.42 2.31 10.55 2.44 ;
 RECT 9.94 1.53 10.07 1.66 ;
 RECT 9.94 1.79 10.07 1.92 ;
 RECT 10.505 0.625 10.635 0.755 ;
 RECT 10.035 0.56 10.165 0.69 ;
 RECT 2.93 0.555 3.06 0.685 ;
 RECT 5.205 0.505 5.335 0.635 ;
 RECT 6.495 1.9 6.625 2.03 ;
 RECT 6.495 0.87 6.625 1 ;
 RECT 6.805 1.28 6.935 1.41 ;
 RECT 8.25 0.87 8.38 1 ;
 RECT 8.265 2.115 8.395 2.245 ;
 RECT 7.15 0.53 7.28 0.66 ;
 RECT 4.645 1.63 4.775 1.76 ;
 RECT 3.835 1.525 3.965 1.655 ;
 RECT 4.93 2.015 5.06 2.145 ;
 RECT 7.78 0.87 7.91 1 ;
 RECT 1.505 2.13 1.635 2.26 ;
 RECT 9.94 2.05 10.07 2.18 ;
 RECT 9.94 2.31 10.07 2.44 ;
 RECT 9.385 2.05 9.515 2.18 ;
 RECT 9.385 2.31 9.515 2.44 ;
 RECT 3.685 0.88 3.815 1.01 ;
 RECT 3.17 2.105 3.3 2.235 ;
 RECT 3.215 0.88 3.345 1.01 ;
 RECT 2.82 0.905 2.95 1.035 ;
 RECT 9.385 0.585 9.515 0.715 ;
 RECT 2.885 1.725 3.015 1.855 ;
 RECT 7.445 1.965 7.575 2.095 ;
 RECT 6.965 1.965 7.095 2.095 ;
 RECT 6.025 0.87 6.155 1 ;
 RECT 6.25 0.505 6.38 0.635 ;
 RECT 1.86 1.555 1.99 1.685 ;
 RECT 1.035 0.845 1.165 0.975 ;
 RECT 7.795 2.11 7.925 2.24 ;
 RECT 9.385 1.79 9.515 1.92 ;
 RECT 8.825 2.13 8.955 2.26 ;
 RECT 8.44 1.76 8.57 1.89 ;
 RECT 6 1.815 6.13 1.945 ;
 RECT 5.49 2.44 5.62 2.57 ;
 RECT 10.075 1.085 10.205 1.215 ;
 RECT 5.66 1.69 5.79 1.82 ;
 RECT 5.42 0.915 5.55 1.045 ;
 RECT 2.355 1.495 2.485 1.625 ;
 RECT 2.225 2.365 2.355 2.495 ;
 RECT 3.665 2.07 3.795 2.2 ;
 RECT 5.095 0.88 5.225 1.01 ;
 RECT 9.385 1.53 9.515 1.66 ;
 RECT 4.47 0.2 4.6 0.33 ;
 RECT 0.545 0.61 0.675 0.74 ;
 RECT 0.545 0.35 0.675 0.48 ;
 RECT 2.755 2.23 2.885 2.36 ;
 RECT 3.57 0.525 3.7 0.655 ;
 RECT 2.125 0.25 2.255 0.38 ;
 RECT 4.545 2.64 4.675 2.77 ;
 RECT 1.32 1.555 1.45 1.685 ;
 RECT 9.105 1.23 9.235 1.36 ;
 RECT 10.42 1.53 10.55 1.66 ;
 RECT 10.42 1.79 10.55 1.92 ;
 RECT 0.545 1.845 0.675 1.975 ;
 LAYER M1 ;
 RECT 2.105 0.805 2.245 1.125 ;
 RECT 2.105 1.125 2.49 1.265 ;
 RECT 2.35 1.265 2.49 2.01 ;
 RECT 1.91 2.01 2.49 2.15 ;
 RECT 6.96 2.1 7.145 2.24 ;
 RECT 7.79 2.03 7.93 2.24 ;
 RECT 6.915 1.96 7.145 2.1 ;
 RECT 6.96 2.24 7.93 2.38 ;
 RECT 6.8 1.21 6.94 1.395 ;
 RECT 8.82 0.38 8.96 0.865 ;
 RECT 8.2 0.865 8.96 1.005 ;
 RECT 8.82 1.005 8.96 1.395 ;
 RECT 6.8 1.395 8.96 1.535 ;
 RECT 8.82 1.535 8.96 2.32 ;
 RECT 9.75 0.38 9.89 1.15 ;
 RECT 8.82 0.24 9.89 0.38 ;
 RECT 10.07 1.02 10.21 1.15 ;
 RECT 9.75 1.15 10.21 1.29 ;
 RECT 0.82 1.26 0.96 2.105 ;
 RECT 0.82 0.98 0.96 1.12 ;
 RECT 0.82 2.105 1.235 2.245 ;
 RECT 0.82 0.84 1.24 0.98 ;
 RECT 0.82 1.12 1.965 1.26 ;
 RECT 1.825 0.665 1.965 1.12 ;
 RECT 3.21 0.36 3.35 0.875 ;
 RECT 3.225 1.015 3.365 2.035 ;
 RECT 2.53 0.36 2.67 0.525 ;
 RECT 3.165 2.035 3.365 2.305 ;
 RECT 3.165 0.875 3.42 1.015 ;
 RECT 1.825 0.525 2.67 0.665 ;
 RECT 2.53 0.22 3.35 0.36 ;
 RECT 5.65 1.685 6.16 1.81 ;
 RECT 5.65 1.81 6.2 1.825 ;
 RECT 6.02 0.78 6.16 1.685 ;
 RECT 5.65 1.615 5.79 1.685 ;
 RECT 5.65 1.825 5.79 1.895 ;
 RECT 5.93 1.825 6.2 1.95 ;
 RECT 6.49 1.815 6.7 1.895 ;
 RECT 6.49 0.805 6.63 1.675 ;
 RECT 7.395 1.815 7.625 2.1 ;
 RECT 6.42 1.895 6.7 2.035 ;
 RECT 6.49 1.675 8.68 1.815 ;
 RECT 9.1 1.18 9.24 2.505 ;
 RECT 8.38 1.815 8.68 1.915 ;
 RECT 8.54 1.915 8.68 2.505 ;
 RECT 8.54 2.505 9.24 2.645 ;
 RECT 5.205 1.36 5.345 2.1 ;
 RECT 5.205 2.24 5.345 2.355 ;
 RECT 4.13 2.355 5.345 2.495 ;
 RECT 2.75 2.515 4.27 2.655 ;
 RECT 2.815 0.735 2.955 1.72 ;
 RECT 2.815 1.72 3.065 1.775 ;
 RECT 2.75 1.775 3.065 1.86 ;
 RECT 2.75 1.86 2.955 2.005 ;
 RECT 2.75 2.005 2.89 2.515 ;
 RECT 2.925 0.505 3.065 0.535 ;
 RECT 4.13 2.495 4.27 2.515 ;
 RECT 2.815 0.535 3.065 0.735 ;
 RECT 6.135 2.24 6.75 2.32 ;
 RECT 5.205 2.185 6.75 2.24 ;
 RECT 6.61 2.32 6.75 2.52 ;
 RECT 5.205 2.1 6.275 2.18 ;
 RECT 5.205 2.18 6.745 2.185 ;
 RECT 5.74 0.5 6.455 0.64 ;
 RECT 5.74 0.64 5.88 1.22 ;
 RECT 5.205 1.22 5.88 1.36 ;
 RECT 6.61 2.52 8.105 2.66 ;
 RECT 4.925 1.04 5.6 1.05 ;
 RECT 4.36 0.91 5.6 1.04 ;
 RECT 4.36 0.9 5.23 0.91 ;
 RECT 4.925 1.08 5.065 2.2 ;
 RECT 4.925 1.05 5.23 1.08 ;
 RECT 3.785 1.52 4.5 1.66 ;
 RECT 5.09 0.81 5.23 0.9 ;
 RECT 4.36 1.04 4.5 1.52 ;
 RECT 3.5 0.52 5.41 0.66 ;
 RECT 5.125 0.47 5.41 0.52 ;
 RECT 3.505 1.805 4.78 1.945 ;
 RECT 3.505 1.945 3.87 1.96 ;
 RECT 3.505 1.22 3.82 1.36 ;
 RECT 3.68 0.805 3.82 1.22 ;
 RECT 3.59 1.96 3.87 2.215 ;
 RECT 3.505 1.36 3.645 1.805 ;
 RECT 4.64 1.56 4.78 1.805 ;
 END
END DFFASX1

MACRO DFFASX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.84 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.84 2.96 ;
 RECT 2.155 2.42 2.405 2.8 ;
 RECT 4.495 2.635 4.755 2.8 ;
 RECT 9.38 1.48 9.52 2.8 ;
 RECT 5.485 2.38 5.625 2.8 ;
 RECT 10.415 1.48 10.555 2.8 ;
 RECT 11.36 1.48 11.5 2.8 ;
 RECT 1.5 2.16 1.64 2.8 ;
 RECT 0.54 1.76 0.68 2.8 ;
 RECT 8.26 2.055 8.4 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.84 0.08 ;
 RECT 1.5 0.08 1.64 1.05 ;
 RECT 10.285 0.08 10.565 0.245 ;
 RECT 2.075 0.08 2.305 0.385 ;
 RECT 4.465 0.08 4.605 0.38 ;
 RECT 9.315 0.08 9.455 0.655 ;
 RECT 0.54 0.08 0.68 0.795 ;
 RECT 7.775 0.08 7.915 1.07 ;
 RECT 11.355 0.08 11.495 0.85 ;
 END
 END VSS

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.04 0.475 7.635 0.795 ;
 END
 ANTENNAGATEAREA 0.088 ;
 END SETB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.64 1.48 2.04 1.88 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 1.16 0.875 1.4 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.8 2.11 10.04 2.36 ;
 RECT 9.88 2.36 10.02 2.51 ;
 RECT 9.88 0.675 10.02 2.11 ;
 END
 ANTENNADIFFAREA 0.714 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.76 1.79 11.025 2.04 ;
 RECT 10.885 2.04 11.025 2.51 ;
 RECT 10.885 0.58 11.025 1.79 ;
 END
 ANTENNADIFFAREA 0.622 ;
 END Q

 OBS
 LAYER PO ;
 RECT 2.92 0.285 3.02 0.5 ;
 RECT 2.92 0.185 4.35 0.285 ;
 RECT 4.25 0.285 4.35 1.24 ;
 RECT 2.88 0.5 3.11 0.735 ;
 RECT 5.525 1.095 5.625 1.64 ;
 RECT 5.525 1.64 5.84 1.87 ;
 RECT 5.355 0.865 5.625 1.095 ;
 RECT 9.065 1.18 10.295 1.28 ;
 RECT 9.065 1.28 9.275 1.415 ;
 RECT 9.645 0.145 9.745 1.18 ;
 RECT 9.645 1.28 9.745 2.79 ;
 RECT 10.195 1.28 10.295 2.79 ;
 RECT 10.135 0.14 10.235 1.18 ;
 RECT 2.285 1.44 2.635 1.69 ;
 RECT 2.535 1.355 2.635 1.44 ;
 RECT 2.535 1.69 2.635 2.685 ;
 RECT 3.465 0.705 3.565 1.255 ;
 RECT 4.22 1.795 4.32 2.685 ;
 RECT 3.465 0.47 3.75 0.705 ;
 RECT 2.535 2.685 4.32 2.785 ;
 RECT 2.535 1.255 3.565 1.355 ;
 RECT 2.6 0.515 2.7 1.255 ;
 RECT 5.155 0.575 5.905 0.675 ;
 RECT 5.805 0.675 5.905 1.35 ;
 RECT 7.56 0.265 7.66 1.32 ;
 RECT 5.805 0.265 5.905 0.575 ;
 RECT 5.155 0.455 5.385 0.575 ;
 RECT 5.155 0.675 5.385 0.685 ;
 RECT 6.25 1.545 6.35 2.435 ;
 RECT 5.805 0.165 7.66 0.265 ;
 RECT 5.805 1.35 6.095 1.445 ;
 RECT 5.805 1.445 6.35 1.45 ;
 RECT 5.995 1.45 6.35 1.545 ;
 RECT 8.03 1.53 8.615 1.63 ;
 RECT 8.39 1.63 8.615 1.94 ;
 RECT 8.03 0.65 8.13 1.53 ;
 RECT 8.515 1.94 8.615 2.56 ;
 RECT 4.575 0.625 4.675 1.58 ;
 RECT 4.705 1.82 4.805 2.39 ;
 RECT 4.575 1.58 4.815 1.82 ;
 RECT 3.42 1.77 3.52 2.495 ;
 RECT 2.815 1.77 3.06 1.92 ;
 RECT 2.815 1.67 3.52 1.77 ;
 RECT 1.285 0.195 1.385 1.23 ;
 RECT 1.285 1.33 1.385 2.59 ;
 RECT 0.64 1.175 0.87 1.23 ;
 RECT 0.64 1.33 0.87 1.385 ;
 RECT 0.64 1.23 1.385 1.33 ;
 RECT 3.915 1.43 4.015 1.475 ;
 RECT 3.915 1.71 4.015 2.505 ;
 RECT 3.935 0.65 4.035 1.33 ;
 RECT 3.915 1.33 4.035 1.43 ;
 RECT 3.785 1.475 4.015 1.71 ;
 RECT 7.83 2.47 8.145 2.71 ;
 RECT 8.045 1.88 8.145 2.47 ;
 RECT 6.745 0.645 6.845 1.24 ;
 RECT 6.745 1.24 6.99 1.45 ;
 RECT 6.745 1.45 6.845 2.37 ;
 RECT 6.275 0.685 6.375 1.23 ;
 RECT 6.2 0.455 6.43 0.685 ;
 RECT 5.195 1.375 5.295 2.69 ;
 RECT 4.875 1.275 5.295 1.375 ;
 RECT 5.195 2.69 7.32 2.79 ;
 RECT 7.22 0.755 7.32 2.69 ;
 RECT 7.08 0.525 7.32 0.755 ;
 RECT 4.875 0.635 4.975 1.275 ;
 RECT 1.76 0.675 1.86 1.5 ;
 RECT 1.76 1.5 2.03 1.74 ;
 RECT 1.76 1.74 1.86 2.585 ;
 RECT 11.14 0.14 11.24 1.135 ;
 RECT 11.14 1.235 11.24 2.79 ;
 RECT 10.56 1.07 10.77 1.135 ;
 RECT 10.56 1.235 10.77 1.305 ;
 RECT 10.56 1.135 11.24 1.235 ;
 RECT 10.67 0.14 10.77 1.07 ;
 RECT 10.67 1.305 10.77 2.79 ;
 LAYER CO ;
 RECT 4.645 1.63 4.775 1.76 ;
 RECT 3.835 1.525 3.965 1.655 ;
 RECT 4.545 2.64 4.675 2.77 ;
 RECT 10.6 1.12 10.73 1.25 ;
 RECT 11.36 0.65 11.49 0.78 ;
 RECT 11.365 1.79 11.495 1.92 ;
 RECT 11.365 2.05 11.495 2.18 ;
 RECT 11.365 2.31 11.495 2.44 ;
 RECT 7.895 2.525 8.025 2.655 ;
 RECT 10.89 1.79 11.02 1.92 ;
 RECT 10.89 1.53 11.02 1.66 ;
 RECT 10.89 2.31 11.02 2.44 ;
 RECT 5.66 1.69 5.79 1.82 ;
 RECT 5.42 0.915 5.55 1.045 ;
 RECT 5.205 0.505 5.335 0.635 ;
 RECT 6.495 1.9 6.625 2.03 ;
 RECT 6.495 0.87 6.625 1 ;
 RECT 7.445 1.965 7.575 2.095 ;
 RECT 7.78 0.87 7.91 1 ;
 RECT 6.25 0.505 6.38 0.635 ;
 RECT 6.805 1.28 6.935 1.41 ;
 RECT 10.42 1.53 10.55 1.66 ;
 RECT 10.42 1.79 10.55 1.92 ;
 RECT 10.42 2.05 10.55 2.18 ;
 RECT 10.42 2.31 10.55 2.44 ;
 RECT 7.15 0.575 7.28 0.705 ;
 RECT 3.665 2.07 3.795 2.2 ;
 RECT 3.685 0.88 3.815 1.01 ;
 RECT 3.17 2.105 3.3 2.235 ;
 RECT 2.93 0.555 3.06 0.685 ;
 RECT 5.095 0.88 5.225 1.01 ;
 RECT 4.47 0.2 4.6 0.33 ;
 RECT 2.755 2.335 2.885 2.465 ;
 RECT 3.57 0.525 3.7 0.655 ;
 RECT 1.035 0.895 1.165 1.025 ;
 RECT 0.545 2.105 0.675 2.235 ;
 RECT 2.11 0.895 2.24 1.025 ;
 RECT 9.32 0.475 9.45 0.605 ;
 RECT 9.885 1.79 10.015 1.92 ;
 RECT 9.885 1.53 10.015 1.66 ;
 RECT 9.885 2.05 10.015 2.18 ;
 RECT 9.885 2.31 10.015 2.44 ;
 RECT 9.885 0.725 10.015 0.855 ;
 RECT 9.105 1.23 9.235 1.36 ;
 RECT 0.545 1.845 0.675 1.975 ;
 RECT 1.505 2.235 1.635 2.365 ;
 RECT 2.355 1.495 2.485 1.625 ;
 RECT 2.225 2.47 2.355 2.6 ;
 RECT 3.215 0.88 3.345 1.01 ;
 RECT 2.82 0.905 2.95 1.035 ;
 RECT 6 1.815 6.13 1.945 ;
 RECT 5.49 2.44 5.62 2.57 ;
 RECT 6.965 1.965 7.095 2.095 ;
 RECT 6.025 0.87 6.155 1 ;
 RECT 8.25 0.87 8.38 1 ;
 RECT 8.265 2.115 8.395 2.245 ;
 RECT 7.795 2.11 7.925 2.24 ;
 RECT 8.825 2.13 8.955 2.26 ;
 RECT 8.44 1.76 8.57 1.89 ;
 RECT 9.385 1.53 9.515 1.66 ;
 RECT 9.385 1.79 9.515 1.92 ;
 RECT 9.385 2.05 9.515 2.18 ;
 RECT 9.385 2.31 9.515 2.44 ;
 RECT 4.93 2.015 5.06 2.145 ;
 RECT 2.125 0.25 2.255 0.38 ;
 RECT 2.885 1.725 3.015 1.855 ;
 RECT 0.545 0.61 0.675 0.74 ;
 RECT 0.545 0.35 0.675 0.48 ;
 RECT 1.505 0.87 1.635 1 ;
 RECT 1.86 1.555 1.99 1.685 ;
 RECT 11.365 1.53 11.495 1.66 ;
 RECT 10.89 2.05 11.02 2.18 ;
 RECT 1.035 2.21 1.165 2.34 ;
 RECT 0.545 2.365 0.675 2.495 ;
 RECT 1.98 2.115 2.11 2.245 ;
 RECT 10.89 0.65 11.02 0.78 ;
 RECT 10.355 0.11 10.485 0.24 ;
 RECT 0.69 1.215 0.82 1.345 ;
 LAYER M1 ;
 RECT 3.5 0.52 5.41 0.66 ;
 RECT 5.125 0.47 5.41 0.52 ;
 RECT 2.105 0.845 2.245 1.18 ;
 RECT 2.105 1.18 2.49 1.335 ;
 RECT 2.35 1.335 2.49 2.11 ;
 RECT 1.91 2.11 2.49 2.25 ;
 RECT 4.925 1.04 5.6 1.05 ;
 RECT 4.36 0.91 5.6 1.04 ;
 RECT 4.36 0.9 5.23 0.91 ;
 RECT 4.925 1.08 5.065 2.2 ;
 RECT 4.925 1.05 5.23 1.08 ;
 RECT 3.785 1.52 4.5 1.66 ;
 RECT 5.09 0.81 5.23 0.9 ;
 RECT 4.36 1.04 4.5 1.52 ;
 RECT 5.205 1.36 5.345 2.1 ;
 RECT 5.205 2.24 5.345 2.355 ;
 RECT 4.13 2.355 5.345 2.495 ;
 RECT 2.75 2.515 4.27 2.655 ;
 RECT 2.815 0.735 2.955 1.72 ;
 RECT 2.815 1.72 3.065 1.775 ;
 RECT 2.75 1.775 3.065 1.86 ;
 RECT 2.75 1.86 2.955 2.005 ;
 RECT 2.75 2.005 2.89 2.515 ;
 RECT 2.925 0.505 3.065 0.535 ;
 RECT 4.13 2.495 4.27 2.515 ;
 RECT 2.815 0.535 3.065 0.735 ;
 RECT 6.61 2.32 6.75 2.52 ;
 RECT 5.74 0.5 6.455 0.64 ;
 RECT 5.74 0.64 5.88 1.22 ;
 RECT 5.205 2.1 6.105 2.18 ;
 RECT 5.205 2.18 6.75 2.24 ;
 RECT 5.965 2.24 6.75 2.32 ;
 RECT 5.205 1.22 5.88 1.36 ;
 RECT 6.61 2.52 8.105 2.66 ;
 RECT 3.505 1.805 4.78 1.945 ;
 RECT 3.505 1.945 3.87 1.96 ;
 RECT 3.505 1.22 3.82 1.36 ;
 RECT 3.68 0.805 3.82 1.22 ;
 RECT 3.59 1.96 3.87 2.215 ;
 RECT 3.505 1.36 3.645 1.805 ;
 RECT 4.64 1.56 4.78 1.805 ;
 RECT 6.96 2.1 7.145 2.24 ;
 RECT 7.79 2.03 7.93 2.24 ;
 RECT 6.915 1.96 7.145 2.1 ;
 RECT 6.96 2.24 7.93 2.38 ;
 RECT 6.49 1.815 6.7 1.895 ;
 RECT 6.49 0.805 6.63 1.675 ;
 RECT 7.395 1.815 7.625 2.1 ;
 RECT 6.42 1.895 6.7 2.035 ;
 RECT 6.49 1.675 8.68 1.815 ;
 RECT 9.1 1.18 9.24 2.505 ;
 RECT 8.38 1.815 8.68 1.915 ;
 RECT 8.54 1.915 8.68 2.505 ;
 RECT 8.54 2.505 9.24 2.645 ;
 RECT 5.65 1.685 6.16 1.81 ;
 RECT 5.65 1.81 6.2 1.825 ;
 RECT 6.02 0.78 6.16 1.685 ;
 RECT 5.65 1.615 5.79 1.685 ;
 RECT 5.65 1.825 5.79 1.895 ;
 RECT 5.93 1.825 6.2 1.95 ;
 RECT 6.8 1.21 6.94 1.395 ;
 RECT 8.82 1.005 8.96 1.395 ;
 RECT 8.82 1.535 8.96 2.32 ;
 RECT 6.8 1.395 8.96 1.535 ;
 RECT 9.595 0.535 9.735 0.865 ;
 RECT 8.2 0.865 9.735 1.005 ;
 RECT 9.595 0.395 10.735 0.535 ;
 RECT 10.595 0.535 10.735 1.315 ;
 RECT 1.03 0.825 1.17 1.195 ;
 RECT 1.03 1.335 1.17 2.41 ;
 RECT 1.825 0.665 1.965 1.195 ;
 RECT 1.03 1.195 1.965 1.335 ;
 RECT 3.21 0.36 3.35 0.875 ;
 RECT 3.225 1.015 3.365 2.035 ;
 RECT 2.53 0.36 2.67 0.525 ;
 RECT 3.165 2.035 3.365 2.305 ;
 RECT 3.165 0.875 3.42 1.015 ;
 RECT 1.825 0.525 2.67 0.665 ;
 RECT 2.53 0.22 3.35 0.36 ;
 END
END DFFASX2

MACRO DFFNARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.2 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.2 2.96 ;
 RECT 5.365 2.635 5.625 2.8 ;
 RECT 1.935 2.635 2.185 2.8 ;
 RECT 9.195 2.06 9.335 2.8 ;
 RECT 10.72 1.73 10.86 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.28 1.98 1.42 2.8 ;
 RECT 8.015 1.955 8.155 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.2 0.08 ;
 RECT 4.625 0.08 4.86 0.26 ;
 RECT 1.91 0.08 2.21 0.26 ;
 RECT 8.045 0.08 8.29 0.545 ;
 RECT 1.28 0.08 1.42 1.055 ;
 RECT 9.215 0.08 9.355 0.725 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 10.805 0.08 10.945 0.88 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.295 1.475 1.59 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.67 0.36 7.81 0.93 ;
 RECT 4.02 0.51 5.14 0.65 ;
 RECT 7.67 0.93 8.655 1.07 ;
 RECT 8.435 0.28 8.715 0.42 ;
 RECT 5.96 0.36 6.2 0.66 ;
 RECT 5 0.36 5.14 0.51 ;
 RECT 5 0.22 7.81 0.36 ;
 RECT 8.435 0.42 8.655 0.93 ;
 END
 ANTENNAGATEAREA 0.107 ;
 END RSTB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.78 1.105 10.105 1.425 ;
 RECT 9.78 0.55 9.92 1.105 ;
 RECT 9.78 1.425 9.92 2.35 ;
 END
 ANTENNADIFFAREA 0.575 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.245 2.015 10.56 2.38 ;
 RECT 10.245 0.7 10.385 2.015 ;
 END
 ANTENNADIFFAREA 0.456 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.32 1.16 0.85 1.525 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 3.695 1.71 3.795 2.475 ;
 RECT 3.735 0.65 3.835 1.33 ;
 RECT 3.695 1.475 3.925 1.71 ;
 RECT 9.525 0.21 9.625 1.225 ;
 RECT 9.525 1.455 9.625 2.775 ;
 RECT 9.28 1.225 9.625 1.455 ;
 RECT 10.505 0.33 10.605 1.09 ;
 RECT 10.505 1.325 10.605 2.79 ;
 RECT 10.49 1.09 10.7 1.325 ;
 RECT 2.72 2.33 2.82 2.685 ;
 RECT 4.995 1.79 5.095 2.685 ;
 RECT 2.6 2.09 2.82 2.33 ;
 RECT 2.72 2.685 5.095 2.785 ;
 RECT 5.45 0.575 6.64 0.675 ;
 RECT 6.54 0.675 6.64 1.35 ;
 RECT 7.875 0.265 7.975 1.32 ;
 RECT 5.45 0.46 5.68 0.575 ;
 RECT 5.45 0.675 5.68 0.69 ;
 RECT 6.54 0.265 6.64 0.575 ;
 RECT 6.985 1.545 7.085 2.405 ;
 RECT 6.54 0.165 7.975 0.265 ;
 RECT 6.54 1.35 6.83 1.445 ;
 RECT 6.54 1.445 7.085 1.45 ;
 RECT 6.73 1.45 7.085 1.545 ;
 RECT 3.245 0.705 3.345 1.21 ;
 RECT 2.675 1.16 2.92 1.21 ;
 RECT 2.675 1.21 3.345 1.31 ;
 RECT 2.675 1.31 2.92 1.405 ;
 RECT 3.245 0.47 3.53 0.705 ;
 RECT 1.065 0.175 1.165 1.335 ;
 RECT 1.065 1.435 1.165 2.465 ;
 RECT 0.665 1.335 1.165 1.435 ;
 RECT 0.665 1.275 0.885 1.335 ;
 RECT 0.665 1.435 0.885 1.505 ;
 RECT 7.8 1.64 7.9 2.585 ;
 RECT 6.58 2.47 6.8 2.585 ;
 RECT 6.58 2.585 7.9 2.685 ;
 RECT 6.58 2.685 6.8 2.71 ;
 RECT 3.2 1.685 3.3 2.495 ;
 RECT 1.88 1.52 2.48 1.585 ;
 RECT 1.88 1.585 3.3 1.62 ;
 RECT 1.88 1.62 2.125 1.69 ;
 RECT 2.315 1.62 3.3 1.685 ;
 RECT 2.315 1.685 2.415 2.27 ;
 RECT 1.88 1.44 2.125 1.52 ;
 RECT 2.38 0.685 2.48 1.52 ;
 RECT 2.7 0.285 2.8 0.585 ;
 RECT 2.7 0.185 4.535 0.285 ;
 RECT 4.435 0.285 4.535 1.24 ;
 RECT 2.38 0.585 2.8 0.685 ;
 RECT 1.54 0.655 1.64 1.48 ;
 RECT 1.345 1.48 1.64 1.72 ;
 RECT 1.54 1.72 1.64 2.37 ;
 RECT 7.48 0.645 7.58 1.24 ;
 RECT 7.48 1.45 7.58 2.37 ;
 RECT 7.46 1.24 7.695 1.45 ;
 RECT 7.01 0.685 7.11 1.255 ;
 RECT 6.935 0.455 7.165 0.685 ;
 RECT 5.96 0.875 6.355 1.105 ;
 RECT 6.255 1.105 6.355 1.64 ;
 RECT 6.255 1.64 6.49 1.87 ;
 RECT 8.89 1.32 8.99 2.545 ;
 RECT 8.59 0.47 8.69 1.22 ;
 RECT 8.59 1.22 8.99 1.32 ;
 RECT 8.46 0.23 8.69 0.47 ;
 RECT 4.135 0.695 4.235 1.61 ;
 RECT 4.17 1.71 4.27 2.48 ;
 RECT 4.135 1.61 4.27 1.71 ;
 RECT 4.015 0.465 4.255 0.695 ;
 RECT 8.29 0.65 8.39 1.71 ;
 RECT 8.29 1.71 8.535 1.95 ;
 RECT 8.29 1.95 8.39 2.56 ;
 RECT 5.095 0.635 5.195 1.475 ;
 RECT 5.465 1.705 5.565 2.52 ;
 RECT 5.3 1.61 5.565 1.705 ;
 RECT 5.095 1.475 5.565 1.61 ;
 RECT 3.695 1.33 3.835 1.475 ;
 LAYER CO ;
 RECT 9.22 0.505 9.35 0.635 ;
 RECT 6.31 1.69 6.44 1.82 ;
 RECT 4.395 1.825 4.525 1.955 ;
 RECT 3.915 2.105 4.045 2.235 ;
 RECT 1.94 1.495 2.07 1.625 ;
 RECT 2.005 2.64 2.135 2.77 ;
 RECT 3.445 2.07 3.575 2.2 ;
 RECT 3.465 0.88 3.595 1.01 ;
 RECT 2.95 2.105 3.08 2.235 ;
 RECT 2.995 0.88 3.125 1.01 ;
 RECT 2.73 1.205 2.86 1.335 ;
 RECT 1.81 1.995 1.94 2.125 ;
 RECT 1.89 0.875 2.02 1.005 ;
 RECT 1.285 2.05 1.415 2.18 ;
 RECT 1.285 0.875 1.415 1.005 ;
 RECT 0.815 0.875 0.945 1.005 ;
 RECT 2.03 0.125 2.16 0.255 ;
 RECT 7.23 0.87 7.36 1 ;
 RECT 8.11 0.4 8.24 0.53 ;
 RECT 8.36 1.765 8.49 1.895 ;
 RECT 2.65 2.145 2.78 2.275 ;
 RECT 2.535 1.825 2.665 1.955 ;
 RECT 3.35 0.525 3.48 0.655 ;
 RECT 7.23 0.87 7.36 1 ;
 RECT 6.76 0.87 6.89 1 ;
 RECT 6.985 0.505 7.115 0.635 ;
 RECT 7.51 1.28 7.64 1.41 ;
 RECT 8.81 0.87 8.94 1 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 10.81 0.68 10.94 0.81 ;
 RECT 10.25 1.65 10.38 1.78 ;
 RECT 10.25 1.91 10.38 2.04 ;
 RECT 10.25 2.17 10.38 2.3 ;
 RECT 10.725 2.32 10.855 2.45 ;
 RECT 10.25 0.75 10.38 0.88 ;
 RECT 9.33 1.275 9.46 1.405 ;
 RECT 10.725 1.8 10.855 1.93 ;
 RECT 10.725 2.06 10.855 2.19 ;
 RECT 9.785 0.615 9.915 0.745 ;
 RECT 9.785 1.87 9.915 2 ;
 RECT 9.785 2.13 9.915 2.26 ;
 RECT 0.815 2.06 0.945 2.19 ;
 RECT 5.49 0.51 5.62 0.64 ;
 RECT 6.03 0.915 6.16 1.045 ;
 RECT 8.51 0.285 8.64 0.415 ;
 RECT 4.07 0.515 4.2 0.645 ;
 RECT 4.675 0.12 4.805 0.25 ;
 RECT 7.23 1.99 7.36 2.12 ;
 RECT 2.6 0.905 2.73 1.035 ;
 RECT 1.395 1.535 1.525 1.665 ;
 RECT 8.02 2.03 8.15 2.16 ;
 RECT 9.2 2.13 9.33 2.26 ;
 RECT 8.64 2.13 8.77 2.26 ;
 RECT 5.355 1.515 5.485 1.645 ;
 RECT 3.745 1.525 3.875 1.655 ;
 RECT 5.69 0.88 5.82 1.01 ;
 RECT 5.685 2.015 5.815 2.145 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 5.415 2.64 5.545 2.77 ;
 RECT 4.745 2.125 4.875 2.255 ;
 RECT 6.63 2.525 6.76 2.655 ;
 RECT 6.735 1.815 6.865 1.945 ;
 RECT 10.53 1.14 10.66 1.27 ;
 RECT 0.715 1.325 0.845 1.455 ;
 LAYER M1 ;
 RECT 3.845 2.1 4.945 2.26 ;
 RECT 3.28 0.52 3.88 0.66 ;
 RECT 3.74 0.66 3.88 0.79 ;
 RECT 5.28 0.505 5.68 0.645 ;
 RECT 3.74 0.79 5.42 0.93 ;
 RECT 5.28 0.645 5.42 0.79 ;
 RECT 7.505 1.395 8.945 1.535 ;
 RECT 8.805 0.76 8.945 0.965 ;
 RECT 8.805 1.105 8.945 1.395 ;
 RECT 8.635 1.535 8.775 2.33 ;
 RECT 7.505 1.21 7.645 1.395 ;
 RECT 9.495 0.36 9.635 0.965 ;
 RECT 8.805 0.965 9.635 1.105 ;
 RECT 10.525 0.36 10.665 1.34 ;
 RECT 9.495 0.22 10.665 0.36 ;
 RECT 2.595 1.385 2.735 1.82 ;
 RECT 2.465 1.825 2.785 1.96 ;
 RECT 2.465 1.82 2.735 1.825 ;
 RECT 2.645 1.96 2.785 2.345 ;
 RECT 2.595 0.84 2.735 1.155 ;
 RECT 2.595 1.155 2.865 1.385 ;
 RECT 2.325 2.515 5.225 2.655 ;
 RECT 5.085 2.495 5.225 2.515 ;
 RECT 1.805 1.475 2.145 2.35 ;
 RECT 2.325 2.49 2.465 2.515 ;
 RECT 1.885 0.825 2.025 1.475 ;
 RECT 1.805 2.35 2.465 2.49 ;
 RECT 6.4 0.58 7.19 0.64 ;
 RECT 6.4 0.64 6.86 0.72 ;
 RECT 6.68 0.5 7.19 0.58 ;
 RECT 5.96 1.21 6.54 1.35 ;
 RECT 6.56 2.24 6.7 2.52 ;
 RECT 5.96 1.35 6.1 2.1 ;
 RECT 5.96 2.24 6.1 2.355 ;
 RECT 5.96 2.1 6.7 2.24 ;
 RECT 5.085 2.355 6.1 2.495 ;
 RECT 6.4 0.72 6.54 1.21 ;
 RECT 6.56 2.52 6.83 2.66 ;
 RECT 3.285 1.82 5.49 1.96 ;
 RECT 3.285 1.22 3.6 1.36 ;
 RECT 3.46 0.805 3.6 1.22 ;
 RECT 3.37 1.96 3.65 2.215 ;
 RECT 5.35 1.44 5.49 1.82 ;
 RECT 3.285 1.36 3.425 1.82 ;
 RECT 5.62 0.875 6.23 1.05 ;
 RECT 5.62 1.05 5.82 1.08 ;
 RECT 5.07 1.08 5.82 1.22 ;
 RECT 5.62 1.22 5.82 1.255 ;
 RECT 5.68 1.255 5.82 2.215 ;
 RECT 3.675 1.52 5.21 1.66 ;
 RECT 5.07 1.22 5.21 1.52 ;
 RECT 6.24 1.685 6.965 1.825 ;
 RECT 6.685 0.865 6.965 1.685 ;
 RECT 6.665 1.825 6.965 1.95 ;
 RECT 8.915 1.92 9.055 2.505 ;
 RECT 7.225 1.675 8.495 1.815 ;
 RECT 8.355 2.505 9.055 2.645 ;
 RECT 8.355 1.815 8.495 2.505 ;
 RECT 7.225 1.815 7.435 1.985 ;
 RECT 7.225 0.805 7.365 1.675 ;
 RECT 7.155 1.985 7.435 2.125 ;
 RECT 9.15 1.41 9.29 1.78 ;
 RECT 9.15 1.27 9.53 1.41 ;
 RECT 8.915 1.78 9.29 1.92 ;
 RECT 1 1.01 1.14 1.195 ;
 RECT 1 1.335 1.14 2.055 ;
 RECT 0.745 0.87 1.14 1.01 ;
 RECT 0.745 2.055 1.14 2.195 ;
 RECT 1.56 0.67 1.7 1.195 ;
 RECT 1 1.195 1.7 1.335 ;
 RECT 1.56 0.53 2.51 0.67 ;
 RECT 2.37 0.22 3.13 0.36 ;
 RECT 2.99 0.36 3.13 0.875 ;
 RECT 2.945 2.035 3.145 2.305 ;
 RECT 3.005 1.015 3.145 2.035 ;
 RECT 2.37 0.36 2.51 0.53 ;
 RECT 2.925 0.875 3.2 1.015 ;
 END
END DFFNARX1

MACRO DFFNARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.84 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.84 2.96 ;
 RECT 5.355 2.635 5.615 2.8 ;
 RECT 1.84 2.625 2.09 2.8 ;
 RECT 1.27 1.98 1.41 2.8 ;
 RECT 8.005 1.955 8.145 2.8 ;
 RECT 9.185 2.06 9.325 2.8 ;
 RECT 11.285 1.73 11.425 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 10.32 2.01 10.46 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.84 0.08 ;
 RECT 1.27 0.08 1.41 0.98 ;
 RECT 4.615 0.08 4.85 0.495 ;
 RECT 11.595 0.08 11.735 0.94 ;
 RECT 9.205 0.08 9.345 0.67 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 8.1 0.08 8.24 0.6 ;
 RECT 2.015 0.08 2.155 0.39 ;
 RECT 10.475 0.08 10.615 0.3 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.265 1.415 1.58 1.84 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.66 0.36 7.8 0.785 ;
 RECT 4.055 0.635 5.13 0.775 ;
 RECT 7.66 0.785 8.635 0.925 ;
 RECT 8.495 0.225 8.635 0.785 ;
 RECT 5.96 0.36 6.2 0.6 ;
 RECT 4.99 0.36 5.13 0.635 ;
 RECT 4.99 0.22 7.8 0.36 ;
 RECT 4.055 0.445 4.195 0.635 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.85 0.72 9.99 2.07 ;
 RECT 9.64 2.07 9.99 2.57 ;
 END
 ANTENNADIFFAREA 0.578 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.6 2.015 10.95 2.38 ;
 RECT 10.81 0.845 11.11 0.985 ;
 RECT 10.81 2.38 10.95 2.61 ;
 RECT 10.97 0.72 11.11 0.845 ;
 RECT 10.81 0.985 10.95 2.015 ;
 END
 ANTENNADIFFAREA 0.6 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.31 1.135 0.655 1.52 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END D

 OBS
 LAYER PO ;
 RECT 5.455 1.745 5.555 2.52 ;
 RECT 5.085 0.635 5.185 1.44 ;
 RECT 5.085 1.44 5.555 1.54 ;
 RECT 3.685 1.33 3.825 1.475 ;
 RECT 3.685 1.71 3.785 2.475 ;
 RECT 3.725 0.65 3.825 1.33 ;
 RECT 3.685 1.475 3.915 1.71 ;
 RECT 5.43 0.59 6.63 0.69 ;
 RECT 6.53 0.69 6.63 1.35 ;
 RECT 7.865 0.265 7.965 1.22 ;
 RECT 5.43 0.46 5.66 0.59 ;
 RECT 6.53 0.265 6.63 0.59 ;
 RECT 6.975 1.545 7.075 2.455 ;
 RECT 6.53 0.165 7.965 0.265 ;
 RECT 6.53 1.35 6.82 1.445 ;
 RECT 6.53 1.445 7.075 1.45 ;
 RECT 6.72 1.45 7.075 1.545 ;
 RECT 1.055 0.65 1.155 1.2 ;
 RECT 1.055 1.45 1.155 2.61 ;
 RECT 0.345 1.2 1.155 1.45 ;
 RECT 11.38 0.46 11.48 1.165 ;
 RECT 11.07 1.265 11.48 1.425 ;
 RECT 11.07 1.425 11.17 2.79 ;
 RECT 10.575 1.165 11.48 1.265 ;
 RECT 10.755 0.46 10.855 1.165 ;
 RECT 10.575 1.265 10.675 2.79 ;
 RECT 9.27 1.05 9.735 1.09 ;
 RECT 9.27 1.09 10.205 1.19 ;
 RECT 9.635 0.135 9.735 1.05 ;
 RECT 9.635 1.28 9.735 2.79 ;
 RECT 9.27 1.19 9.735 1.28 ;
 RECT 10.105 0.135 10.205 1.09 ;
 RECT 10.105 1.19 10.205 2.79 ;
 RECT 7.79 1.575 7.89 2.635 ;
 RECT 6.57 2.635 7.89 2.735 ;
 RECT 6.57 2.4 6.79 2.635 ;
 RECT 1.87 1.52 2.47 1.585 ;
 RECT 1.87 1.585 3.29 1.62 ;
 RECT 1.87 1.62 2.115 1.69 ;
 RECT 3.19 1.685 3.29 2.48 ;
 RECT 2.305 1.685 2.405 2.3 ;
 RECT 1.87 1.44 2.115 1.52 ;
 RECT 2.37 0.285 2.47 1.52 ;
 RECT 2.305 1.62 3.29 1.685 ;
 RECT 2.37 0.185 4.525 0.285 ;
 RECT 4.425 0.285 4.525 1.24 ;
 RECT 1.53 0.655 1.63 1.495 ;
 RECT 1.335 1.495 1.63 1.745 ;
 RECT 1.53 1.745 1.63 2.37 ;
 RECT 4.985 1.79 5.085 2.68 ;
 RECT 2.61 2.075 2.82 2.68 ;
 RECT 2.61 2.68 5.085 2.78 ;
 RECT 3.235 0.705 3.335 1.16 ;
 RECT 3.235 0.47 3.52 0.705 ;
 RECT 2.65 1.16 3.335 1.265 ;
 RECT 2.65 1.265 2.895 1.405 ;
 RECT 5.95 0.875 6.345 1.105 ;
 RECT 6.245 1.105 6.345 1.64 ;
 RECT 6.245 1.64 6.48 1.87 ;
 RECT 8.88 1.32 8.98 2.77 ;
 RECT 8.58 0.47 8.68 1.22 ;
 RECT 8.58 1.22 8.98 1.32 ;
 RECT 8.45 0.23 8.68 0.47 ;
 RECT 4.125 0.695 4.225 1.61 ;
 RECT 4.16 1.71 4.26 2.48 ;
 RECT 4.125 1.61 4.26 1.71 ;
 RECT 4.005 0.465 4.245 0.695 ;
 RECT 7.47 0.645 7.57 1.18 ;
 RECT 7.47 1.39 7.57 2.165 ;
 RECT 7.45 1.18 7.685 1.39 ;
 RECT 7 0.685 7.1 1.255 ;
 RECT 6.925 0.455 7.155 0.685 ;
 RECT 8.28 0.65 8.38 1.71 ;
 RECT 8.28 1.71 8.525 1.95 ;
 RECT 8.28 1.95 8.38 2.765 ;
 RECT 5.29 1.54 5.555 1.745 ;
 LAYER CO ;
 RECT 6.3 1.69 6.43 1.82 ;
 RECT 4.385 1.825 4.515 1.955 ;
 RECT 3.905 2.125 4.035 2.255 ;
 RECT 1.93 1.495 2.06 1.625 ;
 RECT 1.91 2.63 2.04 2.76 ;
 RECT 3.435 2.07 3.565 2.2 ;
 RECT 3.455 0.88 3.585 1.01 ;
 RECT 2.94 2.105 3.07 2.235 ;
 RECT 2.985 0.88 3.115 1.01 ;
 RECT 2.705 1.205 2.835 1.335 ;
 RECT 2.59 0.905 2.72 1.035 ;
 RECT 1.275 2.05 1.405 2.18 ;
 RECT 1.275 0.8 1.405 0.93 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 0.805 2.115 0.935 2.245 ;
 RECT 10.48 0.12 10.61 0.25 ;
 RECT 10.325 2.085 10.455 2.215 ;
 RECT 10.325 2.35 10.455 2.48 ;
 RECT 0.405 1.255 0.535 1.385 ;
 RECT 1.395 1.55 1.525 1.68 ;
 RECT 10.815 1.565 10.945 1.695 ;
 RECT 10.815 1.83 10.945 1.96 ;
 RECT 10.815 2.09 10.945 2.22 ;
 RECT 10.815 2.39 10.945 2.52 ;
 RECT 9.855 2.085 9.985 2.215 ;
 RECT 2.65 2.13 2.78 2.26 ;
 RECT 5.47 0.51 5.6 0.64 ;
 RECT 8.35 1.765 8.48 1.895 ;
 RECT 8.01 2.01 8.14 2.14 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 6.62 2.465 6.75 2.595 ;
 RECT 6.725 1.815 6.855 1.945 ;
 RECT 11.13 1.24 11.26 1.37 ;
 RECT 11.6 0.755 11.73 0.885 ;
 RECT 9.855 2.35 9.985 2.48 ;
 RECT 11.29 2.32 11.42 2.45 ;
 RECT 10.975 0.77 11.105 0.9 ;
 RECT 9.32 1.1 9.45 1.23 ;
 RECT 11.29 1.8 11.42 1.93 ;
 RECT 11.29 2.06 11.42 2.19 ;
 RECT 9.855 0.77 9.985 0.9 ;
 RECT 9.21 0.485 9.34 0.615 ;
 RECT 6.02 0.915 6.15 1.045 ;
 RECT 8.5 0.285 8.63 0.415 ;
 RECT 8.105 0.4 8.235 0.53 ;
 RECT 4.06 0.515 4.19 0.645 ;
 RECT 4.665 0.36 4.795 0.49 ;
 RECT 7.22 1.815 7.35 1.945 ;
 RECT 7.22 0.87 7.35 1 ;
 RECT 6.75 0.87 6.88 1 ;
 RECT 6.975 0.505 7.105 0.635 ;
 RECT 7.5 1.22 7.63 1.35 ;
 RECT 8.8 0.87 8.93 1 ;
 RECT 1.75 1.995 1.88 2.125 ;
 RECT 1.88 0.875 2.01 1.005 ;
 RECT 9.19 2.19 9.32 2.32 ;
 RECT 8.63 2.17 8.76 2.3 ;
 RECT 5.345 1.555 5.475 1.685 ;
 RECT 3.735 1.525 3.865 1.655 ;
 RECT 5.68 0.88 5.81 1.01 ;
 RECT 5.675 2.015 5.805 2.145 ;
 RECT 2.02 0.21 2.15 0.34 ;
 RECT 5.405 2.64 5.535 2.77 ;
 RECT 4.735 2.125 4.865 2.255 ;
 RECT 2.525 1.825 2.655 1.955 ;
 RECT 3.34 0.525 3.47 0.655 ;
 LAYER M1 ;
 RECT 3.835 2.12 4.935 2.26 ;
 RECT 5.67 1.05 5.81 1.195 ;
 RECT 4.395 1.195 5.81 1.335 ;
 RECT 5.67 1.335 5.81 2.215 ;
 RECT 5.61 0.91 6.22 1.015 ;
 RECT 5.61 0.875 5.88 0.91 ;
 RECT 5.67 1.015 6.22 1.05 ;
 RECT 3.665 1.52 4.535 1.66 ;
 RECT 4.395 1.335 4.535 1.52 ;
 RECT 3.27 0.52 3.915 0.66 ;
 RECT 3.775 0.66 3.915 0.915 ;
 RECT 3.775 0.915 5.41 1.055 ;
 RECT 5.27 0.505 5.66 0.645 ;
 RECT 5.27 0.645 5.41 0.915 ;
 RECT 2.585 1.155 2.84 1.385 ;
 RECT 2.585 1.385 2.785 1.82 ;
 RECT 2.585 1.96 2.785 2.335 ;
 RECT 2.585 0.845 2.725 1.155 ;
 RECT 2.455 1.82 2.785 1.96 ;
 RECT 7.495 1.17 7.635 1.395 ;
 RECT 7.495 1.395 8.935 1.535 ;
 RECT 8.795 0.955 8.935 1.395 ;
 RECT 8.625 1.535 8.765 2.36 ;
 RECT 9.485 0.58 9.625 0.815 ;
 RECT 8.795 0.815 9.625 0.955 ;
 RECT 11.25 0.58 11.39 1.17 ;
 RECT 11.125 1.17 11.39 1.235 ;
 RECT 9.485 0.44 11.39 0.58 ;
 RECT 11.125 1.375 11.39 1.44 ;
 RECT 11.09 1.235 11.39 1.375 ;
 RECT 7.215 1.815 7.425 1.87 ;
 RECT 7.215 0.805 7.355 1.675 ;
 RECT 7.145 1.87 7.425 2.01 ;
 RECT 8.905 1.92 9.045 2.505 ;
 RECT 7.215 1.675 8.485 1.815 ;
 RECT 8.345 2.505 9.045 2.645 ;
 RECT 8.345 1.815 8.485 2.505 ;
 RECT 9.14 1.235 9.28 1.78 ;
 RECT 9.14 1.095 9.52 1.235 ;
 RECT 8.905 1.78 9.28 1.92 ;
 RECT 6.23 1.685 6.885 1.81 ;
 RECT 6.745 1.005 6.885 1.685 ;
 RECT 6.23 1.81 6.925 1.825 ;
 RECT 6.655 1.825 6.925 1.95 ;
 RECT 6.675 0.865 6.955 1.005 ;
 RECT 0.8 0.81 0.94 1.125 ;
 RECT 0.8 1.265 0.94 2.315 ;
 RECT 2.98 0.665 3.12 2.035 ;
 RECT 1.55 0.67 1.69 1.125 ;
 RECT 1.55 0.53 3.12 0.665 ;
 RECT 0.8 1.125 1.69 1.265 ;
 RECT 1.55 0.665 2.435 0.67 ;
 RECT 2.295 0.525 3.12 0.53 ;
 RECT 2.935 2.035 3.12 2.17 ;
 RECT 2.935 2.17 3.075 2.305 ;
 RECT 2.23 2.51 5.215 2.65 ;
 RECT 5.075 2.495 5.215 2.51 ;
 RECT 1.79 1.475 2.135 1.63 ;
 RECT 1.79 1.63 1.93 1.99 ;
 RECT 1.875 0.825 2.015 1.475 ;
 RECT 1.79 2.13 1.93 2.345 ;
 RECT 1.68 1.99 1.93 2.13 ;
 RECT 1.79 2.345 2.37 2.485 ;
 RECT 2.23 2.485 2.37 2.51 ;
 RECT 5.075 2.355 6.09 2.495 ;
 RECT 5.95 1.35 6.09 2.1 ;
 RECT 5.95 2.1 6.69 2.24 ;
 RECT 5.95 2.24 6.09 2.355 ;
 RECT 6.55 2.24 6.69 2.46 ;
 RECT 5.95 1.21 6.53 1.35 ;
 RECT 6.55 2.46 6.82 2.6 ;
 RECT 6.67 0.5 7.18 0.58 ;
 RECT 6.39 0.58 7.18 0.64 ;
 RECT 6.39 0.64 6.85 0.72 ;
 RECT 6.39 0.72 6.53 1.21 ;
 RECT 3.275 1.82 5.48 1.96 ;
 RECT 3.275 1.22 3.59 1.36 ;
 RECT 3.45 0.805 3.59 1.22 ;
 RECT 3.36 1.96 3.64 2.215 ;
 RECT 5.34 1.485 5.48 1.82 ;
 RECT 3.275 1.36 3.415 1.82 ;
 END
END DFFNARX2

MACRO DFFNASRNX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.2 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.2 2.96 ;
 RECT 1.935 2.635 2.185 2.8 ;
 RECT 5.365 2.635 5.625 2.8 ;
 RECT 1.28 1.98 1.42 2.8 ;
 RECT 9.175 2.085 9.315 2.8 ;
 RECT 10.295 2.06 10.435 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 6.385 2.38 6.525 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.2 0.08 ;
 RECT 1.91 0.08 2.21 0.26 ;
 RECT 4.625 0.08 4.86 0.26 ;
 RECT 8.645 0.08 8.9 0.285 ;
 RECT 1.28 0.08 1.42 1.055 ;
 RECT 10.315 0.08 10.455 0.725 ;
 RECT 0.3 0.08 0.44 0.775 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.58 1.475 1.91 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.295 0.36 8.435 0.505 ;
 RECT 4.02 0.51 5.175 0.65 ;
 RECT 8.295 0.505 9.28 0.645 ;
 RECT 9.06 0.28 9.34 0.42 ;
 RECT 6.02 0.36 6.43 0.6 ;
 RECT 5.035 0.22 8.435 0.36 ;
 RECT 5.035 0.36 5.175 0.51 ;
 RECT 9.14 0.225 9.28 0.28 ;
 RECT 9.06 0.42 9.28 0.505 ;
 END
 ANTENNAGATEAREA 0.117 ;
 END RSTB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.92 1.475 1.275 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.88 0.5 8.155 0.76 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.88 1.075 11.02 2.35 ;
 RECT 10.595 0.755 11.02 1.075 ;
 RECT 10.88 0.55 11.02 0.755 ;
 END
 ANTENNADIFFAREA 0.544 ;
 END QN

 OBS
 LAYER PO ;
 RECT 6.44 1.64 6.675 1.87 ;
 RECT 9.295 1.63 9.53 1.745 ;
 RECT 9.43 1.745 9.53 2.56 ;
 RECT 8.915 0.65 9.015 1.53 ;
 RECT 8.915 1.53 9.53 1.63 ;
 RECT 3.245 0.705 3.345 1.21 ;
 RECT 3.245 0.47 3.53 0.705 ;
 RECT 2.675 1.16 2.92 1.21 ;
 RECT 2.675 1.31 2.92 1.405 ;
 RECT 2.675 1.21 3.345 1.31 ;
 RECT 1.54 0.655 1.64 1.48 ;
 RECT 1.54 1.48 1.85 1.72 ;
 RECT 1.54 1.72 1.64 2.37 ;
 RECT 2.065 1.44 2.48 1.585 ;
 RECT 2.065 1.585 3.3 1.685 ;
 RECT 3.2 1.685 3.3 2.495 ;
 RECT 2.315 1.69 2.415 2.27 ;
 RECT 2.38 0.685 2.48 1.44 ;
 RECT 2.065 1.685 2.415 1.69 ;
 RECT 4.435 0.285 4.535 1.24 ;
 RECT 2.7 0.185 4.535 0.285 ;
 RECT 2.7 0.285 2.8 0.585 ;
 RECT 2.38 0.585 2.8 0.685 ;
 RECT 4.995 1.79 5.095 2.685 ;
 RECT 2.72 2.33 2.82 2.685 ;
 RECT 2.72 2.685 5.095 2.785 ;
 RECT 2.6 2.09 2.82 2.33 ;
 RECT 3.695 1.33 3.835 1.475 ;
 RECT 3.695 1.71 3.795 2.475 ;
 RECT 3.735 0.65 3.835 1.33 ;
 RECT 3.695 1.475 3.925 1.71 ;
 RECT 5.3 1.61 5.565 1.82 ;
 RECT 5.465 1.82 5.565 2.49 ;
 RECT 4.895 0.625 4.995 1.51 ;
 RECT 4.895 1.51 5.565 1.61 ;
 RECT 8.745 2.47 9.06 2.71 ;
 RECT 8.96 1.83 9.06 2.47 ;
 RECT 10.63 0.13 10.73 1.17 ;
 RECT 10.63 1.4 10.73 2.775 ;
 RECT 10.27 1.17 10.73 1.4 ;
 RECT 9.99 1.32 10.09 2.545 ;
 RECT 9.215 0.47 9.315 1.22 ;
 RECT 9.215 1.22 10.09 1.32 ;
 RECT 9.085 0.23 9.315 0.47 ;
 RECT 4.135 0.695 4.235 1.61 ;
 RECT 4.17 1.71 4.27 2.48 ;
 RECT 4.135 1.61 4.27 1.71 ;
 RECT 4.015 0.465 4.255 0.695 ;
 RECT 7.66 0.645 7.76 1.24 ;
 RECT 7.66 1.24 7.905 1.45 ;
 RECT 7.66 1.45 7.76 2.37 ;
 RECT 7.19 0.685 7.29 1.255 ;
 RECT 7.115 0.455 7.345 0.685 ;
 RECT 1.065 0.635 1.165 1.495 ;
 RECT 1.065 1.725 1.165 2.465 ;
 RECT 0.985 1.495 1.205 1.725 ;
 RECT 5.77 1.33 5.87 1.565 ;
 RECT 6.16 1.665 6.26 2.69 ;
 RECT 8.135 0.73 8.235 2.69 ;
 RECT 7.94 0.635 8.235 0.73 ;
 RECT 7.94 0.5 8.17 0.635 ;
 RECT 5.25 0.635 5.35 1.23 ;
 RECT 5.25 1.23 5.87 1.33 ;
 RECT 5.77 1.565 6.26 1.665 ;
 RECT 6.16 2.69 8.235 2.79 ;
 RECT 6.72 0.265 6.82 0.585 ;
 RECT 6.72 0.685 6.82 1.35 ;
 RECT 7.165 1.545 7.265 2.295 ;
 RECT 8.475 0.265 8.575 1.32 ;
 RECT 5.615 0.455 5.845 0.585 ;
 RECT 5.615 0.585 6.82 0.685 ;
 RECT 6.72 0.165 8.575 0.265 ;
 RECT 6.91 1.45 7.265 1.545 ;
 RECT 6.72 1.35 7.01 1.445 ;
 RECT 6.72 1.445 7.265 1.45 ;
 RECT 6.145 0.865 6.54 1.095 ;
 RECT 6.44 1.095 6.54 1.64 ;
 LAYER CO ;
 RECT 9.35 1.57 9.48 1.7 ;
 RECT 5.355 1.63 5.485 1.76 ;
 RECT 2.535 1.825 2.665 1.955 ;
 RECT 4.745 2.125 4.875 2.255 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 10.885 0.615 11.015 0.745 ;
 RECT 10.885 1.87 11.015 2 ;
 RECT 10.885 2.13 11.015 2.26 ;
 RECT 10.32 0.505 10.45 0.635 ;
 RECT 3.445 2.07 3.575 2.2 ;
 RECT 3.465 0.88 3.595 1.01 ;
 RECT 6.215 0.915 6.345 1.045 ;
 RECT 2.135 1.495 2.265 1.625 ;
 RECT 8.72 0.15 8.85 0.28 ;
 RECT 5.665 0.505 5.795 0.635 ;
 RECT 7.41 1.9 7.54 2.03 ;
 RECT 7.41 0.87 7.54 1 ;
 RECT 8.36 1.92 8.49 2.05 ;
 RECT 0.815 2.055 0.945 2.185 ;
 RECT 2.6 0.905 2.73 1.035 ;
 RECT 7.88 1.965 8.01 2.095 ;
 RECT 6.94 0.87 7.07 1 ;
 RECT 7.165 0.505 7.295 0.635 ;
 RECT 9.435 0.87 9.565 1 ;
 RECT 9.18 2.17 9.31 2.3 ;
 RECT 8.71 2.135 8.84 2.265 ;
 RECT 10.3 2.13 10.43 2.26 ;
 RECT 3.35 0.525 3.48 0.655 ;
 RECT 1.025 1.545 1.155 1.675 ;
 RECT 3.745 1.525 3.875 1.655 ;
 RECT 5.69 0.88 5.82 1.01 ;
 RECT 5.685 2.015 5.815 2.145 ;
 RECT 2.03 0.125 2.16 0.255 ;
 RECT 5.415 2.64 5.545 2.77 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 7.99 0.55 8.12 0.68 ;
 RECT 8.81 2.525 8.94 2.655 ;
 RECT 6.915 1.815 7.045 1.945 ;
 RECT 6.39 2.44 6.52 2.57 ;
 RECT 10.32 1.225 10.45 1.355 ;
 RECT 6.495 1.69 6.625 1.82 ;
 RECT 4.395 1.82 4.525 1.95 ;
 RECT 3.915 2.105 4.045 2.235 ;
 RECT 2.005 2.64 2.135 2.77 ;
 RECT 4.07 0.515 4.2 0.645 ;
 RECT 4.675 0.12 4.805 0.25 ;
 RECT 2.95 2.105 3.08 2.235 ;
 RECT 2.995 0.88 3.125 1.01 ;
 RECT 2.73 1.205 2.86 1.335 ;
 RECT 9.135 0.285 9.265 0.415 ;
 RECT 1.68 1.535 1.81 1.665 ;
 RECT 1.81 1.995 1.94 2.125 ;
 RECT 1.89 0.875 2.02 1.005 ;
 RECT 1.285 2.05 1.415 2.18 ;
 RECT 1.285 0.875 1.415 1.005 ;
 RECT 0.815 0.875 0.945 1.005 ;
 RECT 9.74 2.13 9.87 2.26 ;
 RECT 2.65 2.145 2.78 2.275 ;
 RECT 7.72 1.28 7.85 1.41 ;
 LAYER M1 ;
 RECT 3.845 2.12 4.945 2.24 ;
 RECT 3.845 2.1 4.115 2.12 ;
 RECT 3.91 2.24 4.945 2.26 ;
 RECT 3.28 0.52 3.88 0.66 ;
 RECT 3.74 0.66 3.88 0.79 ;
 RECT 3.74 0.79 5.455 0.93 ;
 RECT 5.315 0.5 5.865 0.64 ;
 RECT 5.315 0.64 5.455 0.79 ;
 RECT 7.715 1.21 7.855 1.245 ;
 RECT 7.715 1.385 7.855 1.48 ;
 RECT 9.735 1.105 9.875 1.245 ;
 RECT 7.715 1.245 9.875 1.385 ;
 RECT 9.735 1.385 9.875 2.33 ;
 RECT 9.43 0.76 9.57 0.965 ;
 RECT 9.43 0.965 9.875 1.105 ;
 RECT 6.025 1.35 6.165 2.1 ;
 RECT 6.025 2.24 6.165 2.295 ;
 RECT 5.085 2.295 6.165 2.435 ;
 RECT 7.525 2.32 7.665 2.52 ;
 RECT 6.025 2.18 7.595 2.185 ;
 RECT 6.025 2.185 7.665 2.24 ;
 RECT 6.58 0.5 7.37 0.64 ;
 RECT 6.88 2.24 7.665 2.32 ;
 RECT 6.025 2.1 7.02 2.18 ;
 RECT 6.58 0.64 6.72 1.21 ;
 RECT 6.025 1.21 6.72 1.35 ;
 RECT 2.325 2.515 5.225 2.655 ;
 RECT 5.085 2.435 5.225 2.515 ;
 RECT 1.885 0.825 2.025 1.135 ;
 RECT 1.805 1.925 1.945 1.99 ;
 RECT 1.805 2.13 1.945 2.35 ;
 RECT 2.325 2.49 2.465 2.515 ;
 RECT 1.885 1.135 2.27 1.275 ;
 RECT 2.13 1.275 2.27 1.99 ;
 RECT 1.735 1.99 2.27 2.13 ;
 RECT 1.805 2.35 2.465 2.49 ;
 RECT 7.525 2.52 9.02 2.66 ;
 RECT 5.68 1.015 6.415 1.05 ;
 RECT 5.68 1.05 5.82 1.185 ;
 RECT 5.07 1.185 5.82 1.325 ;
 RECT 5.68 1.325 5.82 2.01 ;
 RECT 5.62 0.91 6.415 1.015 ;
 RECT 5.62 0.875 5.89 0.91 ;
 RECT 3.675 1.52 5.21 1.66 ;
 RECT 5.07 1.325 5.21 1.52 ;
 RECT 5.63 2.01 5.885 2.15 ;
 RECT 0.58 1.195 1.7 1.335 ;
 RECT 1.56 0.67 1.7 1.195 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.05 ;
 RECT 0.58 2.05 1.015 2.19 ;
 RECT 0.58 0.87 1.015 1.01 ;
 RECT 1.56 0.53 2.51 0.67 ;
 RECT 2.37 0.22 3.13 0.36 ;
 RECT 2.99 0.36 3.13 0.875 ;
 RECT 3.005 1.015 3.145 2.035 ;
 RECT 2.945 2.035 3.145 2.17 ;
 RECT 2.945 2.17 3.085 2.305 ;
 RECT 2.37 0.36 2.51 0.53 ;
 RECT 2.925 0.875 3.2 1.015 ;
 RECT 7.875 2.1 8.06 2.22 ;
 RECT 8.705 2.065 8.845 2.22 ;
 RECT 7.83 1.96 8.06 2.1 ;
 RECT 7.875 2.22 8.845 2.36 ;
 RECT 3.285 1.82 5.49 1.945 ;
 RECT 3.285 1.945 4.595 1.96 ;
 RECT 4.31 1.805 5.49 1.82 ;
 RECT 3.285 1.22 3.6 1.36 ;
 RECT 3.46 0.805 3.6 1.22 ;
 RECT 3.37 1.96 3.65 2.215 ;
 RECT 5.35 1.56 5.49 1.805 ;
 RECT 3.285 1.36 3.425 1.82 ;
 RECT 2.595 1.385 2.735 1.82 ;
 RECT 2.465 1.825 2.785 1.96 ;
 RECT 2.465 1.82 2.735 1.825 ;
 RECT 2.645 1.96 2.785 2.345 ;
 RECT 2.595 0.84 2.735 1.155 ;
 RECT 2.595 1.155 2.865 1.385 ;
 RECT 6.935 1.005 7.075 1.685 ;
 RECT 6.425 1.685 7.075 1.81 ;
 RECT 6.425 1.81 7.115 1.825 ;
 RECT 6.845 1.825 7.115 1.95 ;
 RECT 6.865 0.865 7.145 1.005 ;
 RECT 7.405 1.675 9.595 1.815 ;
 RECT 9.295 1.815 9.595 1.935 ;
 RECT 9.02 1.565 9.595 1.675 ;
 RECT 9.455 1.935 9.595 2.505 ;
 RECT 10.015 1.92 10.155 2.505 ;
 RECT 9.455 2.505 10.155 2.645 ;
 RECT 7.405 0.805 7.545 1.675 ;
 RECT 7.405 1.815 7.615 1.895 ;
 RECT 8.31 1.815 8.54 2.055 ;
 RECT 7.335 1.895 7.615 2.035 ;
 RECT 10.25 1.45 10.39 1.78 ;
 RECT 10.015 1.78 10.39 1.92 ;
 RECT 10.25 1.215 10.595 1.45 ;
 END
END DFFNASRNX1

MACRO DFFNASRNX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.84 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.84 2.96 ;
 RECT 5.345 2.635 5.605 2.8 ;
 RECT 1.865 2.625 2.11 2.8 ;
 RECT 9.155 2.15 9.295 2.8 ;
 RECT 10.275 2.06 10.415 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.26 1.93 1.4 2.8 ;
 RECT 6.365 2.38 6.505 2.8 ;
 RECT 11.33 1.56 11.47 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.84 0.08 ;
 RECT 1.26 0.08 1.4 1.055 ;
 RECT 1.96 0.08 2.19 0.39 ;
 RECT 4.605 0.08 4.84 0.37 ;
 RECT 8.625 0.08 8.88 1.005 ;
 RECT 10.295 0.08 10.435 0.725 ;
 RECT 0.28 0.08 0.42 0.775 ;
 RECT 11.33 0.08 11.47 0.885 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.275 1.475 1.575 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4 0.51 5.155 0.65 ;
 RECT 6.085 0.36 6.41 0.6 ;
 RECT 5.015 0.36 5.155 0.51 ;
 RECT 9.12 1.155 9.575 1.185 ;
 RECT 8.345 1.185 9.575 1.295 ;
 RECT 8.345 0.36 8.485 1.185 ;
 RECT 5.015 0.22 8.485 0.36 ;
 RECT 8.345 1.295 9.26 1.325 ;
 END
 ANTENNAGATEAREA 0.117 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.865 0.5 8.17 0.74 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.585 2.085 11 2.405 ;
 RECT 10.86 2.405 11 2.62 ;
 RECT 10.86 0.69 11 2.085 ;
 END
 ANTENNADIFFAREA 0.676 ;
 END QN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.31 1.16 0.805 1.49 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END D

 OBS
 LAYER PO ;
 RECT 1.335 1.48 1.62 1.72 ;
 RECT 1.52 1.72 1.62 2.37 ;
 RECT 8.95 1.53 9.51 1.63 ;
 RECT 9.285 1.63 9.51 1.94 ;
 RECT 8.95 0.65 9.05 1.53 ;
 RECT 9.41 1.94 9.51 2.695 ;
 RECT 6.125 0.865 6.52 1.095 ;
 RECT 6.42 1.095 6.52 1.64 ;
 RECT 6.42 1.64 6.655 1.87 ;
 RECT 3.675 1.33 3.815 1.475 ;
 RECT 3.675 1.71 3.775 2.475 ;
 RECT 3.715 0.65 3.815 1.33 ;
 RECT 3.675 1.475 3.905 1.71 ;
 RECT 4.115 0.695 4.215 1.61 ;
 RECT 4.15 1.71 4.25 2.48 ;
 RECT 4.115 1.61 4.25 1.71 ;
 RECT 3.995 0.465 4.235 0.695 ;
 RECT 4.975 1.79 5.075 2.685 ;
 RECT 2.6 2.12 2.81 2.685 ;
 RECT 2.6 2.685 5.075 2.785 ;
 RECT 5.75 1.33 5.85 1.565 ;
 RECT 6.14 1.665 6.24 2.69 ;
 RECT 8.115 0.74 8.215 2.69 ;
 RECT 8.115 0.495 8.215 0.5 ;
 RECT 7.935 0.5 8.215 0.74 ;
 RECT 5.23 0.635 5.33 1.23 ;
 RECT 5.23 1.23 5.85 1.33 ;
 RECT 5.75 1.565 6.24 1.665 ;
 RECT 6.14 2.69 8.215 2.79 ;
 RECT 6.7 0.56 6.8 1.35 ;
 RECT 8.455 0.265 8.555 1.32 ;
 RECT 5.715 0.56 5.945 0.69 ;
 RECT 5.715 0.46 6.8 0.56 ;
 RECT 6.7 0.265 6.8 0.46 ;
 RECT 7.145 1.545 7.245 2.495 ;
 RECT 6.7 0.165 8.555 0.265 ;
 RECT 6.7 1.35 6.99 1.445 ;
 RECT 6.7 1.445 7.245 1.45 ;
 RECT 6.89 1.45 7.245 1.545 ;
 RECT 0.6 1.185 1.145 1.425 ;
 RECT 1.045 0.655 1.145 1.185 ;
 RECT 1.045 1.425 1.145 2.685 ;
 RECT 10.36 1.125 10.71 1.19 ;
 RECT 10.36 1.29 10.71 1.355 ;
 RECT 10.61 0.21 10.71 1.125 ;
 RECT 10.61 1.355 10.71 2.79 ;
 RECT 10.36 1.19 11.215 1.29 ;
 RECT 11.115 0.21 11.215 1.19 ;
 RECT 11.115 1.29 11.215 2.79 ;
 RECT 8.725 2.47 9.04 2.71 ;
 RECT 8.94 1.95 9.04 2.47 ;
 RECT 9.97 1.345 10.07 2.69 ;
 RECT 9.39 0.635 9.49 1.105 ;
 RECT 9.32 1.105 9.55 1.245 ;
 RECT 9.32 1.245 10.07 1.345 ;
 RECT 5.28 1.61 5.545 1.82 ;
 RECT 5.445 1.82 5.545 2.52 ;
 RECT 4.875 0.625 4.975 1.51 ;
 RECT 4.875 1.51 5.545 1.61 ;
 RECT 1.86 1.52 2.46 1.62 ;
 RECT 2.32 1.645 3.28 1.745 ;
 RECT 2.32 1.62 2.46 1.645 ;
 RECT 2.36 0.285 2.46 1.52 ;
 RECT 2.32 1.745 2.42 2.355 ;
 RECT 4.415 0.285 4.515 1.24 ;
 RECT 2.36 0.185 4.515 0.285 ;
 RECT 1.86 1.44 2.105 1.52 ;
 RECT 1.86 1.62 2.105 1.69 ;
 RECT 3.18 1.745 3.28 2.495 ;
 RECT 3.18 1.615 3.28 1.645 ;
 RECT 7.64 0.645 7.74 1.24 ;
 RECT 7.64 1.24 7.885 1.45 ;
 RECT 7.64 1.45 7.74 2.37 ;
 RECT 7.17 0.685 7.27 1.255 ;
 RECT 7.095 0.455 7.325 0.685 ;
 RECT 2.655 1.155 3.325 1.31 ;
 RECT 2.655 1.31 2.9 1.465 ;
 RECT 3.225 0.47 3.51 0.705 ;
 RECT 3.225 0.705 3.325 1.155 ;
 RECT 1.52 0.655 1.62 1.48 ;
 LAYER CO ;
 RECT 8.79 2.525 8.92 2.655 ;
 RECT 10.865 1.605 10.995 1.735 ;
 RECT 10.865 1.865 10.995 1.995 ;
 RECT 6.195 0.915 6.325 1.045 ;
 RECT 9.37 1.16 9.5 1.29 ;
 RECT 8.7 0.87 8.83 1 ;
 RECT 11.335 0.665 11.465 0.795 ;
 RECT 11.335 1.61 11.465 1.74 ;
 RECT 5.765 0.51 5.895 0.64 ;
 RECT 4.375 1.825 4.505 1.955 ;
 RECT 3.895 2.105 4.025 2.235 ;
 RECT 1.92 1.495 2.05 1.625 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 8.69 2.19 8.82 2.32 ;
 RECT 10.28 2.13 10.41 2.26 ;
 RECT 9.72 2.13 9.85 2.26 ;
 RECT 9.335 1.76 9.465 1.89 ;
 RECT 5.335 1.63 5.465 1.76 ;
 RECT 1.87 0.875 2 1.005 ;
 RECT 5.665 2.015 5.795 2.145 ;
 RECT 2.01 0.255 2.14 0.385 ;
 RECT 5.395 2.64 5.525 2.77 ;
 RECT 4.725 2.125 4.855 2.255 ;
 RECT 10.865 0.765 10.995 0.895 ;
 RECT 10.865 2.15 10.995 2.28 ;
 RECT 10.865 2.41 10.995 2.54 ;
 RECT 2.58 1.87 2.71 2 ;
 RECT 3.33 0.525 3.46 0.655 ;
 RECT 7.39 1.825 7.52 1.955 ;
 RECT 0.285 0.59 0.415 0.72 ;
 RECT 0.285 0.33 0.415 0.46 ;
 RECT 7.145 0.505 7.275 0.635 ;
 RECT 7.7 1.28 7.83 1.41 ;
 RECT 9.785 0.87 9.915 1 ;
 RECT 9.16 2.2 9.29 2.33 ;
 RECT 2.93 2.105 3.06 2.235 ;
 RECT 2.975 0.88 3.105 1.01 ;
 RECT 2.71 1.28 2.84 1.41 ;
 RECT 2.58 0.905 2.71 1.035 ;
 RECT 1.385 1.535 1.515 1.665 ;
 RECT 1.74 1.995 1.87 2.125 ;
 RECT 1.265 1.995 1.395 2.125 ;
 RECT 1.265 0.875 1.395 1.005 ;
 RECT 0.795 2.095 0.925 2.225 ;
 RECT 10.3 0.525 10.43 0.655 ;
 RECT 6.475 1.69 6.605 1.82 ;
 RECT 0.645 1.245 0.775 1.375 ;
 RECT 4.05 0.515 4.18 0.645 ;
 RECT 4.655 0.235 4.785 0.365 ;
 RECT 7.39 0.87 7.52 1 ;
 RECT 8.34 1.925 8.47 2.055 ;
 RECT 7.86 2.04 7.99 2.17 ;
 RECT 6.92 0.87 7.05 1 ;
 RECT 1.925 2.63 2.055 2.76 ;
 RECT 2.64 2.175 2.77 2.305 ;
 RECT 3.425 2.07 3.555 2.2 ;
 RECT 3.445 0.88 3.575 1.01 ;
 RECT 7.995 0.55 8.125 0.68 ;
 RECT 3.725 1.525 3.855 1.655 ;
 RECT 5.67 0.88 5.8 1.01 ;
 RECT 6.895 1.815 7.025 1.945 ;
 RECT 6.37 2.44 6.5 2.57 ;
 RECT 10.41 1.175 10.54 1.305 ;
 RECT 0.785 0.875 0.915 1.005 ;
 RECT 11.335 1.87 11.465 2 ;
 RECT 11.335 2.155 11.465 2.285 ;
 RECT 11.335 2.415 11.465 2.545 ;
 LAYER M1 ;
 RECT 3.825 2.12 4.925 2.24 ;
 RECT 3.825 2.1 4.095 2.12 ;
 RECT 3.89 2.24 4.925 2.26 ;
 RECT 5.66 1.325 5.8 2.01 ;
 RECT 5.66 1.05 5.8 1.185 ;
 RECT 5.05 1.185 5.8 1.325 ;
 RECT 5.66 1.015 6.395 1.05 ;
 RECT 3.655 1.52 5.19 1.66 ;
 RECT 5.05 1.325 5.19 1.52 ;
 RECT 5.61 2.01 5.865 2.15 ;
 RECT 5.6 0.875 6.395 1.015 ;
 RECT 7.695 1.21 7.835 1.475 ;
 RECT 9.715 1.615 9.855 2.325 ;
 RECT 7.695 1.475 9.92 1.615 ;
 RECT 9.78 0.8 9.92 1.475 ;
 RECT 3.26 0.52 3.86 0.66 ;
 RECT 3.72 0.66 3.86 0.79 ;
 RECT 5.295 0.505 5.945 0.645 ;
 RECT 3.72 0.79 5.435 0.93 ;
 RECT 5.295 0.645 5.435 0.79 ;
 RECT 2.575 1.23 2.845 1.46 ;
 RECT 2.575 0.84 2.715 1.23 ;
 RECT 2.575 1.46 2.775 2.375 ;
 RECT 7.81 2.22 8.825 2.36 ;
 RECT 7.81 2.035 8.04 2.22 ;
 RECT 8.685 2.14 8.825 2.22 ;
 RECT 8.685 2.36 8.825 2.375 ;
 RECT 0.98 1.01 1.12 1.195 ;
 RECT 0.98 1.335 1.12 1.945 ;
 RECT 0.79 2.085 0.93 2.305 ;
 RECT 0.715 0.87 1.12 1.01 ;
 RECT 0.79 1.945 1.12 2.085 ;
 RECT 1.54 0.67 1.68 1.195 ;
 RECT 0.98 1.195 1.68 1.335 ;
 RECT 1.54 0.53 3.11 0.67 ;
 RECT 2.97 0.67 3.11 0.975 ;
 RECT 2.985 1.09 3.125 2.005 ;
 RECT 2.92 2.005 3.125 2.295 ;
 RECT 2.97 0.975 3.125 1.09 ;
 RECT 6.005 1.35 6.145 2.1 ;
 RECT 6.005 2.24 6.145 2.295 ;
 RECT 5.065 2.295 6.145 2.435 ;
 RECT 7.505 2.32 7.645 2.52 ;
 RECT 6.005 2.18 7.645 2.24 ;
 RECT 6.56 0.5 7.35 0.64 ;
 RECT 6.86 2.24 7.645 2.32 ;
 RECT 6.005 2.1 7 2.18 ;
 RECT 6.56 0.64 6.7 1.21 ;
 RECT 6.005 1.21 6.7 1.35 ;
 RECT 2.25 2.52 5.205 2.66 ;
 RECT 5.065 2.435 5.205 2.52 ;
 RECT 1.735 1.63 1.875 2.245 ;
 RECT 1.735 1.475 2.125 1.63 ;
 RECT 1.865 0.825 2.005 1.475 ;
 RECT 2.25 2.385 2.39 2.52 ;
 RECT 1.735 2.245 2.39 2.385 ;
 RECT 7.505 2.52 9 2.66 ;
 RECT 3.265 1.82 5.47 1.96 ;
 RECT 3.35 1.96 3.63 2.215 ;
 RECT 3.44 0.805 3.58 1.22 ;
 RECT 3.265 1.22 3.58 1.36 ;
 RECT 5.33 1.56 5.47 1.82 ;
 RECT 3.265 1.36 3.405 1.82 ;
 RECT 6.405 1.685 7.125 1.825 ;
 RECT 6.825 1.825 7.125 1.95 ;
 RECT 6.915 1.005 7.125 1.685 ;
 RECT 6.845 0.865 7.125 1.005 ;
 RECT 8.29 1.895 8.52 2.06 ;
 RECT 7.315 1.895 7.595 1.96 ;
 RECT 7.385 0.805 7.525 1.755 ;
 RECT 7.315 1.82 9.575 1.895 ;
 RECT 7.385 1.755 9.575 1.82 ;
 RECT 9.995 1.92 10.135 2.505 ;
 RECT 9.435 2.505 10.135 2.645 ;
 RECT 9.435 1.895 9.575 2.505 ;
 RECT 10.23 1.31 10.37 1.78 ;
 RECT 9.995 1.78 10.37 1.92 ;
 RECT 10.23 1.17 10.61 1.31 ;
 END
END DFFNASRNX2

MACRO DFFNASRQX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.2 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.2 2.96 ;
 RECT 1.935 2.635 2.185 2.8 ;
 RECT 5.365 2.635 5.625 2.8 ;
 RECT 10.295 2.06 10.435 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 6.385 2.38 6.525 2.8 ;
 RECT 1.28 1.98 1.42 2.8 ;
 RECT 9.175 2.085 9.315 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.2 0.08 ;
 RECT 1.91 0.08 2.21 0.26 ;
 RECT 1.28 0.08 1.42 1.055 ;
 RECT 4.625 0.08 4.86 0.26 ;
 RECT 8.645 0.08 8.9 0.285 ;
 RECT 10.315 0.08 10.455 0.785 ;
 RECT 0.3 0.08 0.44 0.775 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.58 1.475 1.91 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.02 0.51 5.175 0.65 ;
 RECT 9.06 0.28 9.34 0.42 ;
 RECT 5.94 0.36 6.2 0.6 ;
 RECT 5.035 0.22 8.46 0.225 ;
 RECT 5.035 0.225 8.505 0.36 ;
 RECT 8.365 0.46 9.275 0.6 ;
 RECT 9.135 0.22 9.275 0.28 ;
 RECT 8.365 0.36 8.505 0.46 ;
 RECT 5.035 0.36 5.175 0.51 ;
 RECT 9.06 0.42 9.275 0.46 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.92 1.475 1.275 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.87 0.5 8.195 0.79 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SETB

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.88 2.08 11.02 2.35 ;
 RECT 10.575 1.76 11.02 2.08 ;
 RECT 10.88 0.55 11.02 1.76 ;
 END
 ANTENNADIFFAREA 0.533 ;
 END Q

 OBS
 LAYER PO ;
 RECT 7.66 1.45 7.76 2.37 ;
 RECT 7.19 0.685 7.29 1.255 ;
 RECT 7.115 0.455 7.345 0.685 ;
 RECT 10.38 1.17 10.73 1.4 ;
 RECT 10.63 0.16 10.73 1.17 ;
 RECT 10.63 1.4 10.73 2.775 ;
 RECT 2.72 2.33 2.82 2.685 ;
 RECT 4.995 1.79 5.095 2.685 ;
 RECT 2.6 2.09 2.82 2.33 ;
 RECT 2.72 2.685 5.095 2.785 ;
 RECT 3.695 1.33 3.835 1.475 ;
 RECT 3.695 1.71 3.795 2.475 ;
 RECT 3.735 0.65 3.835 1.33 ;
 RECT 3.695 1.475 3.925 1.71 ;
 RECT 1.065 0.635 1.165 1.495 ;
 RECT 1.065 1.725 1.165 2.465 ;
 RECT 0.985 1.495 1.205 1.725 ;
 RECT 2.065 1.44 2.48 1.585 ;
 RECT 2.065 1.585 3.3 1.685 ;
 RECT 3.2 1.685 3.3 2.495 ;
 RECT 2.315 1.69 2.415 2.27 ;
 RECT 2.065 1.685 2.415 1.69 ;
 RECT 4.435 0.285 4.535 1.24 ;
 RECT 2.7 0.185 4.535 0.285 ;
 RECT 2.38 0.685 2.48 1.44 ;
 RECT 2.7 0.285 2.8 0.585 ;
 RECT 2.38 0.585 2.8 0.685 ;
 RECT 6.72 0.685 6.82 1.35 ;
 RECT 7.165 1.545 7.265 2.43 ;
 RECT 8.475 0.265 8.575 1.32 ;
 RECT 5.53 0.455 5.76 0.585 ;
 RECT 6.72 0.265 6.82 0.585 ;
 RECT 5.53 0.585 6.82 0.685 ;
 RECT 6.72 0.165 8.575 0.265 ;
 RECT 6.91 1.45 7.265 1.545 ;
 RECT 6.72 1.35 7.01 1.445 ;
 RECT 6.72 1.445 7.265 1.45 ;
 RECT 8.745 2.47 9.06 2.71 ;
 RECT 8.96 1.83 9.06 2.47 ;
 RECT 4.135 0.695 4.235 1.61 ;
 RECT 4.17 1.71 4.27 2.48 ;
 RECT 4.135 1.61 4.27 1.71 ;
 RECT 4.015 0.465 4.255 0.695 ;
 RECT 1.54 0.655 1.64 1.48 ;
 RECT 1.54 1.48 1.85 1.72 ;
 RECT 1.54 1.72 1.64 2.37 ;
 RECT 5.77 1.33 5.87 1.565 ;
 RECT 6.16 1.665 6.26 2.69 ;
 RECT 8.135 0.76 8.235 2.69 ;
 RECT 7.94 0.635 8.235 0.76 ;
 RECT 7.94 0.52 8.17 0.635 ;
 RECT 5.25 0.635 5.35 1.23 ;
 RECT 5.25 1.23 5.87 1.33 ;
 RECT 5.77 1.565 6.26 1.665 ;
 RECT 6.16 2.69 8.235 2.79 ;
 RECT 3.245 0.705 3.345 1.21 ;
 RECT 3.245 0.47 3.53 0.705 ;
 RECT 2.675 1.16 2.92 1.21 ;
 RECT 2.675 1.31 2.92 1.405 ;
 RECT 2.675 1.21 3.345 1.31 ;
 RECT 6.145 0.865 6.54 1.095 ;
 RECT 6.44 1.095 6.54 1.64 ;
 RECT 6.44 1.64 6.675 1.87 ;
 RECT 9.99 1.32 10.09 2.545 ;
 RECT 9.215 0.47 9.315 1.22 ;
 RECT 9.215 1.22 10.09 1.32 ;
 RECT 9.085 0.23 9.315 0.47 ;
 RECT 9.305 1.63 9.53 1.94 ;
 RECT 9.43 1.94 9.53 2.56 ;
 RECT 8.915 0.65 9.015 1.53 ;
 RECT 8.915 1.53 9.53 1.63 ;
 RECT 5.3 1.61 5.565 1.82 ;
 RECT 5.465 1.82 5.565 2.49 ;
 RECT 4.895 0.625 4.995 1.51 ;
 RECT 4.895 1.51 5.565 1.61 ;
 RECT 7.66 0.645 7.76 1.24 ;
 RECT 7.66 1.24 7.905 1.45 ;
 LAYER CO ;
 RECT 8.81 2.525 8.94 2.655 ;
 RECT 6.915 1.815 7.045 1.945 ;
 RECT 6.39 2.44 6.52 2.57 ;
 RECT 3.445 2.07 3.575 2.2 ;
 RECT 3.465 0.88 3.595 1.01 ;
 RECT 2.95 2.105 3.08 2.235 ;
 RECT 6.495 1.69 6.625 1.82 ;
 RECT 4.395 1.82 4.525 1.95 ;
 RECT 3.915 2.105 4.045 2.235 ;
 RECT 2.135 1.495 2.265 1.625 ;
 RECT 1.285 0.875 1.415 1.005 ;
 RECT 0.815 0.875 0.945 1.005 ;
 RECT 0.815 2.055 0.945 2.185 ;
 RECT 7.41 0.87 7.54 1 ;
 RECT 8.36 1.92 8.49 2.05 ;
 RECT 2.6 0.905 2.73 1.035 ;
 RECT 1.68 1.535 1.81 1.665 ;
 RECT 1.81 1.995 1.94 2.125 ;
 RECT 1.89 0.875 2.02 1.005 ;
 RECT 1.285 2.05 1.415 2.18 ;
 RECT 3.35 0.525 3.48 0.655 ;
 RECT 5.355 1.63 5.485 1.76 ;
 RECT 2.535 1.825 2.665 1.955 ;
 RECT 5.415 2.64 5.545 2.77 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 8 0.58 8.13 0.71 ;
 RECT 1.025 1.545 1.155 1.675 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 10.43 1.22 10.56 1.35 ;
 RECT 10.885 0.615 11.015 0.745 ;
 RECT 10.885 1.87 11.015 2 ;
 RECT 10.885 2.13 11.015 2.26 ;
 RECT 10.32 0.58 10.45 0.71 ;
 RECT 2.005 2.64 2.135 2.77 ;
 RECT 4.07 0.515 4.2 0.645 ;
 RECT 4.675 0.12 4.805 0.25 ;
 RECT 5.58 0.505 5.71 0.635 ;
 RECT 7.41 1.9 7.54 2.03 ;
 RECT 2.995 0.88 3.125 1.01 ;
 RECT 2.73 1.205 2.86 1.335 ;
 RECT 6.215 0.915 6.345 1.045 ;
 RECT 9.135 0.285 9.265 0.415 ;
 RECT 8.72 0.15 8.85 0.28 ;
 RECT 9.18 2.17 9.31 2.3 ;
 RECT 8.71 2.135 8.84 2.265 ;
 RECT 10.3 2.17 10.43 2.3 ;
 RECT 9.74 2.17 9.87 2.3 ;
 RECT 9.355 1.735 9.485 1.865 ;
 RECT 2.65 2.145 2.78 2.275 ;
 RECT 7.88 1.965 8.01 2.095 ;
 RECT 6.94 0.87 7.07 1 ;
 RECT 7.165 0.505 7.295 0.635 ;
 RECT 7.72 1.28 7.85 1.41 ;
 RECT 9.435 0.87 9.565 1 ;
 RECT 4.745 2.125 4.875 2.255 ;
 RECT 3.745 1.525 3.875 1.655 ;
 RECT 5.69 0.88 5.82 1.01 ;
 RECT 5.685 2.015 5.815 2.145 ;
 RECT 2.03 0.125 2.16 0.255 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 LAYER M1 ;
 RECT 3.845 2.12 4.945 2.24 ;
 RECT 3.845 2.1 4.115 2.12 ;
 RECT 3.91 2.24 4.945 2.26 ;
 RECT 3.28 0.52 3.88 0.66 ;
 RECT 3.74 0.66 3.88 0.79 ;
 RECT 3.74 0.79 5.455 0.93 ;
 RECT 5.315 0.5 5.76 0.64 ;
 RECT 5.315 0.64 5.455 0.79 ;
 RECT 5.68 1.325 5.82 2.01 ;
 RECT 5.68 1.05 5.82 1.185 ;
 RECT 5.07 1.185 5.82 1.325 ;
 RECT 5.62 0.91 6.415 1.015 ;
 RECT 5.62 0.875 5.89 0.91 ;
 RECT 5.68 1.015 6.415 1.05 ;
 RECT 3.675 1.52 5.21 1.66 ;
 RECT 5.07 1.325 5.21 1.52 ;
 RECT 5.63 2.01 5.885 2.15 ;
 RECT 7.715 1.21 7.855 1.395 ;
 RECT 9.735 1.105 9.875 1.34 ;
 RECT 7.715 1.48 9.875 1.535 ;
 RECT 9.735 1.535 9.875 2.365 ;
 RECT 9.43 0.76 9.57 0.965 ;
 RECT 9.43 0.965 9.875 1.105 ;
 RECT 7.715 1.395 10.565 1.48 ;
 RECT 9.735 1.34 10.565 1.395 ;
 RECT 10.425 1.15 10.565 1.34 ;
 RECT 6.025 1.35 6.165 2.1 ;
 RECT 6.025 2.24 6.165 2.295 ;
 RECT 5.085 2.295 6.165 2.435 ;
 RECT 7.525 2.32 7.665 2.52 ;
 RECT 6.025 2.18 7.595 2.185 ;
 RECT 6.025 2.185 7.665 2.24 ;
 RECT 6.88 2.24 7.665 2.32 ;
 RECT 6.025 2.1 7.02 2.18 ;
 RECT 6.58 0.5 7.37 0.64 ;
 RECT 6.025 1.21 6.72 1.35 ;
 RECT 6.58 0.64 6.72 1.21 ;
 RECT 2.325 2.515 5.225 2.655 ;
 RECT 5.085 2.435 5.225 2.515 ;
 RECT 1.885 0.825 2.025 1.125 ;
 RECT 1.805 2.13 1.945 2.35 ;
 RECT 2.325 2.49 2.465 2.515 ;
 RECT 1.885 1.125 2.27 1.265 ;
 RECT 2.13 1.265 2.27 1.99 ;
 RECT 1.735 1.99 2.27 2.13 ;
 RECT 1.805 2.35 2.465 2.49 ;
 RECT 7.525 2.52 9.02 2.66 ;
 RECT 2.595 1.385 2.735 1.82 ;
 RECT 2.465 1.825 2.785 1.96 ;
 RECT 2.465 1.82 2.735 1.825 ;
 RECT 2.645 1.96 2.785 2.345 ;
 RECT 2.595 0.84 2.735 1.155 ;
 RECT 2.595 1.155 2.865 1.385 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.05 ;
 RECT 0.58 2.05 1.015 2.19 ;
 RECT 0.58 0.87 1.015 1.01 ;
 RECT 0.58 1.195 1.7 1.335 ;
 RECT 1.56 0.67 1.7 1.195 ;
 RECT 1.56 0.53 2.51 0.67 ;
 RECT 2.37 0.22 3.13 0.36 ;
 RECT 2.99 0.36 3.13 0.875 ;
 RECT 2.945 2.035 3.145 2.17 ;
 RECT 2.945 2.17 3.085 2.305 ;
 RECT 3.005 1.015 3.145 2.035 ;
 RECT 2.37 0.36 2.51 0.53 ;
 RECT 2.925 0.875 3.2 1.015 ;
 RECT 3.285 1.82 5.49 1.945 ;
 RECT 3.285 1.945 4.595 1.96 ;
 RECT 4.31 1.805 5.49 1.82 ;
 RECT 3.285 1.22 3.6 1.36 ;
 RECT 3.46 0.805 3.6 1.22 ;
 RECT 3.37 1.96 3.65 2.215 ;
 RECT 5.35 1.56 5.49 1.805 ;
 RECT 3.285 1.36 3.425 1.82 ;
 RECT 7.875 2.1 8.06 2.22 ;
 RECT 8.705 2.065 8.845 2.22 ;
 RECT 7.875 2.22 8.845 2.36 ;
 RECT 7.83 1.96 8.06 2.1 ;
 RECT 7.405 1.675 9.525 1.815 ;
 RECT 7.405 0.805 7.545 1.675 ;
 RECT 7.405 1.815 7.615 1.895 ;
 RECT 8.31 1.815 8.54 2.055 ;
 RECT 9.295 1.815 9.525 1.935 ;
 RECT 7.335 1.895 7.615 2.035 ;
 RECT 6.935 1.005 7.075 1.685 ;
 RECT 6.425 1.685 7.075 1.81 ;
 RECT 6.425 1.81 7.115 1.825 ;
 RECT 6.845 1.825 7.115 1.95 ;
 RECT 6.865 0.865 7.145 1.005 ;
 END
END DFFNASRQX1

MACRO DFFNASRQX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.84 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.84 2.96 ;
 RECT 1.865 2.625 2.11 2.8 ;
 RECT 5.345 2.635 5.605 2.8 ;
 RECT 10.275 2.06 10.415 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.26 1.93 1.4 2.8 ;
 RECT 6.365 2.38 6.505 2.8 ;
 RECT 11.33 1.56 11.47 2.8 ;
 RECT 9.155 2.15 9.295 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.84 0.08 ;
 RECT 8.625 0.08 8.88 1.005 ;
 RECT 1.26 0.08 1.4 1.055 ;
 RECT 4.605 0.08 4.84 0.37 ;
 RECT 1.96 0.08 2.19 0.39 ;
 RECT 10.295 0.08 10.435 0.96 ;
 RECT 0.28 0.08 0.42 0.775 ;
 RECT 11.33 0.08 11.47 0.955 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.275 1.475 1.575 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4 0.51 5.155 0.65 ;
 RECT 6.085 0.36 6.41 0.46 ;
 RECT 5.015 0.36 5.155 0.51 ;
 RECT 9.12 1.155 9.575 1.185 ;
 RECT 8.275 1.185 9.575 1.295 ;
 RECT 8.275 0.36 8.415 1.185 ;
 RECT 5.015 0.22 8.415 0.36 ;
 RECT 8.275 1.295 9.26 1.325 ;
 END
 ANTENNAGATEAREA 0.117 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.87 0.5 8.135 0.815 ;
 END
 ANTENNAGATEAREA 0.098 ;
 END SETB

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.585 2.085 11 2.405 ;
 RECT 10.86 2.405 11 2.62 ;
 RECT 10.86 0.69 11 2.085 ;
 END
 ANTENNADIFFAREA 0.596 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.31 1.16 0.805 1.49 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 10.36 1.29 10.71 1.355 ;
 RECT 10.61 0.42 10.71 1.125 ;
 RECT 10.61 1.355 10.71 2.79 ;
 RECT 10.36 1.19 11.215 1.29 ;
 RECT 11.115 0.42 11.215 1.19 ;
 RECT 11.115 1.29 11.215 2.79 ;
 RECT 2.32 1.65 3.28 1.75 ;
 RECT 1.86 1.52 2.46 1.62 ;
 RECT 2.32 1.62 2.46 1.65 ;
 RECT 2.36 0.285 2.46 1.52 ;
 RECT 2.32 1.75 2.42 2.355 ;
 RECT 4.415 0.285 4.515 1.24 ;
 RECT 3.18 1.75 3.28 2.495 ;
 RECT 2.36 0.185 4.515 0.285 ;
 RECT 1.86 1.44 2.105 1.52 ;
 RECT 1.86 1.62 2.105 1.69 ;
 RECT 7.64 0.645 7.74 1.24 ;
 RECT 7.64 1.24 7.885 1.45 ;
 RECT 7.64 1.45 7.74 2.37 ;
 RECT 7.17 0.685 7.27 1.255 ;
 RECT 7.095 0.455 7.325 0.685 ;
 RECT 2.655 1.155 3.325 1.31 ;
 RECT 2.655 1.31 2.9 1.47 ;
 RECT 3.225 0.47 3.51 0.705 ;
 RECT 3.225 0.705 3.325 1.155 ;
 RECT 5.28 1.61 5.545 1.82 ;
 RECT 5.445 1.82 5.545 2.49 ;
 RECT 4.875 0.625 4.975 1.51 ;
 RECT 4.875 1.51 5.545 1.61 ;
 RECT 3.675 1.33 3.815 1.475 ;
 RECT 3.675 1.71 3.775 2.475 ;
 RECT 3.715 0.65 3.815 1.33 ;
 RECT 3.675 1.475 3.905 1.71 ;
 RECT 2.6 2.12 2.81 2.685 ;
 RECT 4.975 1.79 5.075 2.685 ;
 RECT 2.6 2.685 5.075 2.785 ;
 RECT 0.6 1.185 1.145 1.425 ;
 RECT 1.045 0.655 1.145 1.185 ;
 RECT 1.045 1.425 1.145 2.465 ;
 RECT 4.115 0.695 4.215 1.61 ;
 RECT 4.15 1.71 4.25 2.48 ;
 RECT 4.115 1.61 4.25 1.71 ;
 RECT 3.995 0.465 4.235 0.695 ;
 RECT 6.7 0.265 6.8 0.46 ;
 RECT 5.715 0.46 6.8 0.56 ;
 RECT 6.7 0.56 6.8 1.35 ;
 RECT 7.145 1.545 7.245 2.38 ;
 RECT 8.455 0.265 8.555 1.32 ;
 RECT 5.715 0.56 5.945 0.69 ;
 RECT 6.89 1.45 7.245 1.545 ;
 RECT 6.7 1.35 6.99 1.445 ;
 RECT 6.7 1.445 7.245 1.45 ;
 RECT 6.7 0.165 8.555 0.265 ;
 RECT 1.52 0.655 1.62 1.48 ;
 RECT 1.335 1.48 1.62 1.72 ;
 RECT 1.52 1.72 1.62 2.37 ;
 RECT 9.97 1.345 10.07 2.69 ;
 RECT 9.39 0.635 9.49 1.105 ;
 RECT 9.32 1.105 9.55 1.245 ;
 RECT 9.32 1.245 10.07 1.345 ;
 RECT 5.75 1.33 5.85 1.565 ;
 RECT 6.14 1.665 6.24 2.69 ;
 RECT 6.705 2.63 6.935 2.69 ;
 RECT 8.115 0.76 8.215 2.69 ;
 RECT 7.925 0.54 8.215 0.76 ;
 RECT 5.23 0.635 5.33 1.23 ;
 RECT 5.23 1.23 5.85 1.33 ;
 RECT 5.75 1.565 6.24 1.665 ;
 RECT 6.14 2.69 8.215 2.79 ;
 RECT 8.725 2.47 9.04 2.71 ;
 RECT 8.94 1.95 9.04 2.47 ;
 RECT 8.95 1.53 9.51 1.63 ;
 RECT 9.285 1.63 9.51 1.94 ;
 RECT 8.95 0.65 9.05 1.53 ;
 RECT 9.41 1.94 9.51 2.695 ;
 RECT 6.125 0.865 6.52 1.095 ;
 RECT 6.42 1.095 6.52 1.64 ;
 RECT 6.42 1.64 6.655 1.87 ;
 RECT 10.36 1.125 10.71 1.19 ;
 LAYER CO ;
 RECT 2.01 0.255 2.14 0.385 ;
 RECT 5.395 2.64 5.525 2.77 ;
 RECT 10.865 1.605 10.995 1.735 ;
 RECT 10.865 1.865 10.995 1.995 ;
 RECT 10.865 2.15 10.995 2.28 ;
 RECT 10.865 2.41 10.995 2.54 ;
 RECT 10.3 0.745 10.43 0.875 ;
 RECT 0.645 1.245 0.775 1.375 ;
 RECT 2.58 1.87 2.71 2 ;
 RECT 3.33 0.525 3.46 0.655 ;
 RECT 7.7 1.28 7.83 1.41 ;
 RECT 9.785 0.87 9.915 1 ;
 RECT 9.16 2.2 9.29 2.33 ;
 RECT 8.69 2.19 8.82 2.32 ;
 RECT 10.28 2.13 10.41 2.26 ;
 RECT 7.975 0.58 8.105 0.71 ;
 RECT 1.74 1.995 1.87 2.125 ;
 RECT 1.87 0.875 2 1.005 ;
 RECT 1.265 1.995 1.395 2.125 ;
 RECT 1.265 0.875 1.395 1.005 ;
 RECT 0.795 2.095 0.925 2.225 ;
 RECT 6.37 2.44 6.5 2.57 ;
 RECT 10.41 1.175 10.54 1.305 ;
 RECT 6.195 0.915 6.325 1.045 ;
 RECT 9.37 1.16 9.5 1.29 ;
 RECT 11.335 0.73 11.465 0.86 ;
 RECT 11.335 1.61 11.465 1.74 ;
 RECT 11.335 1.87 11.465 2 ;
 RECT 11.335 2.155 11.465 2.285 ;
 RECT 11.335 2.415 11.465 2.545 ;
 RECT 4.375 1.825 4.505 1.955 ;
 RECT 3.895 2.105 4.025 2.235 ;
 RECT 1.92 1.495 2.05 1.625 ;
 RECT 6.92 0.87 7.05 1 ;
 RECT 7.145 0.505 7.275 0.635 ;
 RECT 0.285 0.59 0.415 0.72 ;
 RECT 0.285 0.33 0.415 0.46 ;
 RECT 3.425 2.07 3.555 2.2 ;
 RECT 3.445 0.88 3.575 1.01 ;
 RECT 2.93 2.105 3.06 2.235 ;
 RECT 2.975 0.88 3.105 1.01 ;
 RECT 9.72 2.13 9.85 2.26 ;
 RECT 9.335 1.76 9.465 1.89 ;
 RECT 8.79 2.525 8.92 2.655 ;
 RECT 6.895 1.815 7.025 1.945 ;
 RECT 4.725 2.125 4.855 2.255 ;
 RECT 0.785 0.875 0.915 1.005 ;
 RECT 6.475 1.69 6.605 1.82 ;
 RECT 1.925 2.63 2.055 2.76 ;
 RECT 2.64 2.175 2.77 2.305 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 2.71 1.28 2.84 1.41 ;
 RECT 2.58 0.905 2.71 1.035 ;
 RECT 1.385 1.535 1.515 1.665 ;
 RECT 5.335 1.63 5.465 1.76 ;
 RECT 3.725 1.525 3.855 1.655 ;
 RECT 5.67 0.88 5.8 1.01 ;
 RECT 5.665 2.015 5.795 2.145 ;
 RECT 10.865 0.765 10.995 0.895 ;
 RECT 8.7 0.87 8.83 1 ;
 RECT 4.05 0.515 4.18 0.645 ;
 RECT 4.655 0.235 4.785 0.365 ;
 RECT 5.765 0.51 5.895 0.64 ;
 RECT 7.39 1.825 7.52 1.955 ;
 RECT 7.39 0.87 7.52 1 ;
 RECT 8.34 1.925 8.47 2.055 ;
 RECT 7.86 2.04 7.99 2.17 ;
 LAYER M1 ;
 RECT 3.825 2.12 4.925 2.24 ;
 RECT 3.825 2.1 4.095 2.12 ;
 RECT 3.89 2.24 4.925 2.26 ;
 RECT 7.695 1.21 7.835 1.475 ;
 RECT 9.78 1.31 9.92 1.475 ;
 RECT 7.695 1.475 9.92 1.615 ;
 RECT 9.715 1.615 9.855 2.325 ;
 RECT 9.78 0.8 9.92 1.17 ;
 RECT 9.78 1.17 10.61 1.31 ;
 RECT 3.26 0.52 3.86 0.66 ;
 RECT 3.72 0.66 3.86 0.79 ;
 RECT 5.295 0.505 5.945 0.645 ;
 RECT 3.72 0.79 5.435 0.93 ;
 RECT 5.295 0.645 5.435 0.79 ;
 RECT 5.66 1.325 5.8 2.01 ;
 RECT 5.66 1.05 5.8 1.185 ;
 RECT 5.05 1.185 5.8 1.325 ;
 RECT 5.66 1.015 6.395 1.05 ;
 RECT 3.655 1.52 5.19 1.66 ;
 RECT 5.05 1.325 5.19 1.52 ;
 RECT 5.61 2.01 5.865 2.15 ;
 RECT 5.6 0.875 6.395 1.015 ;
 RECT 6.005 1.35 6.145 2.1 ;
 RECT 6.005 2.24 6.145 2.295 ;
 RECT 5.065 2.295 6.145 2.435 ;
 RECT 2.25 2.52 5.205 2.66 ;
 RECT 5.065 2.435 5.205 2.52 ;
 RECT 7.505 2.32 7.645 2.52 ;
 RECT 6.005 2.18 7.645 2.24 ;
 RECT 6.56 0.5 7.35 0.64 ;
 RECT 6.86 2.24 7.645 2.32 ;
 RECT 6.005 2.1 7 2.18 ;
 RECT 6.56 0.64 6.7 1.21 ;
 RECT 6.005 1.21 6.7 1.35 ;
 RECT 1.735 1.63 1.875 2.245 ;
 RECT 1.735 1.475 2.125 1.63 ;
 RECT 1.865 0.825 2.005 1.475 ;
 RECT 2.25 2.385 2.39 2.52 ;
 RECT 1.735 2.245 2.39 2.385 ;
 RECT 7.505 2.52 9 2.66 ;
 RECT 3.265 1.82 5.47 1.96 ;
 RECT 3.265 1.22 3.58 1.36 ;
 RECT 3.44 0.805 3.58 1.22 ;
 RECT 3.35 1.96 3.63 2.215 ;
 RECT 5.33 1.56 5.47 1.82 ;
 RECT 3.265 1.36 3.405 1.82 ;
 RECT 2.575 1.23 2.845 1.46 ;
 RECT 2.575 0.84 2.715 1.23 ;
 RECT 2.575 1.46 2.775 2.375 ;
 RECT 0.98 1.01 1.12 1.195 ;
 RECT 0.98 1.335 1.12 1.945 ;
 RECT 0.79 2.085 0.93 2.305 ;
 RECT 0.715 0.87 1.12 1.01 ;
 RECT 0.79 1.945 1.12 2.085 ;
 RECT 1.54 0.67 1.68 1.195 ;
 RECT 0.98 1.195 1.68 1.335 ;
 RECT 1.54 0.53 3.11 0.67 ;
 RECT 2.97 0.67 3.11 0.975 ;
 RECT 2.92 2.005 3.125 2.295 ;
 RECT 2.985 1.09 3.125 2.005 ;
 RECT 2.97 0.975 3.125 1.09 ;
 RECT 7.315 1.895 7.595 1.96 ;
 RECT 7.385 0.805 7.525 1.755 ;
 RECT 8.29 1.895 8.52 2.06 ;
 RECT 7.315 1.82 9.575 1.895 ;
 RECT 7.385 1.755 9.575 1.82 ;
 RECT 6.405 1.685 7.125 1.825 ;
 RECT 6.915 1.005 7.125 1.685 ;
 RECT 6.825 1.825 7.125 1.95 ;
 RECT 6.845 0.865 7.125 1.005 ;
 RECT 7.81 2.035 8.04 2.22 ;
 RECT 8.685 2.14 8.825 2.22 ;
 RECT 8.685 2.36 8.825 2.375 ;
 RECT 7.81 2.22 8.825 2.36 ;
 END
END DFFNASRQX2

MACRO DFFNASRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 12.16 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 12.16 2.96 ;
 RECT 1.935 2.635 2.185 2.8 ;
 RECT 5.365 2.635 5.625 2.8 ;
 RECT 1.28 1.98 1.42 2.8 ;
 RECT 9.175 2.085 9.315 2.8 ;
 RECT 10.295 2.06 10.435 2.8 ;
 RECT 11.82 1.73 11.96 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 6.385 2.38 6.525 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 12.16 0.08 ;
 RECT 8.645 0.08 8.9 0.285 ;
 RECT 1.91 0.08 2.21 0.26 ;
 RECT 4.625 0.08 4.86 0.26 ;
 RECT 1.28 0.08 1.42 1.055 ;
 RECT 11.905 0.08 12.045 0.88 ;
 RECT 10.315 0.08 10.455 0.725 ;
 RECT 0.3 0.08 0.44 0.775 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.58 1.475 1.91 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.36 0.36 8.5 0.5 ;
 RECT 4.02 0.51 5.175 0.65 ;
 RECT 9.06 0.28 9.34 0.49 ;
 RECT 5.955 0.36 6.205 0.6 ;
 RECT 5.035 0.22 8.5 0.36 ;
 RECT 5.035 0.36 5.175 0.51 ;
 RECT 8.36 0.635 9.17 0.64 ;
 RECT 9.06 0.49 9.21 0.5 ;
 RECT 8.36 0.5 9.21 0.635 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.92 1.475 1.275 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.88 0.5 8.17 0.765 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.88 1.425 11.02 2.35 ;
 RECT 10.88 1.105 11.19 1.425 ;
 RECT 10.88 0.55 11.02 1.105 ;
 END
 ANTENNADIFFAREA 0.633 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.17 2.015 11.485 2.38 ;
 RECT 11.345 0.7 11.485 2.015 ;
 END
 ANTENNADIFFAREA 0.495 ;
 END Q

 OBS
 LAYER PO ;
 RECT 2.065 1.44 2.48 1.585 ;
 RECT 2.065 1.585 3.3 1.685 ;
 RECT 2.065 1.685 2.415 1.69 ;
 RECT 2.315 1.69 2.415 2.27 ;
 RECT 4.435 0.285 4.535 1.24 ;
 RECT 2.7 0.185 4.535 0.285 ;
 RECT 2.38 0.685 2.48 1.44 ;
 RECT 2.7 0.285 2.8 0.585 ;
 RECT 3.2 1.685 3.3 2.495 ;
 RECT 2.38 0.585 2.8 0.685 ;
 RECT 4.135 0.695 4.235 1.61 ;
 RECT 4.17 1.71 4.27 2.48 ;
 RECT 4.135 1.61 4.27 1.71 ;
 RECT 4.015 0.465 4.255 0.695 ;
 RECT 6.72 0.265 6.82 0.585 ;
 RECT 5.535 0.585 6.82 0.685 ;
 RECT 6.72 0.685 6.82 1.35 ;
 RECT 7.165 1.545 7.265 2.405 ;
 RECT 8.475 0.265 8.575 1.32 ;
 RECT 5.535 0.455 5.765 0.585 ;
 RECT 6.91 1.45 7.265 1.545 ;
 RECT 6.72 0.165 8.575 0.265 ;
 RECT 6.72 1.35 7.01 1.445 ;
 RECT 6.72 1.445 7.265 1.45 ;
 RECT 8.745 2.47 9.06 2.71 ;
 RECT 8.96 1.83 9.06 2.47 ;
 RECT 3.245 0.705 3.345 1.21 ;
 RECT 2.675 1.16 2.92 1.21 ;
 RECT 2.675 1.21 3.345 1.31 ;
 RECT 2.675 1.31 2.92 1.405 ;
 RECT 3.245 0.47 3.53 0.705 ;
 RECT 9.99 1.32 10.09 2.545 ;
 RECT 9.215 0.47 9.315 1.22 ;
 RECT 9.215 1.22 10.09 1.32 ;
 RECT 9.085 0.23 9.315 0.47 ;
 RECT 5.77 1.33 5.87 1.565 ;
 RECT 6.16 1.665 6.26 2.69 ;
 RECT 8.135 0.735 8.235 2.69 ;
 RECT 7.94 0.535 8.235 0.735 ;
 RECT 7.94 0.515 8.17 0.535 ;
 RECT 5.25 0.635 5.35 1.23 ;
 RECT 5.25 1.23 5.87 1.33 ;
 RECT 5.77 1.565 6.26 1.665 ;
 RECT 6.16 2.69 8.235 2.79 ;
 RECT 1.54 0.655 1.64 1.48 ;
 RECT 1.54 1.48 1.85 1.72 ;
 RECT 1.54 1.72 1.64 2.37 ;
 RECT 6.145 0.865 6.54 1.095 ;
 RECT 6.44 1.095 6.54 1.64 ;
 RECT 6.44 1.64 6.675 1.87 ;
 RECT 9.305 1.63 9.53 1.94 ;
 RECT 9.43 1.94 9.53 2.56 ;
 RECT 8.915 0.65 9.015 1.53 ;
 RECT 8.915 1.53 9.53 1.63 ;
 RECT 1.065 0.635 1.165 1.495 ;
 RECT 1.065 1.725 1.165 2.465 ;
 RECT 0.985 1.495 1.205 1.725 ;
 RECT 7.66 0.645 7.76 1.24 ;
 RECT 7.66 1.24 7.905 1.45 ;
 RECT 7.66 1.45 7.76 2.37 ;
 RECT 7.19 0.685 7.29 1.255 ;
 RECT 7.115 0.455 7.345 0.685 ;
 RECT 5.3 1.61 5.565 1.82 ;
 RECT 5.465 1.82 5.565 2.49 ;
 RECT 4.895 0.625 4.995 1.51 ;
 RECT 4.895 1.51 5.565 1.61 ;
 RECT 3.695 1.33 3.835 1.475 ;
 RECT 3.695 1.71 3.795 2.475 ;
 RECT 3.735 0.65 3.835 1.33 ;
 RECT 3.695 1.475 3.925 1.71 ;
 RECT 4.995 1.79 5.095 2.685 ;
 RECT 2.72 2.33 2.82 2.685 ;
 RECT 2.72 2.685 5.095 2.785 ;
 RECT 2.6 2.09 2.82 2.33 ;
 RECT 10.38 1.12 10.73 1.35 ;
 RECT 10.63 0.165 10.73 1.12 ;
 RECT 10.63 1.35 10.73 2.79 ;
 RECT 11.605 0.28 11.705 1.1 ;
 RECT 11.605 1.335 11.705 2.79 ;
 RECT 11.59 1.1 11.8 1.335 ;
 LAYER CO ;
 RECT 3.745 1.525 3.875 1.655 ;
 RECT 5.69 0.88 5.82 1.01 ;
 RECT 5.685 2.015 5.815 2.145 ;
 RECT 2.03 0.125 2.16 0.255 ;
 RECT 10.885 1.87 11.015 2 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 2.995 0.88 3.125 1.01 ;
 RECT 2.73 1.205 2.86 1.335 ;
 RECT 2.6 0.905 2.73 1.035 ;
 RECT 9.435 0.87 9.565 1 ;
 RECT 8.81 2.525 8.94 2.655 ;
 RECT 1.82 1.995 1.95 2.125 ;
 RECT 10.43 1.18 10.56 1.31 ;
 RECT 0.815 0.875 0.945 1.005 ;
 RECT 11.825 1.8 11.955 1.93 ;
 RECT 11.825 2.06 11.955 2.19 ;
 RECT 4.745 2.125 4.875 2.255 ;
 RECT 3.35 0.525 3.48 0.655 ;
 RECT 6.495 1.69 6.625 1.82 ;
 RECT 6.215 0.915 6.345 1.045 ;
 RECT 4.395 1.82 4.525 1.95 ;
 RECT 3.915 2.105 4.045 2.235 ;
 RECT 2.135 1.495 2.265 1.625 ;
 RECT 2.005 2.64 2.135 2.77 ;
 RECT 3.445 2.07 3.575 2.2 ;
 RECT 8.36 1.92 8.49 2.05 ;
 RECT 7.88 1.965 8.01 2.095 ;
 RECT 6.94 0.87 7.07 1 ;
 RECT 7.165 0.505 7.295 0.635 ;
 RECT 7.99 0.565 8.12 0.695 ;
 RECT 1.68 1.535 1.81 1.665 ;
 RECT 9.18 2.17 9.31 2.3 ;
 RECT 8.71 2.135 8.84 2.265 ;
 RECT 10.3 2.13 10.43 2.26 ;
 RECT 6.915 1.815 7.045 1.945 ;
 RECT 6.39 2.44 6.52 2.57 ;
 RECT 11.63 1.15 11.76 1.28 ;
 RECT 11.91 0.68 12.04 0.81 ;
 RECT 11.35 1.65 11.48 1.78 ;
 RECT 11.35 1.91 11.48 2.04 ;
 RECT 11.35 2.17 11.48 2.3 ;
 RECT 11.825 2.32 11.955 2.45 ;
 RECT 11.35 0.75 11.48 0.88 ;
 RECT 5.415 2.64 5.545 2.77 ;
 RECT 2.535 1.825 2.665 1.955 ;
 RECT 10.885 2.13 11.015 2.26 ;
 RECT 10.32 0.505 10.45 0.635 ;
 RECT 3.465 0.88 3.595 1.01 ;
 RECT 2.95 2.105 3.08 2.235 ;
 RECT 7.72 1.28 7.85 1.41 ;
 RECT 1.89 0.875 2.02 1.005 ;
 RECT 1.285 2.05 1.415 2.18 ;
 RECT 1.285 0.875 1.415 1.005 ;
 RECT 9.74 2.13 9.87 2.26 ;
 RECT 9.355 1.76 9.485 1.89 ;
 RECT 5.355 1.63 5.485 1.76 ;
 RECT 0.815 2.055 0.945 2.185 ;
 RECT 2.65 2.145 2.78 2.275 ;
 RECT 10.885 0.615 11.015 0.745 ;
 RECT 1.025 1.545 1.155 1.675 ;
 RECT 9.135 0.285 9.265 0.415 ;
 RECT 8.72 0.15 8.85 0.28 ;
 RECT 4.07 0.515 4.2 0.645 ;
 RECT 4.675 0.12 4.805 0.25 ;
 RECT 5.585 0.505 5.715 0.635 ;
 RECT 7.41 1.9 7.54 2.03 ;
 RECT 7.41 0.87 7.54 1 ;
 LAYER M1 ;
 RECT 3.845 2.12 4.945 2.24 ;
 RECT 3.845 2.1 4.115 2.12 ;
 RECT 3.91 2.24 4.945 2.26 ;
 RECT 5.68 1.325 5.82 2.01 ;
 RECT 5.68 1.05 5.82 1.185 ;
 RECT 5.07 1.185 5.82 1.325 ;
 RECT 5.62 0.91 6.415 1.015 ;
 RECT 5.62 0.875 5.89 0.91 ;
 RECT 5.68 1.015 6.415 1.05 ;
 RECT 3.675 1.52 5.21 1.66 ;
 RECT 5.07 1.325 5.21 1.52 ;
 RECT 5.63 2.01 5.885 2.15 ;
 RECT 3.28 0.52 3.88 0.66 ;
 RECT 3.74 0.66 3.88 0.79 ;
 RECT 3.74 0.79 5.475 0.93 ;
 RECT 5.335 0.5 5.765 0.64 ;
 RECT 5.335 0.64 5.475 0.79 ;
 RECT 9.735 1.105 9.875 1.395 ;
 RECT 9.735 1.535 9.875 2.33 ;
 RECT 7.715 1.395 9.875 1.535 ;
 RECT 9.43 1.005 9.875 1.105 ;
 RECT 9.43 0.76 9.57 0.965 ;
 RECT 7.715 1.21 7.855 1.395 ;
 RECT 10.595 0.36 10.735 0.865 ;
 RECT 9.43 0.965 10.735 1.005 ;
 RECT 9.735 0.865 10.735 0.965 ;
 RECT 10.595 0.22 11.59 0.36 ;
 RECT 11.625 0.56 11.765 1.36 ;
 RECT 11.45 0.36 11.59 0.42 ;
 RECT 11.45 0.42 11.765 0.56 ;
 RECT 6.425 1.685 7.075 1.81 ;
 RECT 6.935 1.005 7.075 1.685 ;
 RECT 6.425 1.81 7.115 1.825 ;
 RECT 6.845 1.825 7.115 1.95 ;
 RECT 6.865 0.865 7.145 1.005 ;
 RECT 6.025 1.35 6.165 2.1 ;
 RECT 6.025 2.24 6.165 2.295 ;
 RECT 5.085 2.295 6.165 2.435 ;
 RECT 2.325 2.515 5.225 2.655 ;
 RECT 5.085 2.435 5.225 2.515 ;
 RECT 1.815 1.925 1.955 1.95 ;
 RECT 1.815 2.18 1.955 2.35 ;
 RECT 2.325 2.49 2.465 2.515 ;
 RECT 1.885 0.825 2.025 1.135 ;
 RECT 1.735 1.95 1.99 1.99 ;
 RECT 1.735 2.13 1.99 2.18 ;
 RECT 1.885 1.135 2.27 1.275 ;
 RECT 1.815 2.35 2.465 2.49 ;
 RECT 2.13 1.275 2.27 1.99 ;
 RECT 1.735 1.99 2.27 2.13 ;
 RECT 7.525 2.32 7.665 2.52 ;
 RECT 6.025 2.18 7.595 2.185 ;
 RECT 6.025 2.185 7.665 2.24 ;
 RECT 6.58 0.5 7.37 0.64 ;
 RECT 6.88 2.24 7.665 2.32 ;
 RECT 6.025 2.1 7.02 2.18 ;
 RECT 6.58 0.64 6.72 1.21 ;
 RECT 6.025 1.21 6.72 1.35 ;
 RECT 7.525 2.52 9.02 2.66 ;
 RECT 2.595 1.385 2.735 1.82 ;
 RECT 2.465 1.825 2.785 1.96 ;
 RECT 2.465 1.82 2.735 1.825 ;
 RECT 2.645 1.96 2.785 2.345 ;
 RECT 2.595 0.84 2.735 1.155 ;
 RECT 2.595 1.155 2.865 1.385 ;
 RECT 3.285 1.82 5.49 1.945 ;
 RECT 3.285 1.945 4.595 1.96 ;
 RECT 4.31 1.805 5.49 1.82 ;
 RECT 3.285 1.22 3.6 1.36 ;
 RECT 3.46 0.805 3.6 1.22 ;
 RECT 3.37 1.96 3.65 2.215 ;
 RECT 5.35 1.56 5.49 1.805 ;
 RECT 3.285 1.36 3.425 1.82 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.05 ;
 RECT 0.58 2.05 1.015 2.19 ;
 RECT 0.58 0.87 1.015 1.01 ;
 RECT 0.58 1.195 1.7 1.335 ;
 RECT 1.56 0.67 1.7 1.195 ;
 RECT 1.56 0.53 2.51 0.67 ;
 RECT 2.37 0.22 3.13 0.36 ;
 RECT 2.99 0.36 3.13 0.875 ;
 RECT 3.005 1.015 3.145 2.035 ;
 RECT 2.945 2.035 3.145 2.17 ;
 RECT 2.945 2.17 3.085 2.305 ;
 RECT 2.37 0.36 2.51 0.53 ;
 RECT 2.925 0.875 3.2 1.015 ;
 RECT 7.405 1.675 9.595 1.815 ;
 RECT 10.015 1.92 10.155 2.505 ;
 RECT 9.295 1.815 9.595 1.935 ;
 RECT 9.455 1.935 9.595 2.505 ;
 RECT 9.455 2.505 10.155 2.645 ;
 RECT 7.405 1.815 7.615 1.895 ;
 RECT 7.405 0.805 7.545 1.675 ;
 RECT 8.31 1.815 8.54 2.055 ;
 RECT 7.335 1.895 7.615 2.035 ;
 RECT 10.25 1.315 10.39 1.78 ;
 RECT 10.25 1.175 10.63 1.315 ;
 RECT 10.015 1.78 10.39 1.92 ;
 RECT 7.875 2.1 8.06 2.22 ;
 RECT 8.705 2.065 8.845 2.22 ;
 RECT 7.83 1.96 8.06 2.1 ;
 RECT 7.875 2.22 8.845 2.36 ;
 END
END DFFNASRX1

MACRO DFFNASRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 12.8 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 12.8 2.96 ;
 RECT 5.345 2.635 5.605 2.8 ;
 RECT 1.83 2.62 2.105 2.8 ;
 RECT 6.365 2.38 6.505 2.8 ;
 RECT 11.33 1.56 11.47 2.8 ;
 RECT 9.155 2.15 9.295 2.8 ;
 RECT 10.275 2.06 10.415 2.8 ;
 RECT 12.28 1.52 12.42 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.26 1.93 1.4 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 12.8 0.08 ;
 RECT 8.625 0.08 8.88 1.005 ;
 RECT 4.605 0.08 4.84 0.37 ;
 RECT 1.26 0.08 1.4 1.055 ;
 RECT 1.96 0.08 2.19 0.39 ;
 RECT 12.555 0.08 12.695 0.94 ;
 RECT 11.535 0.08 11.675 0.885 ;
 RECT 10.295 0.08 10.435 0.725 ;
 RECT 0.28 0.08 0.42 0.775 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.275 1.475 1.575 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4 0.51 5.155 0.65 ;
 RECT 5.92 0.36 6.245 0.63 ;
 RECT 5.015 0.22 8.46 0.36 ;
 RECT 5.015 0.36 5.155 0.51 ;
 RECT 8.32 1.325 8.46 1.33 ;
 RECT 9.12 1.155 9.575 1.185 ;
 RECT 8.32 1.185 9.575 1.295 ;
 RECT 8.32 0.36 8.46 1.185 ;
 RECT 8.32 1.295 9.26 1.325 ;
 END
 ANTENNAGATEAREA 0.117 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.85 0.5 8.18 0.785 ;
 END
 ANTENNAGATEAREA 0.098 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.585 2.085 11 2.405 ;
 RECT 10.86 2.405 11 2.62 ;
 RECT 10.86 0.69 11 2.085 ;
 END
 ANTENNADIFFAREA 0.676 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.805 2.015 12.135 2.38 ;
 RECT 11.805 1.025 12.225 1.165 ;
 RECT 11.805 2.38 11.945 2.61 ;
 RECT 12.085 0.675 12.225 1.025 ;
 RECT 11.805 1.165 11.945 2.015 ;
 END
 ANTENNADIFFAREA 0.55 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.31 1.15 0.805 1.49 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 12.065 1.29 12.165 2.79 ;
 RECT 11.48 1.29 11.69 1.425 ;
 RECT 11.59 1.425 11.69 2.79 ;
 RECT 12.34 0.36 12.44 1.19 ;
 RECT 1.045 0.655 1.145 1.185 ;
 RECT 1.045 1.425 1.145 2.465 ;
 RECT 0.6 1.185 1.145 1.425 ;
 RECT 3.675 1.33 3.815 1.475 ;
 RECT 3.675 1.71 3.775 2.475 ;
 RECT 3.715 0.65 3.815 1.33 ;
 RECT 3.675 1.475 3.905 1.71 ;
 RECT 10.61 0.21 10.71 1.125 ;
 RECT 10.36 1.125 10.71 1.19 ;
 RECT 10.61 1.355 10.71 2.79 ;
 RECT 10.36 1.29 10.71 1.355 ;
 RECT 10.36 1.19 11.215 1.29 ;
 RECT 11.115 0.21 11.215 1.19 ;
 RECT 11.115 1.29 11.215 2.79 ;
 RECT 6.235 1.64 6.655 1.87 ;
 RECT 6.235 1.095 6.44 1.64 ;
 RECT 6.125 0.865 6.44 1.095 ;
 RECT 9.97 1.345 10.07 2.69 ;
 RECT 9.39 0.635 9.49 1.105 ;
 RECT 9.32 1.105 9.55 1.245 ;
 RECT 9.32 1.245 10.07 1.345 ;
 RECT 4.115 0.695 4.215 1.61 ;
 RECT 4.15 1.71 4.25 2.48 ;
 RECT 4.115 1.61 4.25 1.71 ;
 RECT 3.995 0.465 4.235 0.695 ;
 RECT 7.64 0.645 7.74 1.24 ;
 RECT 7.64 1.24 7.885 1.45 ;
 RECT 7.64 1.45 7.74 2.37 ;
 RECT 7.17 0.685 7.27 1.255 ;
 RECT 7.095 0.455 7.325 0.685 ;
 RECT 8.95 1.53 9.51 1.63 ;
 RECT 9.285 1.63 9.51 1.94 ;
 RECT 9.41 1.94 9.51 2.695 ;
 RECT 8.95 0.65 9.05 1.53 ;
 RECT 3.225 0.47 3.51 0.705 ;
 RECT 3.225 0.705 3.325 1.165 ;
 RECT 2.64 1.265 2.885 1.405 ;
 RECT 2.64 1.165 3.325 1.265 ;
 RECT 5.28 1.61 5.545 1.82 ;
 RECT 5.445 1.82 5.545 2.49 ;
 RECT 4.875 0.625 4.975 1.51 ;
 RECT 4.875 1.51 5.545 1.61 ;
 RECT 6.7 0.265 6.8 0.58 ;
 RECT 6.7 0.68 6.8 1.35 ;
 RECT 8.455 0.265 8.555 1.32 ;
 RECT 5.51 0.46 5.74 0.58 ;
 RECT 5.51 0.68 5.74 0.69 ;
 RECT 5.51 0.58 6.8 0.68 ;
 RECT 7.145 1.545 7.245 2.38 ;
 RECT 6.7 0.165 8.555 0.265 ;
 RECT 6.7 1.35 6.99 1.445 ;
 RECT 6.7 1.445 7.245 1.45 ;
 RECT 6.89 1.45 7.245 1.545 ;
 RECT 1.86 1.52 2.46 1.59 ;
 RECT 2.36 0.285 2.46 1.52 ;
 RECT 3.18 1.69 3.28 2.495 ;
 RECT 1.86 1.59 3.28 1.62 ;
 RECT 2.285 1.62 3.28 1.69 ;
 RECT 4.415 0.285 4.515 1.24 ;
 RECT 2.36 0.185 4.515 0.285 ;
 RECT 2.285 1.69 2.385 2.225 ;
 RECT 1.86 1.44 2.105 1.52 ;
 RECT 1.86 1.62 2.105 1.69 ;
 RECT 1.52 0.655 1.62 1.48 ;
 RECT 1.335 1.48 1.62 1.72 ;
 RECT 1.52 1.72 1.62 2.37 ;
 RECT 4.975 1.79 5.075 2.685 ;
 RECT 2.565 2.09 2.81 2.685 ;
 RECT 2.565 2.685 5.075 2.785 ;
 RECT 5.75 1.33 5.85 1.565 ;
 RECT 5.955 1.665 6.055 2.69 ;
 RECT 8.115 0.745 8.215 2.69 ;
 RECT 7.93 0.635 8.215 0.745 ;
 RECT 7.93 0.515 8.16 0.635 ;
 RECT 5.23 0.635 5.33 1.23 ;
 RECT 5.23 1.23 5.85 1.33 ;
 RECT 5.75 1.565 6.055 1.665 ;
 RECT 5.955 2.69 8.215 2.79 ;
 RECT 8.725 2.47 9.04 2.71 ;
 RECT 8.94 1.95 9.04 2.47 ;
 RECT 11.48 1.19 12.44 1.29 ;
 RECT 11.87 0.395 11.97 1.19 ;
 LAYER CO ;
 RECT 2.58 1.81 2.71 1.94 ;
 RECT 3.33 0.525 3.46 0.655 ;
 RECT 0.285 0.59 0.415 0.72 ;
 RECT 0.285 0.33 0.415 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 7.99 0.565 8.12 0.695 ;
 RECT 4.05 0.515 4.18 0.645 ;
 RECT 4.655 0.235 4.785 0.365 ;
 RECT 8.34 1.925 8.47 2.055 ;
 RECT 7.86 2.04 7.99 2.17 ;
 RECT 6.92 0.87 7.05 1 ;
 RECT 6.895 1.815 7.025 1.945 ;
 RECT 6.37 2.44 6.5 2.57 ;
 RECT 7.7 1.28 7.83 1.41 ;
 RECT 9.785 0.87 9.915 1 ;
 RECT 9.16 2.2 9.29 2.33 ;
 RECT 12.09 0.75 12.22 0.88 ;
 RECT 10.41 1.175 10.54 1.305 ;
 RECT 9.72 2.13 9.85 2.26 ;
 RECT 9.335 1.76 9.465 1.89 ;
 RECT 5.335 1.63 5.465 1.76 ;
 RECT 3.725 1.525 3.855 1.655 ;
 RECT 5.67 0.88 5.8 1.01 ;
 RECT 5.665 2.015 5.795 2.145 ;
 RECT 2.01 0.255 2.14 0.385 ;
 RECT 5.395 2.64 5.525 2.77 ;
 RECT 4.725 2.125 4.855 2.255 ;
 RECT 11.335 2.155 11.465 2.285 ;
 RECT 11.335 2.415 11.465 2.545 ;
 RECT 4.375 1.825 4.505 1.955 ;
 RECT 1.915 2.625 2.045 2.755 ;
 RECT 2.93 2.105 3.06 2.235 ;
 RECT 2.975 0.88 3.105 1.01 ;
 RECT 2.695 1.23 2.825 1.36 ;
 RECT 1.385 1.535 1.515 1.665 ;
 RECT 1.74 1.995 1.87 2.125 ;
 RECT 1.87 0.875 2 1.005 ;
 RECT 1.265 1.995 1.395 2.125 ;
 RECT 1.265 0.875 1.395 1.005 ;
 RECT 0.795 2.095 0.925 2.225 ;
 RECT 2.62 2.135 2.75 2.265 ;
 RECT 12.285 1.605 12.415 1.735 ;
 RECT 12.285 1.865 12.415 1.995 ;
 RECT 12.285 2.15 12.415 2.28 ;
 RECT 12.285 2.41 12.415 2.54 ;
 RECT 11.81 1.605 11.94 1.735 ;
 RECT 10.865 1.605 10.995 1.735 ;
 RECT 10.865 1.865 10.995 1.995 ;
 RECT 0.785 0.875 0.915 1.005 ;
 RECT 0.645 1.245 0.775 1.375 ;
 RECT 11.81 1.865 11.94 1.995 ;
 RECT 11.81 2.15 11.94 2.28 ;
 RECT 11.81 2.41 11.94 2.54 ;
 RECT 8.79 2.525 8.92 2.655 ;
 RECT 11.52 1.24 11.65 1.37 ;
 RECT 12.56 0.74 12.69 0.87 ;
 RECT 10.865 0.765 10.995 0.895 ;
 RECT 10.865 2.15 10.995 2.28 ;
 RECT 10.865 2.41 10.995 2.54 ;
 RECT 10.3 0.525 10.43 0.655 ;
 RECT 6.475 1.69 6.605 1.82 ;
 RECT 6.195 0.915 6.325 1.045 ;
 RECT 9.37 1.16 9.5 1.29 ;
 RECT 8.7 0.87 8.83 1 ;
 RECT 11.54 0.665 11.67 0.795 ;
 RECT 11.335 1.61 11.465 1.74 ;
 RECT 11.335 1.87 11.465 2 ;
 RECT 5.56 0.51 5.69 0.64 ;
 RECT 7.39 1.825 7.52 1.955 ;
 RECT 7.39 0.87 7.52 1 ;
 RECT 3.895 2.105 4.025 2.235 ;
 RECT 1.92 1.495 2.05 1.625 ;
 RECT 7.145 0.505 7.275 0.635 ;
 RECT 3.425 2.07 3.555 2.2 ;
 RECT 3.445 0.88 3.575 1.01 ;
 RECT 8.69 2.19 8.82 2.32 ;
 RECT 10.28 2.13 10.41 2.26 ;
 RECT 2.58 0.905 2.71 1.035 ;
 LAYER M1 ;
 RECT 7.695 1.21 7.835 1.475 ;
 RECT 9.78 0.865 10.715 1.005 ;
 RECT 10.575 0.525 10.715 0.865 ;
 RECT 11.165 0.525 11.305 1.1 ;
 RECT 10.575 0.385 11.305 0.525 ;
 RECT 7.695 1.475 9.92 1.615 ;
 RECT 9.78 1.005 9.92 1.475 ;
 RECT 9.78 0.8 9.92 0.865 ;
 RECT 9.715 1.615 9.855 2.325 ;
 RECT 11.515 1.24 11.655 1.42 ;
 RECT 11.165 1.1 11.655 1.24 ;
 RECT 3.26 0.52 3.86 0.66 ;
 RECT 3.72 0.66 3.86 0.79 ;
 RECT 5.295 0.505 5.74 0.645 ;
 RECT 3.72 0.79 5.435 0.93 ;
 RECT 5.295 0.645 5.435 0.79 ;
 RECT 5.66 1.015 6.395 1.05 ;
 RECT 5.66 1.05 5.8 1.185 ;
 RECT 5.66 1.325 5.8 2.01 ;
 RECT 5.05 1.185 5.8 1.325 ;
 RECT 5.6 0.875 6.395 1.015 ;
 RECT 5.61 2.01 5.865 2.15 ;
 RECT 5.05 1.325 5.19 1.52 ;
 RECT 3.655 1.52 5.19 1.66 ;
 RECT 3.825 2.12 4.925 2.24 ;
 RECT 3.825 2.1 4.095 2.12 ;
 RECT 3.89 2.24 4.925 2.26 ;
 RECT 6.005 1.35 6.145 2.1 ;
 RECT 6.005 2.24 6.145 2.295 ;
 RECT 5.065 2.295 6.145 2.435 ;
 RECT 7.505 2.32 7.645 2.52 ;
 RECT 6.005 2.18 7.645 2.24 ;
 RECT 6.56 0.5 7.35 0.64 ;
 RECT 6.86 2.24 7.645 2.32 ;
 RECT 6.005 2.1 7 2.18 ;
 RECT 6.56 0.64 6.7 1.21 ;
 RECT 6.005 1.21 6.7 1.35 ;
 RECT 2.245 2.52 5.205 2.66 ;
 RECT 5.065 2.435 5.205 2.52 ;
 RECT 2.245 2.48 2.385 2.52 ;
 RECT 1.735 1.63 1.875 2.34 ;
 RECT 1.735 1.475 2.125 1.63 ;
 RECT 1.865 0.825 2.005 1.475 ;
 RECT 1.735 2.34 2.385 2.48 ;
 RECT 7.505 2.52 9 2.66 ;
 RECT 0.98 1.01 1.12 1.195 ;
 RECT 0.98 1.335 1.12 1.945 ;
 RECT 0.79 2.085 0.93 2.305 ;
 RECT 0.715 0.87 1.12 1.01 ;
 RECT 0.79 1.945 1.12 2.085 ;
 RECT 2.925 2.035 3.125 2.305 ;
 RECT 1.54 0.67 1.68 1.195 ;
 RECT 0.98 1.195 1.68 1.335 ;
 RECT 1.54 0.53 3.11 0.67 ;
 RECT 2.97 0.67 3.11 0.96 ;
 RECT 2.985 1.085 3.125 2.035 ;
 RECT 2.97 0.96 3.125 1.085 ;
 RECT 6.405 1.685 7.125 1.825 ;
 RECT 6.825 1.825 7.125 1.95 ;
 RECT 6.915 1.005 7.125 1.685 ;
 RECT 6.845 0.865 7.125 1.005 ;
 RECT 3.265 1.82 5.47 1.96 ;
 RECT 3.265 1.22 3.58 1.36 ;
 RECT 3.44 0.805 3.58 1.22 ;
 RECT 3.35 1.96 3.63 2.215 ;
 RECT 5.33 1.56 5.47 1.82 ;
 RECT 3.265 1.36 3.405 1.82 ;
 RECT 8.29 1.895 8.52 2.06 ;
 RECT 7.315 1.895 7.595 1.96 ;
 RECT 7.385 0.805 7.525 1.755 ;
 RECT 7.315 1.82 9.575 1.895 ;
 RECT 7.385 1.755 9.575 1.82 ;
 RECT 9.995 1.92 10.135 2.505 ;
 RECT 9.435 2.505 10.135 2.645 ;
 RECT 9.435 1.895 9.575 2.505 ;
 RECT 10.23 1.31 10.37 1.78 ;
 RECT 9.995 1.78 10.37 1.92 ;
 RECT 10.23 1.17 10.61 1.31 ;
 RECT 7.81 2.035 8.04 2.22 ;
 RECT 8.685 2.14 8.825 2.22 ;
 RECT 8.685 2.36 8.825 2.375 ;
 RECT 7.81 2.22 8.825 2.36 ;
 RECT 2.575 1.41 2.755 2.335 ;
 RECT 2.575 0.84 2.715 1.18 ;
 RECT 2.575 1.18 2.83 1.41 ;
 END
END DFFNASRX2

MACRO DFFNASX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.56 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.56 2.96 ;
 RECT 1.935 2.635 2.185 2.8 ;
 RECT 4.275 2.635 4.535 2.8 ;
 RECT 8.04 2.085 8.18 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 9.64 1.8 9.78 2.8 ;
 RECT 5.265 2.38 5.405 2.8 ;
 RECT 1.28 1.98 1.42 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.56 0.08 ;
 RECT 1.28 0.08 1.42 1.055 ;
 RECT 1.91 0.08 2.21 0.26 ;
 RECT 7.51 0.08 7.765 0.285 ;
 RECT 4.245 0.08 4.385 0.33 ;
 RECT 9.72 0.08 9.86 0.815 ;
 RECT 0.3 0.08 0.44 0.775 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.58 1.475 1.91 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.92 1.475 1.275 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.835 0.42 7.16 0.76 ;
 END
 ANTENNAGATEAREA 0.12 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.16 0.88 9.3 2.33 ;
 RECT 8.955 0.51 9.27 0.52 ;
 RECT 8.955 0.52 9.3 0.88 ;
 END
 ANTENNADIFFAREA 0.596 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.195 2.385 10.335 2.52 ;
 RECT 9.935 2.065 10.335 2.385 ;
 RECT 10.195 0.555 10.335 2.065 ;
 END
 ANTENNADIFFAREA 0.495 ;
 END Q

 OBS
 LAYER PO ;
 RECT 8.295 1.94 8.395 2.56 ;
 RECT 7.78 0.65 7.88 1.53 ;
 RECT 7.78 1.53 8.395 1.63 ;
 RECT 8.83 1.205 9.525 1.44 ;
 RECT 9.425 0.185 9.525 1.205 ;
 RECT 9.425 1.44 9.525 2.79 ;
 RECT 9.975 0.09 10.075 1.19 ;
 RECT 9.975 1.425 10.075 2.79 ;
 RECT 9.815 1.19 10.075 1.425 ;
 RECT 3.245 0.705 3.345 1.21 ;
 RECT 2.675 1.16 2.92 1.21 ;
 RECT 2.675 1.21 3.345 1.31 ;
 RECT 2.675 1.31 2.92 1.405 ;
 RECT 3.245 0.47 3.53 0.705 ;
 RECT 2.065 1.44 2.48 1.585 ;
 RECT 2.065 1.585 3.3 1.685 ;
 RECT 3.2 1.685 3.3 2.495 ;
 RECT 2.065 1.685 2.415 1.69 ;
 RECT 2.315 1.69 2.415 2.27 ;
 RECT 2.38 0.685 2.48 1.44 ;
 RECT 4.03 0.285 4.13 1.24 ;
 RECT 2.7 0.185 4.13 0.285 ;
 RECT 2.7 0.285 2.8 0.585 ;
 RECT 2.38 0.585 2.8 0.685 ;
 RECT 4.935 0.575 5.685 0.675 ;
 RECT 5.585 0.675 5.685 1.35 ;
 RECT 6.03 1.545 6.13 2.325 ;
 RECT 7.34 0.265 7.44 1.32 ;
 RECT 5.585 0.265 5.685 0.575 ;
 RECT 4.935 0.455 5.165 0.575 ;
 RECT 4.935 0.675 5.165 0.685 ;
 RECT 5.585 0.165 7.44 0.265 ;
 RECT 5.775 1.45 6.13 1.545 ;
 RECT 5.585 1.35 5.875 1.445 ;
 RECT 5.585 1.445 6.13 1.45 ;
 RECT 1.065 0.635 1.165 1.495 ;
 RECT 1.065 1.725 1.165 2.465 ;
 RECT 0.985 1.495 1.205 1.725 ;
 RECT 1.54 0.655 1.64 1.48 ;
 RECT 1.54 1.48 1.85 1.72 ;
 RECT 1.54 1.72 1.64 2.37 ;
 RECT 2.72 2.33 2.82 2.685 ;
 RECT 4 1.77 4.1 2.685 ;
 RECT 2.72 2.685 4.1 2.785 ;
 RECT 2.6 2.09 2.82 2.33 ;
 RECT 6.055 0.685 6.155 1.23 ;
 RECT 5.98 0.455 6.21 0.685 ;
 RECT 4.355 0.625 4.455 1.58 ;
 RECT 4.485 1.82 4.585 2.49 ;
 RECT 4.355 1.58 4.595 1.82 ;
 RECT 3.695 1.43 3.795 1.475 ;
 RECT 3.695 1.71 3.795 2.505 ;
 RECT 3.715 0.65 3.815 1.33 ;
 RECT 3.695 1.33 3.815 1.43 ;
 RECT 3.565 1.475 3.795 1.71 ;
 RECT 4.975 1.375 5.075 2.69 ;
 RECT 4.655 1.275 5.075 1.375 ;
 RECT 4.975 2.69 7.1 2.79 ;
 RECT 7 0.715 7.1 2.69 ;
 RECT 4.655 0.635 4.755 1.275 ;
 RECT 6.87 0.485 7.1 0.715 ;
 RECT 7.61 2.47 7.925 2.71 ;
 RECT 7.825 1.83 7.925 2.47 ;
 RECT 5.305 1.095 5.405 1.64 ;
 RECT 5.305 1.64 5.62 1.87 ;
 RECT 5.135 0.865 5.405 1.095 ;
 RECT 6.525 0.645 6.625 1.24 ;
 RECT 6.525 1.24 6.77 1.45 ;
 RECT 6.525 1.45 6.625 2.37 ;
 RECT 8.17 1.63 8.395 1.94 ;
 LAYER CO ;
 RECT 2.6 0.905 2.73 1.035 ;
 RECT 1.68 1.535 1.81 1.665 ;
 RECT 1.81 1.995 1.94 2.125 ;
 RECT 1.89 0.875 2.02 1.005 ;
 RECT 10.2 1.8 10.33 1.93 ;
 RECT 10.2 2.06 10.33 2.19 ;
 RECT 1.285 0.875 1.415 1.005 ;
 RECT 5.44 1.69 5.57 1.82 ;
 RECT 5.2 0.915 5.33 1.045 ;
 RECT 7.585 0.15 7.715 0.28 ;
 RECT 4.25 0.15 4.38 0.28 ;
 RECT 6.275 1.9 6.405 2.03 ;
 RECT 6.275 0.87 6.405 1 ;
 RECT 7.225 1.92 7.355 2.05 ;
 RECT 2.65 2.145 2.78 2.275 ;
 RECT 2.535 1.825 2.665 1.955 ;
 RECT 3.35 0.525 3.48 0.655 ;
 RECT 6.585 1.28 6.715 1.41 ;
 RECT 8 0.87 8.13 1 ;
 RECT 8.605 2.13 8.735 2.26 ;
 RECT 8.22 1.76 8.35 1.89 ;
 RECT 4.425 1.63 4.555 1.76 ;
 RECT 3.615 1.525 3.745 1.655 ;
 RECT 4.71 2.015 4.84 2.145 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 6.93 0.535 7.06 0.665 ;
 RECT 7.675 2.525 7.805 2.655 ;
 RECT 5.78 1.815 5.91 1.945 ;
 RECT 5.27 2.44 5.4 2.57 ;
 RECT 9.855 1.24 9.985 1.37 ;
 RECT 10.2 0.625 10.33 0.755 ;
 RECT 10.2 2.32 10.33 2.45 ;
 RECT 8.885 1.245 9.015 1.375 ;
 RECT 9.725 0.56 9.855 0.69 ;
 RECT 9.645 1.87 9.775 2 ;
 RECT 9.645 2.13 9.775 2.26 ;
 RECT 2.135 1.495 2.265 1.625 ;
 RECT 2.005 2.64 2.135 2.77 ;
 RECT 4.985 0.505 5.115 0.635 ;
 RECT 3.445 2.07 3.575 2.2 ;
 RECT 3.465 0.88 3.595 1.01 ;
 RECT 2.95 2.105 3.08 2.235 ;
 RECT 2.995 0.88 3.125 1.01 ;
 RECT 2.73 1.205 2.86 1.335 ;
 RECT 6.745 1.965 6.875 2.095 ;
 RECT 5.805 0.87 5.935 1 ;
 RECT 6.03 0.505 6.16 0.635 ;
 RECT 1.285 2.05 1.415 2.18 ;
 RECT 8.045 2.17 8.175 2.3 ;
 RECT 7.575 2.135 7.705 2.265 ;
 RECT 9.165 2.13 9.295 2.26 ;
 RECT 9.165 0.585 9.295 0.715 ;
 RECT 4.875 0.88 5.005 1.01 ;
 RECT 9.165 1.795 9.295 1.925 ;
 RECT 2.03 0.125 2.16 0.255 ;
 RECT 4.325 2.64 4.455 2.77 ;
 RECT 0.815 0.875 0.945 1.005 ;
 RECT 0.815 2.055 0.945 2.185 ;
 RECT 1.025 1.545 1.155 1.675 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 LAYER M1 ;
 RECT 6.58 1.21 6.72 1.395 ;
 RECT 7.93 0.965 8.74 1.005 ;
 RECT 8.295 1.005 8.74 1.105 ;
 RECT 7.93 0.865 8.435 0.965 ;
 RECT 8.6 0.37 8.74 0.965 ;
 RECT 8.6 1.105 8.74 1.395 ;
 RECT 6.58 1.395 8.74 1.535 ;
 RECT 8.6 1.535 8.74 2.33 ;
 RECT 9.44 0.37 9.58 1.235 ;
 RECT 8.6 0.23 9.58 0.37 ;
 RECT 9.85 1.175 9.99 1.235 ;
 RECT 9.85 1.375 9.99 1.44 ;
 RECT 9.44 1.235 9.995 1.375 ;
 RECT 3.91 2.355 5.125 2.495 ;
 RECT 4.985 2.24 5.125 2.355 ;
 RECT 4.985 1.36 5.125 2.1 ;
 RECT 1.885 0.825 2.025 1.125 ;
 RECT 1.805 2.13 1.945 2.35 ;
 RECT 2.325 2.49 2.465 2.515 ;
 RECT 2.325 2.515 4.05 2.655 ;
 RECT 1.885 1.125 2.27 1.265 ;
 RECT 2.13 1.265 2.27 1.99 ;
 RECT 1.735 1.99 2.27 2.13 ;
 RECT 1.805 2.35 2.465 2.49 ;
 RECT 3.91 2.495 4.05 2.515 ;
 RECT 6.39 2.32 6.53 2.52 ;
 RECT 5.52 0.5 6.235 0.64 ;
 RECT 5.52 0.64 5.66 1.22 ;
 RECT 4.985 2.1 5.885 2.18 ;
 RECT 4.985 2.18 6.53 2.24 ;
 RECT 5.745 2.24 6.53 2.32 ;
 RECT 4.985 1.22 5.66 1.36 ;
 RECT 6.39 2.52 7.885 2.66 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.05 ;
 RECT 0.58 2.05 1.015 2.19 ;
 RECT 0.58 0.87 1.015 1.01 ;
 RECT 0.58 1.195 1.7 1.335 ;
 RECT 1.56 0.67 1.7 1.195 ;
 RECT 1.56 0.53 2.51 0.67 ;
 RECT 2.37 0.22 3.13 0.36 ;
 RECT 2.99 0.36 3.13 0.875 ;
 RECT 3.005 1.015 3.145 2.035 ;
 RECT 2.945 2.035 3.145 2.17 ;
 RECT 2.945 2.17 3.085 2.305 ;
 RECT 2.37 0.36 2.51 0.53 ;
 RECT 2.925 0.875 3.2 1.015 ;
 RECT 3.285 1.805 4.56 1.945 ;
 RECT 3.285 1.945 3.65 1.96 ;
 RECT 3.285 1.22 3.6 1.36 ;
 RECT 3.46 0.805 3.6 1.22 ;
 RECT 3.37 1.96 3.65 2.215 ;
 RECT 3.285 1.36 3.425 1.805 ;
 RECT 4.42 1.56 4.56 1.805 ;
 RECT 6.74 2.1 6.925 2.22 ;
 RECT 7.57 2.065 7.71 2.22 ;
 RECT 6.695 1.96 6.925 2.1 ;
 RECT 6.74 2.22 7.71 2.36 ;
 RECT 5.43 1.685 5.94 1.81 ;
 RECT 5.8 0.78 5.94 1.685 ;
 RECT 5.43 1.825 5.57 1.895 ;
 RECT 5.43 1.615 5.57 1.685 ;
 RECT 5.43 1.81 5.98 1.825 ;
 RECT 5.71 1.825 5.98 1.95 ;
 RECT 6.27 0.805 6.41 1.675 ;
 RECT 6.27 1.815 6.48 1.895 ;
 RECT 7.175 1.815 7.405 2.055 ;
 RECT 6.2 1.895 6.48 2.035 ;
 RECT 6.27 1.675 8.46 1.815 ;
 RECT 8.16 1.815 8.46 1.935 ;
 RECT 8.32 1.935 8.46 2.505 ;
 RECT 8.88 1.175 9.02 2.505 ;
 RECT 8.32 2.505 9.02 2.645 ;
 RECT 2.595 1.385 2.735 1.82 ;
 RECT 2.465 1.825 2.785 1.96 ;
 RECT 2.465 1.82 2.735 1.825 ;
 RECT 2.645 1.96 2.785 2.345 ;
 RECT 2.595 0.84 2.735 1.155 ;
 RECT 2.595 1.155 2.865 1.385 ;
 RECT 4.705 1.04 5.38 1.05 ;
 RECT 4.14 0.91 5.38 1.04 ;
 RECT 4.14 0.9 5.01 0.91 ;
 RECT 4.705 1.08 4.845 2.2 ;
 RECT 4.705 1.05 5.01 1.08 ;
 RECT 3.565 1.52 4.28 1.66 ;
 RECT 4.87 0.81 5.01 0.9 ;
 RECT 4.14 1.04 4.28 1.52 ;
 RECT 3.28 0.52 5.19 0.66 ;
 RECT 4.905 0.47 5.19 0.52 ;
 END
END DFFNASX1

MACRO SDFFASX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 13.76 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 13.76 2.96 ;
 RECT 6.415 2.635 6.675 2.8 ;
 RECT 4.075 2.36 4.325 2.8 ;
 RECT 1.51 2.085 1.65 2.8 ;
 RECT 11.305 1.48 11.445 2.8 ;
 RECT 7.405 2.38 7.545 2.8 ;
 RECT 12.25 1.48 12.39 2.8 ;
 RECT 13.22 1.435 13.36 2.8 ;
 RECT 3.42 2 3.56 2.8 ;
 RECT 0.54 1.76 0.68 2.8 ;
 RECT 10.18 2.055 10.32 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 13.76 0.08 ;
 RECT 11.185 0.08 11.455 0.245 ;
 RECT 12.2 0.08 12.47 0.245 ;
 RECT 3.42 0.08 3.56 0.505 ;
 RECT 3.995 0.08 4.225 0.385 ;
 RECT 6.385 0.08 6.525 0.38 ;
 RECT 0.54 0.08 0.68 0.83 ;
 RECT 9.695 0.08 9.835 1.07 ;
 RECT 13.215 0.08 13.355 0.825 ;
 RECT 1.51 0.08 1.65 1.075 ;
 END
 END VSS

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.925 0.475 9.285 0.81 ;
 END
 ANTENNAGATEAREA 0.088 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.515 1.495 1.925 1.905 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.9 2.115 2.255 2.385 ;
 RECT 2.815 1.635 2.955 1.74 ;
 RECT 2.115 1.74 2.955 1.91 ;
 RECT 2.115 1.91 2.255 2.115 ;
 RECT 2.115 1.13 2.255 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.485 1.155 2.84 1.435 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.48 1.47 3.885 1.765 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.665 2.08 12.02 2.375 ;
 RECT 11.78 2.375 11.92 2.51 ;
 RECT 11.78 0.665 11.92 2.08 ;
 END
 ANTENNADIFFAREA 0.616 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.635 2.08 12.965 2.375 ;
 RECT 12.745 2.375 12.885 2.51 ;
 RECT 12.745 0.595 12.885 2.08 ;
 END
 ANTENNADIFFAREA 0.622 ;
 END Q

 OBS
 LAYER PO ;
 RECT 7.275 0.865 7.545 1.095 ;
 RECT 7.725 0.265 7.825 0.575 ;
 RECT 7.075 0.575 7.825 0.675 ;
 RECT 7.725 0.675 7.825 1.35 ;
 RECT 8.17 1.545 8.27 2.445 ;
 RECT 9.48 0.265 9.58 1.32 ;
 RECT 7.075 0.455 7.305 0.575 ;
 RECT 7.075 0.675 7.305 0.685 ;
 RECT 7.915 1.45 8.27 1.545 ;
 RECT 7.725 0.165 9.58 0.265 ;
 RECT 7.725 1.35 8.015 1.445 ;
 RECT 7.725 1.445 8.27 1.45 ;
 RECT 4.84 0.285 4.94 0.5 ;
 RECT 4.84 0.185 6.27 0.285 ;
 RECT 6.17 0.285 6.27 1.24 ;
 RECT 4.8 0.5 5.03 0.735 ;
 RECT 5.34 1.77 5.44 2.495 ;
 RECT 4.735 1.77 4.98 1.92 ;
 RECT 4.735 1.67 5.44 1.77 ;
 RECT 2.485 1.43 2.585 1.665 ;
 RECT 2.905 0.675 3.005 1.2 ;
 RECT 2.485 1.2 3.005 1.43 ;
 RECT 2.435 1.665 2.585 1.765 ;
 RECT 2.435 1.765 2.535 2.49 ;
 RECT 1.295 1.495 1.865 1.77 ;
 RECT 1.765 0.675 1.865 1.495 ;
 RECT 1.765 1.77 1.865 2.485 ;
 RECT 1.295 0.655 1.395 1.495 ;
 RECT 1.295 1.77 1.395 2.485 ;
 RECT 3 0.195 3.305 0.425 ;
 RECT 3.205 0.425 3.305 2.485 ;
 RECT 2.765 1.655 3.005 1.885 ;
 RECT 2.905 1.885 3.005 2.5 ;
 RECT 6.795 1.275 7.2 1.375 ;
 RECT 7.1 1.375 7.2 2.69 ;
 RECT 7.1 2.69 9.24 2.79 ;
 RECT 9.14 0.705 9.24 2.69 ;
 RECT 6.795 0.635 6.895 1.275 ;
 RECT 9.01 0.495 9.24 0.705 ;
 RECT 8.665 0.645 8.765 1.24 ;
 RECT 8.665 1.24 8.91 1.45 ;
 RECT 8.665 1.45 8.765 2.37 ;
 RECT 8.195 0.685 8.295 1.23 ;
 RECT 8.12 0.455 8.35 0.685 ;
 RECT 6.495 0.625 6.595 1.58 ;
 RECT 6.625 1.82 6.725 2.39 ;
 RECT 6.495 1.58 6.735 1.82 ;
 RECT 5.835 1.43 5.935 1.475 ;
 RECT 5.835 1.71 5.935 2.505 ;
 RECT 5.855 0.65 5.955 1.33 ;
 RECT 5.835 1.33 5.955 1.43 ;
 RECT 5.705 1.475 5.935 1.71 ;
 RECT 3.68 0.675 3.78 1.5 ;
 RECT 3.485 1.5 3.78 1.74 ;
 RECT 3.68 1.74 3.78 2.39 ;
 RECT 2.1 0.66 2.2 1.165 ;
 RECT 2.06 1.165 2.305 1.405 ;
 RECT 4.205 1.44 4.555 1.69 ;
 RECT 4.455 1.69 4.555 2.685 ;
 RECT 4.455 1.355 4.555 1.44 ;
 RECT 5.385 0.705 5.485 1.255 ;
 RECT 6.14 1.795 6.24 2.685 ;
 RECT 4.455 2.685 6.24 2.785 ;
 RECT 4.455 1.255 5.485 1.355 ;
 RECT 5.385 0.47 5.67 0.705 ;
 RECT 4.52 0.515 4.62 1.255 ;
 RECT 12.415 1.1 12.63 1.18 ;
 RECT 12.415 1.18 13.1 1.28 ;
 RECT 12.415 1.28 12.63 1.335 ;
 RECT 13 0.145 13.1 1.18 ;
 RECT 13 1.28 13.1 2.79 ;
 RECT 12.53 0.145 12.63 1.1 ;
 RECT 12.53 1.335 12.63 2.79 ;
 RECT 10.985 1.18 12.135 1.28 ;
 RECT 10.985 1.28 11.195 1.415 ;
 RECT 11.565 0.145 11.665 1.18 ;
 RECT 11.565 1.28 11.665 2.79 ;
 RECT 12.035 0.145 12.135 1.18 ;
 RECT 12.035 1.28 12.135 2.79 ;
 RECT 9.75 2.47 10.065 2.71 ;
 RECT 9.965 1.88 10.065 2.47 ;
 RECT 9.95 1.53 10.535 1.63 ;
 RECT 10.31 1.63 10.535 1.94 ;
 RECT 9.95 0.65 10.05 1.53 ;
 RECT 10.435 1.94 10.535 2.565 ;
 RECT 7.38 1.64 7.76 1.87 ;
 RECT 7.38 1.095 7.545 1.64 ;
 LAYER CO ;
 RECT 5.755 1.525 5.885 1.655 ;
 RECT 6.85 2.015 6.98 2.145 ;
 RECT 4.045 0.25 4.175 0.38 ;
 RECT 12.255 1.79 12.385 1.92 ;
 RECT 12.255 2.05 12.385 2.18 ;
 RECT 12.255 2.31 12.385 2.44 ;
 RECT 11.255 0.11 11.385 0.24 ;
 RECT 12.455 1.15 12.585 1.28 ;
 RECT 13.22 0.625 13.35 0.755 ;
 RECT 11.785 1.79 11.915 1.92 ;
 RECT 11.785 1.53 11.915 1.66 ;
 RECT 11.785 2.05 11.915 2.18 ;
 RECT 9.7 0.87 9.83 1 ;
 RECT 11.025 1.23 11.155 1.36 ;
 RECT 11.31 1.53 11.44 1.66 ;
 RECT 3.425 0.26 3.555 0.39 ;
 RECT 3.05 0.245 3.18 0.375 ;
 RECT 4.85 0.555 4.98 0.685 ;
 RECT 2.655 2.135 2.785 2.265 ;
 RECT 2.64 1.25 2.77 1.38 ;
 RECT 0.545 2.365 0.675 2.495 ;
 RECT 3.9 2.015 4.03 2.145 ;
 RECT 1.515 0.895 1.645 1.025 ;
 RECT 0.545 2.105 0.675 2.235 ;
 RECT 4.03 0.895 4.16 1.025 ;
 RECT 0.545 1.845 0.675 1.975 ;
 RECT 1.515 2.135 1.645 2.265 ;
 RECT 1.52 1.57 1.65 1.7 ;
 RECT 3.425 2.07 3.555 2.2 ;
 RECT 4.275 1.495 4.405 1.625 ;
 RECT 4.145 2.365 4.275 2.495 ;
 RECT 5.585 2.07 5.715 2.2 ;
 RECT 5.605 0.88 5.735 1.01 ;
 RECT 5.09 2.105 5.22 2.235 ;
 RECT 5.135 0.88 5.265 1.01 ;
 RECT 4.74 0.905 4.87 1.035 ;
 RECT 4.675 2.23 4.805 2.36 ;
 RECT 5.49 0.525 5.62 0.655 ;
 RECT 7.015 0.88 7.145 1.01 ;
 RECT 6.39 0.2 6.52 0.33 ;
 RECT 9.815 2.525 9.945 2.655 ;
 RECT 7.92 1.815 8.05 1.945 ;
 RECT 7.41 2.44 7.54 2.57 ;
 RECT 7.58 1.69 7.71 1.82 ;
 RECT 7.34 0.915 7.47 1.045 ;
 RECT 8.415 0.87 8.545 1 ;
 RECT 9.365 1.965 9.495 2.095 ;
 RECT 8.885 1.965 9.015 2.095 ;
 RECT 6.465 2.64 6.595 2.77 ;
 RECT 8.725 1.28 8.855 1.41 ;
 RECT 10.17 0.87 10.3 1 ;
 RECT 10.185 2.115 10.315 2.245 ;
 RECT 9.715 2.11 9.845 2.24 ;
 RECT 13.225 1.53 13.355 1.66 ;
 RECT 13.225 1.79 13.355 1.92 ;
 RECT 13.225 2.05 13.355 2.18 ;
 RECT 13.225 2.31 13.355 2.44 ;
 RECT 12.75 1.79 12.88 1.92 ;
 RECT 12.75 1.53 12.88 1.66 ;
 RECT 12.75 2.05 12.88 2.18 ;
 RECT 12.75 0.645 12.88 0.775 ;
 RECT 12.75 2.31 12.88 2.44 ;
 RECT 12.28 0.11 12.41 0.24 ;
 RECT 12.255 1.53 12.385 1.66 ;
 RECT 11.31 1.79 11.44 1.92 ;
 RECT 11.31 2.05 11.44 2.18 ;
 RECT 11.31 2.31 11.44 2.44 ;
 RECT 11.785 0.715 11.915 0.845 ;
 RECT 11.785 2.31 11.915 2.44 ;
 RECT 4.805 1.725 4.935 1.855 ;
 RECT 1.045 2.075 1.175 2.205 ;
 RECT 0.545 0.63 0.675 0.76 ;
 RECT 2.12 1.215 2.25 1.345 ;
 RECT 0.545 0.37 0.675 0.5 ;
 RECT 1.045 0.895 1.175 1.025 ;
 RECT 3.535 1.555 3.665 1.685 ;
 RECT 2.46 0.545 2.59 0.675 ;
 RECT 2.82 1.705 2.95 1.835 ;
 RECT 9.06 0.535 9.19 0.665 ;
 RECT 7.125 0.505 7.255 0.635 ;
 RECT 8.415 1.9 8.545 2.03 ;
 RECT 7.945 0.87 8.075 1 ;
 RECT 8.17 0.505 8.3 0.635 ;
 RECT 10.745 2.13 10.875 2.26 ;
 RECT 10.36 1.76 10.49 1.89 ;
 RECT 6.565 1.63 6.695 1.76 ;
 LAYER M1 ;
 RECT 7.125 1.36 7.265 2.1 ;
 RECT 7.125 2.24 7.265 2.355 ;
 RECT 6.05 2.355 7.265 2.495 ;
 RECT 4.67 2.515 6.19 2.655 ;
 RECT 4.735 0.735 4.875 1.72 ;
 RECT 4.735 1.72 4.985 1.775 ;
 RECT 4.67 1.775 4.985 1.86 ;
 RECT 4.67 1.86 4.875 2.005 ;
 RECT 4.67 2.005 4.81 2.515 ;
 RECT 4.845 0.505 4.985 0.535 ;
 RECT 6.05 2.495 6.19 2.515 ;
 RECT 4.735 0.535 4.985 0.735 ;
 RECT 8.53 2.32 8.67 2.52 ;
 RECT 7.66 0.5 8.375 0.64 ;
 RECT 7.66 0.64 7.8 1.22 ;
 RECT 7.125 2.1 8.025 2.18 ;
 RECT 7.125 2.18 8.67 2.24 ;
 RECT 7.885 2.24 8.67 2.32 ;
 RECT 7.125 1.22 7.8 1.36 ;
 RECT 8.53 2.52 10.025 2.66 ;
 RECT 4.025 0.845 4.165 1.125 ;
 RECT 4.025 1.125 4.41 1.265 ;
 RECT 4.27 1.265 4.41 2.01 ;
 RECT 3.83 2.01 4.41 2.15 ;
 RECT 6.845 1.04 7.52 1.05 ;
 RECT 6.28 0.91 7.52 1.04 ;
 RECT 6.28 0.9 7.15 0.91 ;
 RECT 6.845 1.08 6.985 2.2 ;
 RECT 6.845 1.05 7.15 1.08 ;
 RECT 5.705 1.52 6.42 1.66 ;
 RECT 7.01 0.81 7.15 0.9 ;
 RECT 6.28 1.04 6.42 1.52 ;
 RECT 1.04 0.82 1.18 1.215 ;
 RECT 1.04 1.355 1.18 2.325 ;
 RECT 1.825 0.38 1.965 1.215 ;
 RECT 1.04 1.215 1.965 1.355 ;
 RECT 1.825 0.24 3.25 0.38 ;
 RECT 5.42 0.52 7.33 0.66 ;
 RECT 7.045 0.47 7.33 0.52 ;
 RECT 8.41 0.805 8.55 1.675 ;
 RECT 8.41 1.815 8.62 1.895 ;
 RECT 8.34 1.895 8.62 2.035 ;
 RECT 9.315 1.815 9.545 2.1 ;
 RECT 8.41 1.675 10.6 1.815 ;
 RECT 11.02 1.18 11.16 2.505 ;
 RECT 10.3 1.815 10.6 1.915 ;
 RECT 10.46 1.915 10.6 2.505 ;
 RECT 10.46 2.505 11.16 2.645 ;
 RECT 8.88 2.1 9.065 2.24 ;
 RECT 9.71 2.03 9.85 2.24 ;
 RECT 8.835 1.96 9.065 2.1 ;
 RECT 8.88 2.24 9.85 2.38 ;
 RECT 7.57 1.685 8.08 1.81 ;
 RECT 7.94 0.78 8.08 1.685 ;
 RECT 7.57 1.615 7.71 1.685 ;
 RECT 7.57 1.825 7.71 1.895 ;
 RECT 7.57 1.81 8.12 1.825 ;
 RECT 7.85 1.825 8.12 1.95 ;
 RECT 5.425 1.805 6.7 1.945 ;
 RECT 5.425 1.945 5.79 1.96 ;
 RECT 5.425 1.22 5.74 1.36 ;
 RECT 5.6 0.805 5.74 1.22 ;
 RECT 5.51 1.96 5.79 2.215 ;
 RECT 5.425 1.36 5.565 1.805 ;
 RECT 6.56 1.56 6.7 1.805 ;
 RECT 10.74 0.745 11.63 0.865 ;
 RECT 10.12 0.865 11.63 0.885 ;
 RECT 11.49 0.525 11.63 0.745 ;
 RECT 10.12 0.885 10.88 1.005 ;
 RECT 10.74 1.005 10.88 1.395 ;
 RECT 10.74 1.535 10.88 2.32 ;
 RECT 8.72 1.395 10.88 1.535 ;
 RECT 8.72 1.21 8.86 1.395 ;
 RECT 11.49 0.385 12.59 0.525 ;
 RECT 12.45 0.525 12.59 1.34 ;
 RECT 3.095 1.025 3.235 2.13 ;
 RECT 3.095 0.68 3.235 0.885 ;
 RECT 2.585 2.13 3.235 2.27 ;
 RECT 2.395 0.54 3.235 0.68 ;
 RECT 3.7 0.665 3.84 0.885 ;
 RECT 3.095 0.885 3.84 1.025 ;
 RECT 5.13 0.36 5.27 0.875 ;
 RECT 5.145 1.015 5.285 2.035 ;
 RECT 3.7 0.525 4.59 0.665 ;
 RECT 4.45 0.36 4.59 0.525 ;
 RECT 5.085 2.035 5.285 2.305 ;
 RECT 5.085 0.875 5.34 1.015 ;
 RECT 4.45 0.22 5.27 0.36 ;
 END
END SDFFASX2

MACRO SDFFNARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 13.12 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 13.12 2.96 ;
 RECT 3.835 2.635 4.085 2.8 ;
 RECT 1.27 2.005 1.41 2.8 ;
 RECT 7.265 2.635 7.525 2.8 ;
 RECT 3.18 1.98 3.32 2.8 ;
 RECT 9.915 1.955 10.055 2.8 ;
 RECT 11.095 2.06 11.235 2.8 ;
 RECT 12.62 1.73 12.76 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 13.12 0.08 ;
 RECT 9.92 0.08 10.175 0.285 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 3.81 0.08 4.11 0.26 ;
 RECT 6.525 0.08 6.76 0.26 ;
 RECT 12.705 0.08 12.845 0.88 ;
 RECT 11.115 0.08 11.255 0.64 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 1.055 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.515 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.335 0.28 10.615 0.42 ;
 RECT 5.92 0.51 7.04 0.65 ;
 RECT 9.285 0.36 9.71 0.505 ;
 RECT 9.285 0.505 10.555 0.645 ;
 RECT 6.9 0.36 7.04 0.51 ;
 RECT 10.415 0.225 10.555 0.28 ;
 RECT 6.9 0.22 9.71 0.36 ;
 RECT 10.335 0.42 10.555 0.505 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.84 1.75 2.24 1.855 ;
 RECT 1.84 1.48 2.24 1.61 ;
 RECT 2.575 1.75 2.715 1.78 ;
 RECT 1.84 1.61 2.715 1.75 ;
 RECT 2.575 1.505 2.715 1.61 ;
 RECT 1.875 1.11 2.015 1.48 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.205 2.275 2.56 2.66 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.655 1.105 12.005 1.425 ;
 RECT 11.68 1.425 11.82 2.35 ;
 RECT 11.68 0.55 11.82 1.105 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.09 2.015 12.465 2.38 ;
 RECT 12.145 0.7 12.285 2.015 ;
 END
 ANTENNADIFFAREA 0.456 ;
 END Q

 OBS
 LAYER PO ;
 RECT 5.595 1.475 5.825 1.71 ;
 RECT 11.43 0.16 11.53 1.17 ;
 RECT 11.43 1.4 11.53 2.62 ;
 RECT 11.18 1.17 11.53 1.4 ;
 RECT 2.665 1.755 2.765 2.48 ;
 RECT 2.525 1.525 2.765 1.755 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 7.86 0.875 8.255 1.105 ;
 RECT 8.155 1.105 8.255 1.64 ;
 RECT 8.155 1.64 8.39 1.87 ;
 RECT 10.79 1.32 10.89 2.545 ;
 RECT 10.49 0.47 10.59 1.22 ;
 RECT 10.49 1.22 10.89 1.32 ;
 RECT 10.36 0.23 10.59 0.47 ;
 RECT 6.035 0.695 6.135 1.61 ;
 RECT 6.07 1.71 6.17 2.48 ;
 RECT 6.035 1.61 6.17 1.71 ;
 RECT 5.915 0.465 6.155 0.695 ;
 RECT 8.44 0.265 8.54 0.575 ;
 RECT 8.44 0.675 8.54 1.35 ;
 RECT 7.635 0.575 8.54 0.675 ;
 RECT 8.885 1.545 8.985 2.405 ;
 RECT 9.775 0.265 9.875 1.32 ;
 RECT 7.635 0.46 7.865 0.575 ;
 RECT 7.635 0.675 7.865 0.69 ;
 RECT 8.63 1.45 8.985 1.545 ;
 RECT 8.44 0.165 9.875 0.265 ;
 RECT 8.44 1.35 8.73 1.445 ;
 RECT 8.44 1.445 8.985 1.45 ;
 RECT 9.38 0.645 9.48 1.24 ;
 RECT 9.38 1.45 9.48 2.37 ;
 RECT 9.36 1.24 9.595 1.45 ;
 RECT 8.91 0.685 9.01 1.255 ;
 RECT 8.835 0.455 9.065 0.685 ;
 RECT 10.19 0.65 10.29 1.71 ;
 RECT 10.19 1.71 10.435 1.95 ;
 RECT 10.19 1.95 10.29 2.56 ;
 RECT 7.2 1.61 7.465 1.82 ;
 RECT 7.365 1.82 7.465 2.52 ;
 RECT 6.995 0.635 7.095 1.51 ;
 RECT 6.995 1.51 7.465 1.61 ;
 RECT 12.405 0.355 12.505 1.05 ;
 RECT 12.405 1.285 12.505 2.79 ;
 RECT 12.39 1.05 12.6 1.285 ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 5.145 0.705 5.245 1.21 ;
 RECT 5.145 0.47 5.43 0.705 ;
 RECT 4.575 1.16 4.82 1.21 ;
 RECT 4.575 1.31 4.82 1.405 ;
 RECT 4.575 1.21 5.245 1.31 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.245 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 2.665 0.655 2.765 1.245 ;
 RECT 2.245 1.345 2.345 1.645 ;
 RECT 2.195 1.745 2.295 2.44 ;
 RECT 2.195 2.44 2.445 2.67 ;
 RECT 2.245 1.245 2.765 1.345 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 9.7 1.64 9.8 2.585 ;
 RECT 8.48 2.47 8.7 2.585 ;
 RECT 8.48 2.585 9.8 2.685 ;
 RECT 8.48 2.685 8.7 2.71 ;
 RECT 5.1 1.685 5.2 2.495 ;
 RECT 3.78 1.52 4.38 1.585 ;
 RECT 3.78 1.585 5.2 1.62 ;
 RECT 3.78 1.62 4.025 1.69 ;
 RECT 4.215 1.62 5.2 1.685 ;
 RECT 4.215 1.685 4.315 2.27 ;
 RECT 3.78 1.44 4.025 1.52 ;
 RECT 4.28 0.685 4.38 1.52 ;
 RECT 4.6 0.285 4.7 0.585 ;
 RECT 4.6 0.185 6.435 0.285 ;
 RECT 6.335 0.285 6.435 1.24 ;
 RECT 4.28 0.585 4.7 0.685 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 6.895 1.79 6.995 2.685 ;
 RECT 4.62 2.33 4.72 2.685 ;
 RECT 4.62 2.685 6.995 2.785 ;
 RECT 4.5 2.09 4.72 2.33 ;
 RECT 5.595 1.33 5.735 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.635 0.65 5.735 1.33 ;
 LAYER CO ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 8.53 2.525 8.66 2.655 ;
 RECT 9.13 0.87 9.26 1 ;
 RECT 12.15 1.91 12.28 2.04 ;
 RECT 9.92 2.01 10.05 2.14 ;
 RECT 11.1 2.13 11.23 2.26 ;
 RECT 10.54 2.13 10.67 2.26 ;
 RECT 7.255 1.63 7.385 1.76 ;
 RECT 5.645 1.525 5.775 1.655 ;
 RECT 7.59 0.88 7.72 1.01 ;
 RECT 7.585 2.015 7.715 2.145 ;
 RECT 3.93 0.125 4.06 0.255 ;
 RECT 7.315 2.64 7.445 2.77 ;
 RECT 6.645 2.125 6.775 2.255 ;
 RECT 6.295 1.82 6.425 1.95 ;
 RECT 5.815 2.105 5.945 2.235 ;
 RECT 3.905 2.64 4.035 2.77 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 4.63 1.205 4.76 1.335 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 3.295 1.535 3.425 1.665 ;
 RECT 3.71 1.995 3.84 2.125 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2 2.545 2.13 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 7.675 0.51 7.805 0.64 ;
 RECT 10.26 1.765 10.39 1.895 ;
 RECT 8.635 1.815 8.765 1.945 ;
 RECT 4.55 2.145 4.68 2.275 ;
 RECT 9.13 1.9 9.26 2.03 ;
 RECT 12.43 1.1 12.56 1.23 ;
 RECT 4.435 1.825 4.565 1.955 ;
 RECT 12.71 0.68 12.84 0.81 ;
 RECT 12.15 1.65 12.28 1.78 ;
 RECT 5.25 0.525 5.38 0.655 ;
 RECT 12.15 2.17 12.28 2.3 ;
 RECT 12.15 0.75 12.28 0.88 ;
 RECT 11.23 1.22 11.36 1.35 ;
 RECT 12.625 1.8 12.755 1.93 ;
 RECT 12.625 2.06 12.755 2.19 ;
 RECT 11.685 0.615 11.815 0.745 ;
 RECT 11.685 1.87 11.815 2 ;
 RECT 11.685 2.13 11.815 2.26 ;
 RECT 11.12 0.435 11.25 0.565 ;
 RECT 2.58 1.575 2.71 1.705 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 8.21 1.69 8.34 1.82 ;
 RECT 7.93 0.915 8.06 1.045 ;
 RECT 10.41 0.285 10.54 0.415 ;
 RECT 9.995 0.15 10.125 0.28 ;
 RECT 5.97 0.515 6.1 0.645 ;
 RECT 6.575 0.12 6.705 0.25 ;
 RECT 8.66 0.87 8.79 1 ;
 RECT 8.885 0.505 9.015 0.635 ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 9.41 1.28 9.54 1.41 ;
 RECT 10.71 0.87 10.84 1 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 2.265 2.49 2.395 2.62 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 LAYER M1 ;
 RECT 9.405 1.21 9.545 1.395 ;
 RECT 9.405 1.395 10.675 1.535 ;
 RECT 10.535 1.105 10.675 1.395 ;
 RECT 10.535 1.535 10.675 2.33 ;
 RECT 10.705 0.92 10.845 0.965 ;
 RECT 10.535 0.965 10.845 1.105 ;
 RECT 10.705 0.78 11.535 0.92 ;
 RECT 11.395 0.36 11.535 0.78 ;
 RECT 11.395 0.22 12.39 0.36 ;
 RECT 12.425 0.56 12.565 1.41 ;
 RECT 12.25 0.36 12.39 0.42 ;
 RECT 12.25 0.42 12.565 0.56 ;
 RECT 5.18 0.52 5.78 0.66 ;
 RECT 5.64 0.66 5.78 0.79 ;
 RECT 7.18 0.505 7.855 0.645 ;
 RECT 5.64 0.79 7.32 0.93 ;
 RECT 7.18 0.645 7.32 0.79 ;
 RECT 7.58 1.015 8.13 1.05 ;
 RECT 7.58 1.05 7.72 1.185 ;
 RECT 7.52 0.91 8.13 1.015 ;
 RECT 7.52 0.875 7.79 0.91 ;
 RECT 6.97 1.185 7.72 1.325 ;
 RECT 7.58 1.325 7.72 2.215 ;
 RECT 6.97 1.325 7.11 1.52 ;
 RECT 5.575 1.52 7.11 1.66 ;
 RECT 5.745 2.12 6.845 2.24 ;
 RECT 5.745 2.1 6.015 2.12 ;
 RECT 5.81 2.24 6.845 2.26 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 10.815 1.92 10.955 2.505 ;
 RECT 9.125 1.675 10.395 1.815 ;
 RECT 10.255 2.505 10.955 2.645 ;
 RECT 10.255 1.815 10.395 2.505 ;
 RECT 9.125 1.815 9.335 1.895 ;
 RECT 9.125 0.805 9.265 1.675 ;
 RECT 9.055 1.895 9.335 2.035 ;
 RECT 11.05 1.355 11.19 1.78 ;
 RECT 11.05 1.215 11.43 1.355 ;
 RECT 10.815 1.78 11.19 1.92 ;
 RECT 4.495 1.385 4.635 1.82 ;
 RECT 4.365 1.825 4.685 1.96 ;
 RECT 4.365 1.82 4.635 1.825 ;
 RECT 4.545 1.96 4.685 2.345 ;
 RECT 4.495 0.84 4.635 1.155 ;
 RECT 4.495 1.155 4.765 1.385 ;
 RECT 4.225 2.65 6.33 2.655 ;
 RECT 4.225 2.49 4.365 2.515 ;
 RECT 3.705 1.63 3.845 2.35 ;
 RECT 3.705 1.475 4.045 1.63 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.705 2.35 4.365 2.49 ;
 RECT 4.225 2.515 7.125 2.65 ;
 RECT 6.19 2.51 7.125 2.515 ;
 RECT 6.985 2.495 7.125 2.51 ;
 RECT 8.3 0.58 9.09 0.64 ;
 RECT 8.3 0.64 8.76 0.72 ;
 RECT 8.58 0.5 9.09 0.58 ;
 RECT 7.86 1.21 8.44 1.35 ;
 RECT 7.86 1.35 8 2.1 ;
 RECT 7.86 2.1 8.6 2.24 ;
 RECT 7.86 2.24 8 2.355 ;
 RECT 8.46 2.24 8.6 2.52 ;
 RECT 6.985 2.355 8 2.495 ;
 RECT 8.46 2.52 8.73 2.66 ;
 RECT 8.3 0.72 8.44 1.21 ;
 RECT 8.14 1.685 8.795 1.81 ;
 RECT 8.655 1.005 8.795 1.685 ;
 RECT 8.14 1.81 8.835 1.825 ;
 RECT 8.565 1.825 8.835 1.95 ;
 RECT 8.585 0.865 8.865 1.005 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 1.995 ;
 RECT 2.855 2.135 2.995 2.195 ;
 RECT 2.365 1.995 2.995 2.135 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 3.46 0.53 4.41 0.67 ;
 RECT 4.27 0.22 5.03 0.36 ;
 RECT 4.89 0.36 5.03 0.875 ;
 RECT 4.905 1.015 5.045 2.035 ;
 RECT 4.845 2.035 5.045 2.17 ;
 RECT 4.845 2.17 4.985 2.305 ;
 RECT 4.27 0.36 4.41 0.53 ;
 RECT 4.825 0.875 5.1 1.015 ;
 RECT 5.185 1.82 7.39 1.945 ;
 RECT 5.185 1.945 6.495 1.96 ;
 RECT 6.21 1.805 7.39 1.82 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 5.36 0.805 5.5 1.22 ;
 RECT 7.25 1.56 7.39 1.805 ;
 RECT 5.185 1.36 5.325 1.82 ;
 END
END SDFFNARX1

MACRO DFFNX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.88 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.88 2.96 ;
 RECT 4.405 2.635 4.665 2.8 ;
 RECT 2.045 2.625 2.295 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 8.595 1.54 8.735 2.8 ;
 RECT 9.615 1.54 9.755 2.8 ;
 RECT 10.555 1.54 10.695 2.8 ;
 RECT 1.39 1.98 1.53 2.8 ;
 RECT 7.315 1.955 7.455 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.88 0.08 ;
 RECT 1.39 0.08 1.53 1.055 ;
 RECT 2.02 0.08 2.32 0.39 ;
 RECT 7.32 0.08 7.575 0.535 ;
 RECT 9.545 0.08 9.8 0.3 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.34 0.08 4.48 0.58 ;
 RECT 8.58 0.08 8.72 0.6 ;
 RECT 10.555 0.08 10.695 0.685 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.495 1.475 2.025 1.735 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.95 2.12 9.28 2.39 ;
 RECT 9.14 2.39 9.28 2.575 ;
 RECT 9.14 0.72 9.28 2.12 ;
 END
 ANTENNADIFFAREA 0.748 ;
 END QN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.95 1.475 1.32 1.785 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.895 2.1 10.225 2.35 ;
 RECT 10.085 2.35 10.225 2.575 ;
 RECT 10.085 0.72 10.225 2.1 ;
 END
 ANTENNADIFFAREA 0.622 ;
 END Q

 OBS
 LAYER PO ;
 RECT 3.825 0.65 3.925 1.33 ;
 RECT 5.84 0.525 5.94 1.35 ;
 RECT 7.175 0.265 7.275 1.32 ;
 RECT 5.84 0.265 5.94 0.295 ;
 RECT 5.035 0.295 5.94 0.525 ;
 RECT 6.285 1.51 6.385 2.48 ;
 RECT 5.84 0.165 7.275 0.265 ;
 RECT 5.84 1.35 6.13 1.41 ;
 RECT 5.84 1.41 6.385 1.45 ;
 RECT 6.03 1.45 6.385 1.51 ;
 RECT 2.28 1.49 2.59 1.56 ;
 RECT 2.49 0.285 2.59 1.49 ;
 RECT 2.49 0.185 4.225 0.285 ;
 RECT 2.425 1.735 2.525 2.21 ;
 RECT 3.31 1.66 3.41 2.49 ;
 RECT 2.28 1.56 3.41 1.66 ;
 RECT 2.28 1.66 2.525 1.735 ;
 RECT 3.31 1.53 3.41 1.56 ;
 RECT 4.125 0.285 4.225 1.26 ;
 RECT 10.34 0.2 10.44 1.225 ;
 RECT 9.87 1.325 9.97 2.79 ;
 RECT 10.34 1.325 10.44 2.79 ;
 RECT 9.76 1.225 10.44 1.27 ;
 RECT 9.76 1.035 9.97 1.225 ;
 RECT 9.87 1.27 10.44 1.325 ;
 RECT 9.87 0.2 9.97 1.035 ;
 RECT 8.115 1.12 8.95 1.225 ;
 RECT 8.115 1.225 9.495 1.325 ;
 RECT 8.85 0.195 8.95 1.12 ;
 RECT 8.85 1.35 8.95 2.79 ;
 RECT 8.115 1.325 8.95 1.35 ;
 RECT 9.395 0.2 9.495 1.225 ;
 RECT 9.395 1.325 9.495 2.79 ;
 RECT 3.355 0.705 3.455 1.155 ;
 RECT 3.355 0.47 3.645 0.705 ;
 RECT 2.77 1.255 3.015 1.38 ;
 RECT 2.77 1.155 3.455 1.255 ;
 RECT 7.1 1.64 7.2 2.69 ;
 RECT 5.88 2.47 6.1 2.69 ;
 RECT 5.88 2.69 7.2 2.79 ;
 RECT 1.65 0.655 1.75 1.48 ;
 RECT 1.455 1.48 1.75 1.72 ;
 RECT 1.65 1.72 1.75 2.37 ;
 RECT 7.59 0.65 7.69 1.48 ;
 RECT 7.59 1.72 7.69 2.56 ;
 RECT 7.495 1.48 7.725 1.72 ;
 RECT 4.565 0.635 4.665 1.415 ;
 RECT 4.565 1.415 4.885 1.645 ;
 RECT 4.565 1.645 4.665 2.49 ;
 RECT 4.125 1.53 4.225 2.685 ;
 RECT 2.71 2.075 2.92 2.685 ;
 RECT 2.71 2.685 4.225 2.785 ;
 RECT 1.175 0.655 1.275 1.515 ;
 RECT 1.175 1.745 1.275 2.735 ;
 RECT 1.055 1.515 1.275 1.745 ;
 RECT 5.49 1.105 5.59 1.64 ;
 RECT 5.26 0.875 5.59 1.105 ;
 RECT 5.49 1.64 5.725 1.87 ;
 RECT 6.78 0.645 6.88 1.24 ;
 RECT 6.78 1.45 6.88 2.505 ;
 RECT 6.76 1.24 6.995 1.45 ;
 RECT 6.31 0.685 6.41 1.22 ;
 RECT 6.235 0.455 6.465 0.685 ;
 RECT 3.805 1.64 3.925 1.71 ;
 RECT 3.805 1.71 3.905 2.49 ;
 RECT 3.805 1.33 3.925 1.405 ;
 RECT 3.69 1.405 3.925 1.64 ;
 LAYER CO ;
 RECT 1.505 1.535 1.635 1.665 ;
 RECT 1.92 1.995 2.05 2.125 ;
 RECT 2 0.875 2.13 1.005 ;
 RECT 1.395 2.05 1.525 2.18 ;
 RECT 1.395 0.875 1.525 1.005 ;
 RECT 7.81 0.87 7.94 1 ;
 RECT 7.32 2.01 7.45 2.14 ;
 RECT 4.7 1.455 4.83 1.585 ;
 RECT 10.56 1.85 10.69 1.98 ;
 RECT 10.56 2.115 10.69 2.245 ;
 RECT 10.56 2.375 10.69 2.505 ;
 RECT 10.09 1.85 10.22 1.98 ;
 RECT 10.09 2.115 10.22 2.245 ;
 RECT 10.09 2.375 10.22 2.505 ;
 RECT 10.09 1.59 10.22 1.72 ;
 RECT 10.09 0.77 10.22 0.9 ;
 RECT 9.62 0.165 9.75 0.295 ;
 RECT 9.62 1.59 9.75 1.72 ;
 RECT 9.62 1.85 9.75 1.98 ;
 RECT 9.145 2.375 9.275 2.505 ;
 RECT 9.145 0.77 9.275 0.9 ;
 RECT 5.33 0.915 5.46 1.045 ;
 RECT 7.395 0.4 7.525 0.53 ;
 RECT 0.925 0.875 1.055 1.005 ;
 RECT 0.925 2.05 1.055 2.18 ;
 RECT 8.6 1.85 8.73 1.98 ;
 RECT 8.6 2.115 8.73 2.245 ;
 RECT 8.6 2.375 8.73 2.505 ;
 RECT 9.145 1.59 9.275 1.72 ;
 RECT 9.145 1.85 9.275 1.98 ;
 RECT 2.645 1.825 2.775 1.955 ;
 RECT 2.75 2.13 2.88 2.26 ;
 RECT 1.105 1.565 1.235 1.695 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 5.93 2.525 6.06 2.655 ;
 RECT 6.035 1.815 6.165 1.945 ;
 RECT 9.8 1.085 9.93 1.215 ;
 RECT 8.165 1.17 8.295 1.3 ;
 RECT 9.145 2.115 9.275 2.245 ;
 RECT 2.115 2.63 2.245 2.76 ;
 RECT 5.545 1.69 5.675 1.82 ;
 RECT 3.06 2.105 3.19 2.235 ;
 RECT 3.105 0.88 3.235 1.01 ;
 RECT 4.345 0.38 4.475 0.51 ;
 RECT 6.53 1.9 6.66 2.03 ;
 RECT 6.53 0.87 6.66 1 ;
 RECT 6.06 0.87 6.19 1 ;
 RECT 6.285 0.505 6.415 0.635 ;
 RECT 6.81 1.28 6.94 1.41 ;
 RECT 2.335 1.535 2.465 1.665 ;
 RECT 3.465 0.525 3.595 0.655 ;
 RECT 7.88 2.13 8.01 2.26 ;
 RECT 5.075 0.345 5.205 0.475 ;
 RECT 7.55 1.535 7.68 1.665 ;
 RECT 3.74 1.46 3.87 1.59 ;
 RECT 4.99 0.88 5.12 1.01 ;
 RECT 4.985 2.015 5.115 2.145 ;
 RECT 2.14 0.235 2.27 0.365 ;
 RECT 4.455 2.64 4.585 2.77 ;
 RECT 9.62 2.115 9.75 2.245 ;
 RECT 9.62 2.375 9.75 2.505 ;
 RECT 8.585 0.42 8.715 0.55 ;
 RECT 8.6 1.59 8.73 1.72 ;
 RECT 3.555 2.07 3.685 2.2 ;
 RECT 3.575 0.88 3.705 1.01 ;
 RECT 2.825 1.2 2.955 1.33 ;
 RECT 2.715 0.885 2.845 1.015 ;
 RECT 1.395 2.31 1.525 2.44 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 10.56 0.505 10.69 0.635 ;
 RECT 10.56 1.59 10.69 1.72 ;
 RECT 0.305 1.825 0.435 1.955 ;
 LAYER M1 ;
 RECT 4.98 0.875 5.53 1.005 ;
 RECT 3.69 1.455 4.335 1.595 ;
 RECT 4.195 1.005 5.53 1.05 ;
 RECT 4.98 0.805 5.12 0.875 ;
 RECT 4.98 1.145 5.12 2.215 ;
 RECT 4.195 1.05 5.12 1.145 ;
 RECT 4.16 1.595 4.335 1.66 ;
 RECT 4.195 1.145 4.335 1.455 ;
 RECT 3.39 0.52 4.2 0.66 ;
 RECT 4.06 0.66 4.2 0.725 ;
 RECT 4.62 0.34 5.275 0.48 ;
 RECT 4.06 0.725 4.76 0.865 ;
 RECT 4.62 0.48 4.76 0.725 ;
 RECT 2.745 1.965 2.895 2.33 ;
 RECT 2.71 1.41 2.9 1.82 ;
 RECT 2.71 1.96 2.9 1.965 ;
 RECT 2.575 1.82 2.9 1.96 ;
 RECT 2.71 0.81 2.85 1.15 ;
 RECT 2.71 1.15 2.96 1.41 ;
 RECT 0.67 1.01 0.81 1.195 ;
 RECT 0.67 1.335 0.81 2.045 ;
 RECT 0.67 0.87 1.125 1.01 ;
 RECT 0.67 2.045 1.125 2.185 ;
 RECT 1.67 0.67 1.81 1.195 ;
 RECT 0.67 1.195 1.81 1.335 ;
 RECT 1.67 0.53 3.25 0.67 ;
 RECT 3.1 0.67 3.25 1.07 ;
 RECT 3.11 1.07 3.25 2.035 ;
 RECT 3.05 2.035 3.25 2.305 ;
 RECT 6.525 1.815 6.735 1.895 ;
 RECT 6.525 0.805 6.665 1.675 ;
 RECT 6.455 1.895 6.735 2.035 ;
 RECT 6.525 1.675 7.385 1.815 ;
 RECT 7.245 1.67 7.385 1.675 ;
 RECT 8.16 1.12 8.3 2.505 ;
 RECT 7.245 1.53 7.735 1.67 ;
 RECT 7.595 2.505 8.3 2.645 ;
 RECT 7.595 1.67 7.735 2.505 ;
 RECT 5.54 1.685 6.195 1.81 ;
 RECT 6.055 1.005 6.195 1.685 ;
 RECT 5.54 1.81 6.235 1.825 ;
 RECT 5.54 1.825 5.68 1.89 ;
 RECT 5.54 1.62 5.68 1.685 ;
 RECT 5.965 1.825 6.235 1.95 ;
 RECT 5.985 0.865 6.265 1.005 ;
 RECT 8.86 0.58 9 0.84 ;
 RECT 7.805 0.84 9 0.98 ;
 RECT 6.805 1.245 8.015 1.385 ;
 RECT 7.875 1.105 8.015 1.245 ;
 RECT 7.875 1.385 8.015 2.33 ;
 RECT 7.805 0.76 7.945 0.84 ;
 RECT 7.805 0.98 8.015 1.105 ;
 RECT 6.805 1.21 6.945 1.245 ;
 RECT 6.805 1.385 6.945 1.465 ;
 RECT 9.795 0.58 9.935 1.29 ;
 RECT 8.86 0.44 9.935 0.58 ;
 RECT 1.995 1.045 2.305 1.185 ;
 RECT 2.165 1.185 2.305 1.53 ;
 RECT 1.995 0.81 2.135 1.045 ;
 RECT 2.295 1.67 2.435 1.99 ;
 RECT 2.295 2.13 2.435 2.345 ;
 RECT 2.465 2.51 3.97 2.65 ;
 RECT 2.165 1.53 2.57 1.67 ;
 RECT 1.85 1.99 2.435 2.13 ;
 RECT 2.295 2.345 2.605 2.485 ;
 RECT 2.465 2.485 2.605 2.51 ;
 RECT 3.83 2.495 3.97 2.51 ;
 RECT 3.83 2.355 5.4 2.495 ;
 RECT 5.86 2.24 6 2.52 ;
 RECT 5.26 2.24 5.4 2.355 ;
 RECT 5.26 1.35 5.4 2.1 ;
 RECT 5.26 2.1 6 2.24 ;
 RECT 5.26 1.21 5.84 1.35 ;
 RECT 5.86 2.52 6.13 2.66 ;
 RECT 5.98 0.5 6.49 0.58 ;
 RECT 5.7 0.58 6.49 0.64 ;
 RECT 5.7 0.64 6.16 0.72 ;
 RECT 5.7 0.72 5.84 1.21 ;
 RECT 3.395 1.82 4.835 1.915 ;
 RECT 3.48 1.96 3.76 2.215 ;
 RECT 3.48 1.915 4.835 1.96 ;
 RECT 3.395 1.775 3.69 1.82 ;
 RECT 3.57 1.015 3.71 1.175 ;
 RECT 4.695 1.385 4.835 1.82 ;
 RECT 3.5 0.875 3.78 1.015 ;
 RECT 3.395 1.175 3.71 1.315 ;
 RECT 3.395 1.315 3.535 1.775 ;
 END
END DFFNX2

MACRO DFFSSRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.52 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.52 2.96 ;
 RECT 4.34 2.38 4.59 2.8 ;
 RECT 6.7 2.635 6.96 2.8 ;
 RECT 1.505 1.98 1.645 2.8 ;
 RECT 8.815 1.955 8.955 2.8 ;
 RECT 3.685 1.95 3.825 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 10.29 1.51 10.43 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.52 0.08 ;
 RECT 1.4 0.08 1.7 0.26 ;
 RECT 4.315 0.08 4.615 0.26 ;
 RECT 8.57 0.08 8.825 0.285 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 6.635 0.08 6.775 0.58 ;
 RECT 10.34 0.08 10.48 0.815 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.02 1.475 4.44 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.715 2.085 10.145 2.39 ;
 RECT 9.775 2.39 9.915 2.575 ;
 RECT 9.775 0.56 9.915 2.085 ;
 END
 ANTENNADIFFAREA 0.527 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.775 2.08 11.15 2.385 ;
 RECT 10.82 2.385 10.96 2.575 ;
 RECT 10.82 0.61 10.96 2.08 ;
 END
 ANTENNADIFFAREA 0.47 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.115 1.455 2.495 1.735 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.22 1.48 1.535 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SETB

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.48 0.22 3.74 0.6 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END RSTB

 OBS
 LAYER PO ;
 RECT 5.105 0.185 6.52 0.285 ;
 RECT 5.105 0.285 5.205 0.525 ;
 RECT 6.42 0.285 6.52 1.26 ;
 RECT 5.065 0.525 5.295 0.76 ;
 RECT 2.23 0.745 2.33 1.475 ;
 RECT 2.23 1.71 2.33 2.465 ;
 RECT 2.185 1.475 2.415 1.71 ;
 RECT 5.605 1.675 5.705 2.495 ;
 RECT 5.08 1.49 5.325 1.575 ;
 RECT 5.08 1.675 5.325 1.735 ;
 RECT 5.08 1.575 5.705 1.675 ;
 RECT 4.18 1.3 4.28 1.48 ;
 RECT 4.18 1.2 4.565 1.3 ;
 RECT 4.465 0.64 4.565 1.2 ;
 RECT 3.945 1.72 4.045 2.37 ;
 RECT 3.945 1.48 4.29 1.72 ;
 RECT 8.6 1.64 8.7 2.69 ;
 RECT 7.225 2.385 7.445 2.69 ;
 RECT 7.225 2.69 8.7 2.79 ;
 RECT 2.7 0.745 2.8 1.28 ;
 RECT 2.7 1.28 3.21 1.515 ;
 RECT 6.86 0.66 6.96 1.59 ;
 RECT 6.86 1.82 6.96 2.49 ;
 RECT 6.81 1.59 7.05 1.82 ;
 RECT 1.29 0.74 1.39 1.485 ;
 RECT 1.29 1.72 1.39 2.465 ;
 RECT 1.255 1.485 1.485 1.72 ;
 RECT 8.84 1.205 10.13 1.365 ;
 RECT 9.27 1.135 10.13 1.205 ;
 RECT 8.84 1.365 9.765 1.44 ;
 RECT 8.88 0.5 8.98 1.205 ;
 RECT 9.09 1.44 9.19 2.695 ;
 RECT 10.03 0.195 10.13 1.135 ;
 RECT 10.03 1.365 10.13 2.79 ;
 RECT 1.76 1.775 1.86 2.675 ;
 RECT 0.845 2.375 1.075 2.675 ;
 RECT 0.845 2.675 1.86 2.775 ;
 RECT 10.605 0.245 10.705 1.035 ;
 RECT 10.405 1.035 10.705 1.27 ;
 RECT 10.605 1.27 10.705 2.79 ;
 RECT 7.63 1.505 7.73 2.27 ;
 RECT 7.63 2.27 8.15 2.51 ;
 RECT 7.655 0.685 7.755 1.255 ;
 RECT 7.52 0.455 7.755 0.685 ;
 RECT 6.1 1.33 6.22 1.475 ;
 RECT 6.1 1.71 6.2 2.475 ;
 RECT 5.985 1.475 6.22 1.71 ;
 RECT 6.12 0.65 6.22 1.33 ;
 RECT 8.425 0.265 8.525 1.16 ;
 RECT 6.89 0.265 7.2 0.435 ;
 RECT 8.425 1.16 8.66 1.37 ;
 RECT 6.89 0.165 8.525 0.265 ;
 RECT 7.95 0.445 8.225 0.655 ;
 RECT 8.125 0.655 8.225 2.09 ;
 RECT 3.395 0.46 3.495 0.465 ;
 RECT 1.76 0.465 3.495 0.565 ;
 RECT 3.395 0.565 3.495 1.71 ;
 RECT 1.76 0.565 1.86 1.325 ;
 RECT 2.7 1.81 2.8 2.465 ;
 RECT 2.7 1.71 3.495 1.81 ;
 RECT 3.395 0.225 3.73 0.46 ;
 RECT 4.575 1.49 4.885 1.62 ;
 RECT 4.785 1.255 4.885 1.49 ;
 RECT 4.72 1.735 4.82 2.685 ;
 RECT 6.42 1.78 6.52 2.685 ;
 RECT 4.575 1.62 4.82 1.735 ;
 RECT 5.65 0.705 5.75 1.155 ;
 RECT 4.785 0.685 4.885 1.155 ;
 RECT 5.65 0.47 5.94 0.705 ;
 RECT 4.72 2.685 6.52 2.785 ;
 RECT 4.785 1.155 5.75 1.255 ;
 LAYER CO ;
 RECT 6.035 1.525 6.165 1.655 ;
 RECT 7.28 0.88 7.41 1.01 ;
 RECT 7.28 2.015 7.41 2.145 ;
 RECT 4.435 0.125 4.565 0.255 ;
 RECT 2.45 2.05 2.58 2.18 ;
 RECT 2.45 0.97 2.58 1.1 ;
 RECT 0.895 2.43 1.025 2.56 ;
 RECT 1.51 2.05 1.64 2.18 ;
 RECT 1.98 2.05 2.11 2.18 ;
 RECT 1.98 0.97 2.11 1.1 ;
 RECT 4.215 0.905 4.345 1.035 ;
 RECT 3.69 2 3.82 2.13 ;
 RECT 10.345 0.615 10.475 0.745 ;
 RECT 9.78 2.115 9.91 2.245 ;
 RECT 9.78 2.375 9.91 2.505 ;
 RECT 9.78 0.63 9.91 0.76 ;
 RECT 8.645 0.15 8.775 0.28 ;
 RECT 7.98 2.33 8.11 2.46 ;
 RECT 8.475 1.2 8.605 1.33 ;
 RECT 8 0.485 8.13 0.615 ;
 RECT 9.105 0.87 9.235 1 ;
 RECT 8.82 2.01 8.95 2.14 ;
 RECT 10.825 1.59 10.955 1.72 ;
 RECT 10.295 1.59 10.425 1.72 ;
 RECT 10.295 1.85 10.425 1.98 ;
 RECT 10.295 2.115 10.425 2.245 ;
 RECT 10.295 2.375 10.425 2.505 ;
 RECT 8.895 1.25 9.025 1.38 ;
 RECT 4.94 1.825 5.07 1.955 ;
 RECT 1.52 0.125 1.65 0.255 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 7.275 2.435 7.405 2.565 ;
 RECT 7.28 1.755 7.41 1.885 ;
 RECT 4.41 2.385 4.54 2.515 ;
 RECT 5.85 2.07 5.98 2.2 ;
 RECT 5.87 0.88 6 1.01 ;
 RECT 5.355 2.105 5.485 2.235 ;
 RECT 6.64 0.38 6.77 0.51 ;
 RECT 7.875 1.9 8.005 2.03 ;
 RECT 7.875 0.87 8.005 1 ;
 RECT 7.57 0.505 7.7 0.635 ;
 RECT 3.55 0.28 3.68 0.41 ;
 RECT 9.31 1.965 9.44 2.095 ;
 RECT 9.78 1.59 9.91 1.72 ;
 RECT 9.78 1.85 9.91 1.98 ;
 RECT 4.63 1.535 4.76 1.665 ;
 RECT 5.76 0.525 5.89 0.655 ;
 RECT 7.01 0.255 7.14 0.385 ;
 RECT 6.75 2.64 6.88 2.77 ;
 RECT 5.115 0.58 5.245 0.71 ;
 RECT 2.235 1.53 2.365 1.66 ;
 RECT 10.825 1.85 10.955 1.98 ;
 RECT 10.825 2.115 10.955 2.245 ;
 RECT 10.825 2.375 10.955 2.505 ;
 RECT 5.4 0.88 5.53 1.01 ;
 RECT 5.135 1.535 5.265 1.665 ;
 RECT 5.005 0.905 5.135 1.035 ;
 RECT 4.12 1.535 4.25 1.665 ;
 RECT 4.215 2 4.345 2.13 ;
 RECT 3.03 1.335 3.16 1.465 ;
 RECT 6.865 1.63 6.995 1.76 ;
 RECT 1.305 1.54 1.435 1.67 ;
 RECT 2.92 2.05 3.05 2.18 ;
 RECT 2.92 0.97 3.05 1.1 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 1.04 2.05 1.17 2.18 ;
 RECT 1.04 0.97 1.17 1.1 ;
 RECT 10.445 1.085 10.575 1.215 ;
 RECT 10.825 0.68 10.955 0.81 ;
 LAYER M1 ;
 RECT 5.97 1.52 6.63 1.66 ;
 RECT 6.49 1.185 7.415 1.325 ;
 RECT 7.275 0.81 7.415 1.185 ;
 RECT 7.275 1.325 7.415 2.215 ;
 RECT 6.49 1.325 6.63 1.52 ;
 RECT 1.975 2.465 3.055 2.605 ;
 RECT 2.915 1.98 3.055 2.465 ;
 RECT 1.975 1.98 2.115 2.465 ;
 RECT 0.89 0.54 1.03 0.965 ;
 RECT 0.89 1.105 1.03 2.045 ;
 RECT 0.89 2.185 1.03 2.66 ;
 RECT 0.89 2.045 1.23 2.185 ;
 RECT 0.89 0.965 1.24 1.105 ;
 RECT 2.915 1.33 3.335 1.47 ;
 RECT 3.195 0.54 3.335 1.33 ;
 RECT 0.89 0.4 3.335 0.54 ;
 RECT 5.685 0.52 6.495 0.66 ;
 RECT 6.355 0.66 6.495 0.79 ;
 RECT 6.355 0.79 7.055 0.93 ;
 RECT 6.915 0.25 7.21 0.39 ;
 RECT 6.915 0.39 7.055 0.79 ;
 RECT 1.975 0.825 2.115 0.965 ;
 RECT 1.975 0.685 3.055 0.825 ;
 RECT 2.915 0.825 3.055 1.16 ;
 RECT 1.9 0.965 2.185 1.105 ;
 RECT 8.28 1.195 8.675 1.335 ;
 RECT 8.28 1.335 8.42 2.325 ;
 RECT 7.89 2.325 8.42 2.465 ;
 RECT 7.87 0.82 8.01 0.86 ;
 RECT 7.87 1 8.01 2.135 ;
 RECT 7.87 0.86 8.96 1 ;
 RECT 8.82 1.245 9.095 1.385 ;
 RECT 8.82 1 8.96 1.245 ;
 RECT 4.87 1.82 5.19 1.96 ;
 RECT 5.05 1.96 5.19 2.51 ;
 RECT 5.05 2.51 6.265 2.65 ;
 RECT 5 1.715 5.19 1.82 ;
 RECT 6.125 2.495 6.265 2.51 ;
 RECT 5.11 0.5 5.25 0.84 ;
 RECT 5 0.84 5.25 1.035 ;
 RECT 5 1.035 5.14 1.485 ;
 RECT 5 1.485 5.27 1.715 ;
 RECT 6.125 2.355 7.24 2.43 ;
 RECT 6.125 2.43 7.705 2.495 ;
 RECT 7.1 2.495 7.705 2.57 ;
 RECT 7.565 0.45 7.705 2.43 ;
 RECT 2.635 1.81 2.775 1.9 ;
 RECT 2.445 2.04 2.585 2.255 ;
 RECT 2.37 0.965 2.775 1.105 ;
 RECT 2.635 1.105 2.775 1.67 ;
 RECT 2.445 1.9 2.775 2.04 ;
 RECT 2.635 1.67 3.785 1.81 ;
 RECT 3.645 1.325 3.785 1.67 ;
 RECT 3.925 0.67 4.065 1.185 ;
 RECT 3.645 1.185 4.065 1.325 ;
 RECT 3.925 0.53 4.915 0.67 ;
 RECT 5.395 0.36 5.535 0.8 ;
 RECT 4.775 0.36 4.915 0.53 ;
 RECT 4.775 0.22 5.535 0.36 ;
 RECT 5.395 0.8 5.55 1.095 ;
 RECT 5.41 1.095 5.55 2.035 ;
 RECT 5.35 2.035 5.55 2.305 ;
 RECT 5.775 1.96 6.055 2.215 ;
 RECT 5.865 1.015 6.005 1.22 ;
 RECT 5.69 1.22 6.005 1.36 ;
 RECT 5.69 1.82 7 1.96 ;
 RECT 6.86 1.56 7 1.82 ;
 RECT 5.795 0.875 6.075 1.015 ;
 RECT 5.69 1.36 5.83 1.82 ;
 RECT 4.21 0.835 4.35 1.15 ;
 RECT 4.615 1.29 4.755 1.53 ;
 RECT 4.59 1.675 4.73 1.995 ;
 RECT 4.21 1.15 4.755 1.29 ;
 RECT 4.145 1.995 4.73 2.135 ;
 RECT 4.58 1.53 4.81 1.675 ;
 RECT 9.1 0.965 9.445 1.105 ;
 RECT 9.1 0.63 9.24 0.965 ;
 RECT 9.1 0.36 9.24 0.49 ;
 RECT 7.995 0.49 9.24 0.63 ;
 RECT 9.305 1.105 9.445 2.165 ;
 RECT 7.995 0.425 8.14 0.49 ;
 RECT 7.995 0.63 8.14 0.675 ;
 RECT 10.06 0.36 10.2 1.08 ;
 RECT 9.1 0.22 10.2 0.36 ;
 RECT 10.44 1.01 10.58 1.08 ;
 RECT 10.44 1.22 10.58 1.29 ;
 RECT 10.06 1.08 10.58 1.22 ;
 END
END DFFSSRX1

MACRO DFFSSRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 13.12 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 13.12 2.96 ;
 RECT 4.405 2.38 4.655 2.8 ;
 RECT 6.765 2.635 7.025 2.8 ;
 RECT 10.355 1.765 10.495 2.8 ;
 RECT 1.57 1.98 1.71 2.8 ;
 RECT 12.085 1.765 12.225 2.8 ;
 RECT 8.88 1.955 9.02 2.8 ;
 RECT 3.75 1.95 3.89 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 13.12 0.08 ;
 RECT 4.38 0.08 4.68 0.26 ;
 RECT 12.135 0.08 12.275 0.795 ;
 RECT 1.465 0.08 1.765 0.26 ;
 RECT 8.635 0.08 8.89 0.285 ;
 RECT 10.405 0.08 10.545 0.815 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 6.7 0.08 6.84 0.58 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.085 1.475 4.505 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.84 2.085 10.205 2.39 ;
 RECT 9.84 2.39 9.98 2.575 ;
 RECT 10.965 1.565 11.105 2.575 ;
 RECT 10.965 0.645 11.105 1.425 ;
 RECT 9.84 1.425 11.105 1.565 ;
 RECT 9.84 1.565 9.98 2.085 ;
 RECT 9.84 0.56 9.98 1.425 ;
 END
 ANTENNADIFFAREA 1.089 ;
 END QN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.925 1.455 2.48 1.735 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.285 1.48 1.6 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SETB

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.545 0.22 3.845 0.6 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END RSTB

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.695 0.61 12.835 1.125 ;
 RECT 11.57 1.565 11.71 2.575 ;
 RECT 11.57 0.65 11.71 1.425 ;
 RECT 12.695 1.565 12.835 2.575 ;
 RECT 12.47 1.125 12.835 1.425 ;
 RECT 11.57 1.425 12.835 1.565 ;
 END
 ANTENNADIFFAREA 1.043 ;
 END Q

 OBS
 LAYER PO ;
 RECT 5.145 1.575 5.77 1.675 ;
 RECT 4.245 1.3 4.345 1.48 ;
 RECT 4.245 1.2 4.63 1.3 ;
 RECT 4.53 0.64 4.63 1.2 ;
 RECT 4.01 1.72 4.11 2.37 ;
 RECT 4.01 1.48 4.355 1.72 ;
 RECT 6.925 0.66 7.025 1.59 ;
 RECT 6.925 1.82 7.025 2.49 ;
 RECT 6.875 1.59 7.115 1.82 ;
 RECT 9.335 1.135 10.195 1.205 ;
 RECT 8.905 1.205 10.195 1.325 ;
 RECT 8.905 1.325 10.77 1.365 ;
 RECT 8.905 1.365 9.83 1.44 ;
 RECT 10.095 0.195 10.195 1.135 ;
 RECT 8.945 0.505 9.045 1.205 ;
 RECT 9.155 1.44 9.255 2.695 ;
 RECT 10.095 1.365 10.77 1.425 ;
 RECT 10.095 1.425 10.195 2.79 ;
 RECT 10.67 0.2 10.77 1.325 ;
 RECT 10.67 1.425 10.77 2.79 ;
 RECT 4.64 1.49 4.95 1.62 ;
 RECT 4.785 1.735 4.885 2.685 ;
 RECT 4.85 1.255 4.95 1.49 ;
 RECT 5.715 0.47 6.005 0.705 ;
 RECT 5.715 0.705 5.815 1.155 ;
 RECT 6.485 1.78 6.585 2.685 ;
 RECT 4.85 0.685 4.95 1.155 ;
 RECT 4.64 1.62 4.885 1.735 ;
 RECT 4.785 2.685 6.585 2.785 ;
 RECT 4.85 1.155 5.815 1.255 ;
 RECT 3.46 0.46 3.56 0.465 ;
 RECT 1.825 0.465 3.56 0.565 ;
 RECT 3.46 0.565 3.56 1.71 ;
 RECT 1.825 0.565 1.925 1.325 ;
 RECT 2.765 1.81 2.865 2.465 ;
 RECT 2.765 1.71 3.56 1.81 ;
 RECT 3.46 0.225 3.795 0.46 ;
 RECT 8.015 0.445 8.29 0.655 ;
 RECT 8.19 0.655 8.29 2.09 ;
 RECT 7.72 0.685 7.82 1.255 ;
 RECT 7.585 0.455 7.82 0.685 ;
 RECT 6.185 0.65 6.285 1.475 ;
 RECT 6.185 1.71 6.285 2.475 ;
 RECT 6.05 1.475 6.285 1.71 ;
 RECT 2.765 0.745 2.865 1.28 ;
 RECT 2.765 1.28 3.275 1.515 ;
 RECT 1.825 1.775 1.925 2.675 ;
 RECT 0.91 2.375 1.14 2.675 ;
 RECT 0.91 2.675 1.925 2.775 ;
 RECT 2.295 0.745 2.395 1.475 ;
 RECT 2.295 1.71 2.395 2.465 ;
 RECT 2.25 1.475 2.48 1.71 ;
 RECT 8.665 1.64 8.765 2.69 ;
 RECT 7.29 2.385 7.51 2.69 ;
 RECT 7.29 2.69 8.765 2.79 ;
 RECT 1.355 0.74 1.455 1.485 ;
 RECT 1.355 1.72 1.455 2.465 ;
 RECT 1.32 1.485 1.55 1.72 ;
 RECT 5.17 0.185 6.585 0.285 ;
 RECT 5.17 0.285 5.27 0.525 ;
 RECT 6.485 0.285 6.585 1.26 ;
 RECT 5.13 0.525 5.36 0.76 ;
 RECT 7.695 1.505 7.795 2.27 ;
 RECT 7.695 2.27 8.215 2.51 ;
 RECT 11.825 0.245 11.925 1.325 ;
 RECT 11.825 1.425 11.925 2.79 ;
 RECT 12.4 0.2 12.5 1.325 ;
 RECT 12.4 1.425 12.5 2.79 ;
 RECT 11.185 0.245 11.44 0.48 ;
 RECT 11.825 1.325 12.5 1.425 ;
 RECT 11.185 0.145 11.925 0.245 ;
 RECT 8.49 0.265 8.59 1.16 ;
 RECT 6.955 0.265 7.265 0.435 ;
 RECT 8.49 1.16 8.725 1.37 ;
 RECT 6.955 0.165 8.59 0.265 ;
 RECT 5.67 1.675 5.77 2.495 ;
 RECT 5.145 1.49 5.39 1.575 ;
 RECT 5.145 1.675 5.39 1.735 ;
 LAYER CO ;
 RECT 10.97 2.115 11.1 2.245 ;
 RECT 10.97 2.375 11.1 2.505 ;
 RECT 10.97 1.59 11.1 1.72 ;
 RECT 10.36 1.85 10.49 1.98 ;
 RECT 10.36 2.115 10.49 2.245 ;
 RECT 10.36 2.375 10.49 2.505 ;
 RECT 9.845 1.59 9.975 1.72 ;
 RECT 9.845 1.85 9.975 1.98 ;
 RECT 9.845 0.63 9.975 0.76 ;
 RECT 8.71 0.15 8.84 0.28 ;
 RECT 6.705 0.38 6.835 0.51 ;
 RECT 7.075 0.255 7.205 0.385 ;
 RECT 8.96 1.25 9.09 1.38 ;
 RECT 8.065 0.485 8.195 0.615 ;
 RECT 9.17 0.87 9.3 1 ;
 RECT 6.93 1.63 7.06 1.76 ;
 RECT 6.1 1.525 6.23 1.655 ;
 RECT 7.345 0.88 7.475 1.01 ;
 RECT 7.345 2.015 7.475 2.145 ;
 RECT 4.5 0.125 4.63 0.255 ;
 RECT 7.34 2.435 7.47 2.565 ;
 RECT 7.345 1.755 7.475 1.885 ;
 RECT 5.935 0.88 6.065 1.01 ;
 RECT 5.42 2.105 5.55 2.235 ;
 RECT 5.465 0.88 5.595 1.01 ;
 RECT 5.2 1.535 5.33 1.665 ;
 RECT 4.28 2 4.41 2.13 ;
 RECT 12.09 1.85 12.22 1.98 ;
 RECT 11.575 1.59 11.705 1.72 ;
 RECT 11.575 2.115 11.705 2.245 ;
 RECT 12.7 1.85 12.83 1.98 ;
 RECT 11.575 1.85 11.705 1.98 ;
 RECT 11.575 2.375 11.705 2.505 ;
 RECT 11.575 0.745 11.705 0.875 ;
 RECT 12.7 2.115 12.83 2.245 ;
 RECT 12.7 2.375 12.83 2.505 ;
 RECT 3.095 1.335 3.225 1.465 ;
 RECT 1.585 0.125 1.715 0.255 ;
 RECT 2.515 2.05 2.645 2.18 ;
 RECT 2.515 0.97 2.645 1.1 ;
 RECT 0.96 2.43 1.09 2.56 ;
 RECT 1.105 2.05 1.235 2.18 ;
 RECT 1.105 0.97 1.235 1.1 ;
 RECT 2.3 1.53 2.43 1.66 ;
 RECT 1.37 1.54 1.5 1.67 ;
 RECT 2.985 2.05 3.115 2.18 ;
 RECT 2.985 0.97 3.115 1.1 ;
 RECT 4.695 1.535 4.825 1.665 ;
 RECT 5.825 0.525 5.955 0.655 ;
 RECT 1.575 2.05 1.705 2.18 ;
 RECT 2.045 2.05 2.175 2.18 ;
 RECT 2.045 0.97 2.175 1.1 ;
 RECT 5.005 1.825 5.135 1.955 ;
 RECT 5.18 0.58 5.31 0.71 ;
 RECT 4.28 0.905 4.41 1.035 ;
 RECT 3.755 2 3.885 2.13 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 8.045 2.33 8.175 2.46 ;
 RECT 8.54 1.2 8.67 1.33 ;
 RECT 10.97 1.85 11.1 1.98 ;
 RECT 11.25 0.295 11.38 0.425 ;
 RECT 10.97 0.74 11.1 0.87 ;
 RECT 10.41 0.615 10.54 0.745 ;
 RECT 9.845 2.115 9.975 2.245 ;
 RECT 9.845 2.375 9.975 2.505 ;
 RECT 4.475 2.385 4.605 2.515 ;
 RECT 5.915 2.07 6.045 2.2 ;
 RECT 7.94 1.9 8.07 2.03 ;
 RECT 7.94 0.87 8.07 1 ;
 RECT 7.635 0.505 7.765 0.635 ;
 RECT 5.07 0.905 5.2 1.035 ;
 RECT 4.185 1.535 4.315 1.665 ;
 RECT 8.885 2.01 9.015 2.14 ;
 RECT 9.375 1.965 9.505 2.095 ;
 RECT 12.09 2.115 12.22 2.245 ;
 RECT 12.09 2.375 12.22 2.505 ;
 RECT 12.14 0.615 12.27 0.745 ;
 RECT 6.815 2.64 6.945 2.77 ;
 RECT 12.7 1.59 12.83 1.72 ;
 RECT 12.7 0.68 12.83 0.81 ;
 RECT 3.615 0.28 3.745 0.41 ;
 LAYER M1 ;
 RECT 6.035 1.52 6.695 1.66 ;
 RECT 6.555 1.185 7.48 1.325 ;
 RECT 7.34 0.81 7.48 1.185 ;
 RECT 7.34 1.325 7.48 2.215 ;
 RECT 6.555 1.325 6.695 1.52 ;
 RECT 2.04 2.465 3.12 2.605 ;
 RECT 2.98 1.98 3.12 2.465 ;
 RECT 2.04 1.98 2.18 2.465 ;
 RECT 0.955 0.54 1.095 0.965 ;
 RECT 0.955 1.105 1.095 2.045 ;
 RECT 0.955 2.185 1.095 2.63 ;
 RECT 0.955 2.045 1.295 2.185 ;
 RECT 0.955 0.965 1.305 1.105 ;
 RECT 2.98 1.33 3.4 1.47 ;
 RECT 3.26 0.54 3.4 1.33 ;
 RECT 0.955 0.4 3.4 0.54 ;
 RECT 2.04 0.825 2.18 0.965 ;
 RECT 2.04 0.685 3.12 0.825 ;
 RECT 2.98 0.825 3.12 1.16 ;
 RECT 1.965 0.965 2.25 1.105 ;
 RECT 8.345 1.195 8.74 1.335 ;
 RECT 8.345 1.335 8.485 2.325 ;
 RECT 7.955 2.325 8.485 2.465 ;
 RECT 5.75 0.52 6.56 0.66 ;
 RECT 6.42 0.66 6.56 0.79 ;
 RECT 6.42 0.79 7.12 0.93 ;
 RECT 6.98 0.25 7.275 0.39 ;
 RECT 6.98 0.39 7.12 0.79 ;
 RECT 4.935 1.82 5.255 1.96 ;
 RECT 5.115 1.96 5.255 2.51 ;
 RECT 5.115 2.51 6.33 2.65 ;
 RECT 5.065 1.715 5.255 1.82 ;
 RECT 6.19 2.495 6.33 2.51 ;
 RECT 5.175 0.5 5.315 0.84 ;
 RECT 5.065 0.84 5.315 1.035 ;
 RECT 5.065 1.035 5.205 1.485 ;
 RECT 5.065 1.485 5.335 1.715 ;
 RECT 7.165 2.495 7.77 2.57 ;
 RECT 6.19 2.355 7.305 2.43 ;
 RECT 6.19 2.43 7.77 2.495 ;
 RECT 7.63 0.45 7.77 2.43 ;
 RECT 2.7 1.81 2.84 1.9 ;
 RECT 2.51 2.04 2.65 2.255 ;
 RECT 2.435 0.965 2.84 1.105 ;
 RECT 2.7 1.105 2.84 1.67 ;
 RECT 2.51 1.9 2.84 2.04 ;
 RECT 2.7 1.67 3.85 1.81 ;
 RECT 3.71 1.325 3.85 1.67 ;
 RECT 3.99 0.67 4.13 1.185 ;
 RECT 3.71 1.185 4.13 1.325 ;
 RECT 3.99 0.53 4.98 0.67 ;
 RECT 5.46 0.36 5.6 0.8 ;
 RECT 4.84 0.36 4.98 0.53 ;
 RECT 4.84 0.22 5.6 0.36 ;
 RECT 5.46 0.8 5.615 1.095 ;
 RECT 5.475 1.095 5.615 2.035 ;
 RECT 5.415 2.035 5.615 2.305 ;
 RECT 4.275 0.835 4.415 1.15 ;
 RECT 4.68 1.29 4.82 1.53 ;
 RECT 4.655 1.675 4.795 1.995 ;
 RECT 4.275 1.15 4.82 1.29 ;
 RECT 4.21 1.995 4.795 2.135 ;
 RECT 4.645 1.53 4.875 1.675 ;
 RECT 5.84 1.96 6.12 2.215 ;
 RECT 5.93 1.015 6.07 1.22 ;
 RECT 5.755 1.22 6.07 1.36 ;
 RECT 5.755 1.82 7.065 1.96 ;
 RECT 6.925 1.56 7.065 1.82 ;
 RECT 5.86 0.875 6.14 1.015 ;
 RECT 5.755 1.36 5.895 1.82 ;
 RECT 7.935 0.82 8.075 0.86 ;
 RECT 7.935 1 8.075 2.135 ;
 RECT 7.935 0.86 9.025 1 ;
 RECT 8.885 1.245 9.16 1.385 ;
 RECT 8.885 1 9.025 1.245 ;
 RECT 10.125 0.36 10.265 0.955 ;
 RECT 9.165 0.22 10.265 0.36 ;
 RECT 10.685 0.43 10.825 0.955 ;
 RECT 10.125 0.955 10.825 1.095 ;
 RECT 10.685 0.285 10.825 0.29 ;
 RECT 9.165 0.965 9.51 1.105 ;
 RECT 9.165 0.63 9.305 0.965 ;
 RECT 9.165 0.36 9.305 0.49 ;
 RECT 8.06 0.49 9.305 0.63 ;
 RECT 9.37 1.105 9.51 2.165 ;
 RECT 8.06 0.425 8.205 0.49 ;
 RECT 8.06 0.63 8.205 0.675 ;
 RECT 11.245 0.22 11.385 0.29 ;
 RECT 11.245 0.43 11.385 0.5 ;
 RECT 10.685 0.29 11.485 0.43 ;
 END
END DFFSSRX2

MACRO DFFX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.64 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.64 2.96 ;
 RECT 1.915 2.38 2.165 2.8 ;
 RECT 4.275 2.635 4.535 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 7.865 1.51 8.005 2.8 ;
 RECT 1.26 1.98 1.4 2.8 ;
 RECT 6.39 1.955 6.53 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.64 0.08 ;
 RECT 1.26 0.08 1.4 1.055 ;
 RECT 1.89 0.08 2.19 0.26 ;
 RECT 6.145 0.08 6.4 0.285 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.21 0.08 4.35 0.58 ;
 RECT 7.915 0.08 8.055 0.815 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.595 1.475 1.91 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.35 2.085 7.64 2.39 ;
 RECT 7.35 2.39 7.49 2.575 ;
 RECT 7.35 0.56 7.49 2.085 ;
 END
 ANTENNADIFFAREA 0.527 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.2 2.08 8.535 2.385 ;
 RECT 8.395 2.385 8.535 2.575 ;
 RECT 8.395 0.61 8.535 2.08 ;
 END
 ANTENNADIFFAREA 0.47 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.975 1.475 1.24 1.785 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 OBS
 LAYER PO ;
 RECT 1.52 0.655 1.62 1.48 ;
 RECT 1.52 1.72 1.62 2.37 ;
 RECT 1.52 1.48 1.865 1.72 ;
 RECT 2.68 0.185 4.095 0.285 ;
 RECT 2.68 0.285 2.78 0.525 ;
 RECT 3.995 0.285 4.095 1.26 ;
 RECT 2.64 0.525 2.87 0.76 ;
 RECT 3.18 1.675 3.28 2.495 ;
 RECT 2.655 1.49 2.9 1.575 ;
 RECT 2.655 1.575 3.28 1.675 ;
 RECT 2.655 1.675 2.9 1.735 ;
 RECT 6 0.265 6.1 1.16 ;
 RECT 4.675 0.165 6.1 0.205 ;
 RECT 4.435 0.205 6.1 0.265 ;
 RECT 4.435 0.265 4.775 0.435 ;
 RECT 6 1.16 6.235 1.37 ;
 RECT 5.525 0.445 5.8 0.655 ;
 RECT 5.7 0.655 5.8 2.09 ;
 RECT 5.23 0.685 5.33 1.255 ;
 RECT 5.095 0.455 5.33 0.685 ;
 RECT 4.435 0.66 4.535 1.59 ;
 RECT 4.435 1.82 4.535 2.49 ;
 RECT 4.385 1.59 4.625 1.82 ;
 RECT 3.675 1.33 3.795 1.475 ;
 RECT 3.675 1.71 3.775 2.475 ;
 RECT 3.56 1.475 3.795 1.71 ;
 RECT 3.695 0.65 3.795 1.33 ;
 RECT 6.415 1.205 7.705 1.365 ;
 RECT 6.845 1.135 7.705 1.205 ;
 RECT 6.415 1.365 7.34 1.44 ;
 RECT 6.455 0.65 6.555 1.205 ;
 RECT 6.665 1.44 6.765 2.51 ;
 RECT 7.605 0.195 7.705 1.135 ;
 RECT 7.605 1.365 7.705 2.79 ;
 RECT 8.18 0.26 8.28 1.035 ;
 RECT 8.18 1.27 8.28 2.79 ;
 RECT 7.98 1.035 8.28 1.27 ;
 RECT 2.15 1.49 2.46 1.62 ;
 RECT 2.295 1.735 2.395 2.685 ;
 RECT 2.36 1.255 2.46 1.49 ;
 RECT 3.225 0.47 3.515 0.705 ;
 RECT 3.225 0.705 3.325 1.155 ;
 RECT 3.995 1.78 4.095 2.685 ;
 RECT 2.36 0.685 2.46 1.155 ;
 RECT 2.15 1.62 2.395 1.735 ;
 RECT 2.295 2.685 4.095 2.785 ;
 RECT 2.36 1.155 3.325 1.255 ;
 RECT 5.205 1.465 5.305 2.27 ;
 RECT 5.205 2.27 5.725 2.51 ;
 RECT 1.045 0.655 1.145 1.475 ;
 RECT 1.045 1.71 1.145 2.465 ;
 RECT 1.045 1.475 1.275 1.71 ;
 RECT 6.175 1.64 6.275 2.69 ;
 RECT 4.8 2.385 5.02 2.69 ;
 RECT 4.8 2.69 6.275 2.79 ;
 LAYER CO ;
 RECT 3.445 0.88 3.575 1.01 ;
 RECT 2.93 2.105 3.06 2.235 ;
 RECT 2.975 0.88 3.105 1.01 ;
 RECT 2.71 1.535 2.84 1.665 ;
 RECT 2.58 0.905 2.71 1.035 ;
 RECT 1.695 1.535 1.825 1.665 ;
 RECT 1.79 1.995 1.92 2.125 ;
 RECT 1.87 0.875 2 1.005 ;
 RECT 1.265 2.05 1.395 2.18 ;
 RECT 1.265 0.875 1.395 1.005 ;
 RECT 1.095 1.53 1.225 1.66 ;
 RECT 0.795 2.05 0.925 2.18 ;
 RECT 0.795 0.875 0.925 1.005 ;
 RECT 5.555 2.33 5.685 2.46 ;
 RECT 6.05 1.2 6.18 1.33 ;
 RECT 8.4 1.85 8.53 1.98 ;
 RECT 8.4 2.115 8.53 2.245 ;
 RECT 8.4 2.375 8.53 2.505 ;
 RECT 8.4 1.59 8.53 1.72 ;
 RECT 7.87 1.59 8 1.72 ;
 RECT 7.87 1.85 8 1.98 ;
 RECT 7.87 2.115 8 2.245 ;
 RECT 7.87 2.375 8 2.505 ;
 RECT 7.355 1.59 7.485 1.72 ;
 RECT 7.355 1.85 7.485 1.98 ;
 RECT 2.205 1.535 2.335 1.665 ;
 RECT 3.335 0.525 3.465 0.655 ;
 RECT 4.585 0.255 4.715 0.385 ;
 RECT 6.47 1.25 6.6 1.38 ;
 RECT 2.515 1.825 2.645 1.955 ;
 RECT 2.69 0.58 2.82 0.71 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 4.85 2.435 4.98 2.565 ;
 RECT 4.855 1.755 4.985 1.885 ;
 RECT 8.02 1.085 8.15 1.215 ;
 RECT 8.4 0.68 8.53 0.81 ;
 RECT 7.92 0.615 8.05 0.745 ;
 RECT 7.355 2.115 7.485 2.245 ;
 RECT 7.355 2.375 7.485 2.505 ;
 RECT 7.355 0.63 7.485 0.76 ;
 RECT 6.22 0.15 6.35 0.28 ;
 RECT 4.215 0.38 4.345 0.51 ;
 RECT 5.45 1.9 5.58 2.03 ;
 RECT 5.45 0.87 5.58 1 ;
 RECT 5.145 0.505 5.275 0.635 ;
 RECT 5.575 0.485 5.705 0.615 ;
 RECT 6.68 0.87 6.81 1 ;
 RECT 6.395 2.01 6.525 2.14 ;
 RECT 6.885 1.965 7.015 2.095 ;
 RECT 4.44 1.63 4.57 1.76 ;
 RECT 3.61 1.525 3.74 1.655 ;
 RECT 4.855 0.88 4.985 1.01 ;
 RECT 4.855 2.015 4.985 2.145 ;
 RECT 2.01 0.125 2.14 0.255 ;
 RECT 4.325 2.64 4.455 2.77 ;
 RECT 1.985 2.385 2.115 2.515 ;
 RECT 3.425 2.07 3.555 2.2 ;
 LAYER M1 ;
 RECT 5.855 1.195 6.25 1.335 ;
 RECT 5.855 1.335 5.995 2.325 ;
 RECT 5.465 2.325 5.995 2.465 ;
 RECT 3.26 0.52 4.07 0.66 ;
 RECT 3.93 0.66 4.07 0.79 ;
 RECT 3.93 0.79 4.63 0.93 ;
 RECT 4.49 0.25 4.785 0.39 ;
 RECT 4.49 0.39 4.63 0.79 ;
 RECT 3.545 1.52 4.205 1.66 ;
 RECT 4.065 1.185 4.99 1.325 ;
 RECT 4.85 0.81 4.99 1.185 ;
 RECT 4.85 1.325 4.99 2.215 ;
 RECT 4.065 1.325 4.205 1.52 ;
 RECT 2.19 1.01 2.33 1.53 ;
 RECT 2.165 1.675 2.305 1.99 ;
 RECT 1.82 0.87 2.33 1.01 ;
 RECT 1.72 1.99 2.305 2.13 ;
 RECT 2.155 1.53 2.385 1.675 ;
 RECT 6.675 0.965 7.02 1.105 ;
 RECT 6.675 0.63 6.815 0.965 ;
 RECT 6.675 0.36 6.815 0.49 ;
 RECT 5.57 0.49 6.815 0.63 ;
 RECT 6.88 1.105 7.02 2.165 ;
 RECT 5.57 0.425 5.715 0.49 ;
 RECT 5.57 0.63 5.715 0.675 ;
 RECT 7.635 0.36 7.775 1.08 ;
 RECT 6.675 0.22 7.775 0.36 ;
 RECT 8.015 1.01 8.155 1.08 ;
 RECT 8.015 1.22 8.155 1.29 ;
 RECT 7.635 1.08 8.155 1.22 ;
 RECT 5.445 0.82 5.585 0.86 ;
 RECT 5.445 1 5.585 2.11 ;
 RECT 5.445 0.86 6.535 1 ;
 RECT 6.395 1.245 6.67 1.385 ;
 RECT 6.395 1 6.535 1.245 ;
 RECT 2.445 1.82 2.765 1.96 ;
 RECT 2.625 1.96 2.765 2.51 ;
 RECT 2.625 2.51 3.84 2.65 ;
 RECT 2.575 1.715 2.765 1.82 ;
 RECT 3.7 2.495 3.84 2.51 ;
 RECT 2.685 0.5 2.825 0.84 ;
 RECT 2.575 0.84 2.825 1.035 ;
 RECT 2.575 1.035 2.715 1.485 ;
 RECT 2.575 1.485 2.845 1.715 ;
 RECT 4.675 2.495 5.28 2.57 ;
 RECT 3.7 2.355 4.815 2.43 ;
 RECT 3.7 2.43 5.28 2.495 ;
 RECT 5.14 0.45 5.28 2.43 ;
 RECT 0.58 1.01 0.72 1.195 ;
 RECT 0.58 1.335 0.72 2.045 ;
 RECT 1.54 0.67 1.68 1.195 ;
 RECT 0.58 1.195 1.68 1.335 ;
 RECT 0.58 0.87 1 1.01 ;
 RECT 0.58 2.045 1 2.185 ;
 RECT 1.54 0.53 2.49 0.67 ;
 RECT 2.97 0.36 3.11 0.8 ;
 RECT 2.35 0.36 2.49 0.53 ;
 RECT 2.35 0.22 3.11 0.36 ;
 RECT 2.97 0.8 3.125 1.095 ;
 RECT 2.985 1.095 3.125 2.035 ;
 RECT 2.925 2.035 3.125 2.305 ;
 RECT 3.265 1.82 4.575 1.96 ;
 RECT 3.44 1.015 3.58 1.22 ;
 RECT 4.435 1.56 4.575 1.82 ;
 RECT 3.265 1.22 3.58 1.36 ;
 RECT 3.35 1.96 3.63 2.215 ;
 RECT 3.37 0.875 3.65 1.015 ;
 RECT 3.265 1.36 3.405 1.82 ;
 END
END DFFX1

MACRO DFFX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.88 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.88 2.96 ;
 RECT 2.045 2.38 2.295 2.8 ;
 RECT 4.405 2.635 4.665 2.8 ;
 RECT 1.39 1.98 1.53 2.8 ;
 RECT 7.315 1.955 7.455 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 8.595 1.54 8.735 2.8 ;
 RECT 9.615 1.54 9.755 2.8 ;
 RECT 10.555 1.54 10.695 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.88 0.08 ;
 RECT 2.02 0.08 2.32 0.39 ;
 RECT 7.32 0.08 7.575 0.535 ;
 RECT 9.545 0.08 9.8 0.3 ;
 RECT 1.39 0.08 1.53 1.055 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.34 0.08 4.48 0.58 ;
 RECT 8.58 0.08 8.72 0.6 ;
 RECT 10.555 0.08 10.695 0.685 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.495 1.475 2.025 1.735 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.95 2.12 9.28 2.39 ;
 RECT 9.14 2.39 9.28 2.575 ;
 RECT 9.14 0.72 9.28 2.12 ;
 END
 ANTENNADIFFAREA 0.748 ;
 END QN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.95 1.475 1.32 1.785 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.895 2.1 10.225 2.35 ;
 RECT 10.085 2.35 10.225 2.575 ;
 RECT 10.085 0.72 10.225 2.1 ;
 END
 ANTENNADIFFAREA 0.622 ;
 END Q

 OBS
 LAYER PO ;
 RECT 8.85 1.35 8.95 2.79 ;
 RECT 5.035 0.575 5.94 0.675 ;
 RECT 5.84 0.675 5.94 1.35 ;
 RECT 7.175 0.265 7.275 1.32 ;
 RECT 5.035 0.46 5.265 0.575 ;
 RECT 5.035 0.675 5.265 0.69 ;
 RECT 5.84 0.265 5.94 0.575 ;
 RECT 6.285 1.545 6.385 2.48 ;
 RECT 5.84 0.165 7.275 0.265 ;
 RECT 5.84 1.35 6.13 1.445 ;
 RECT 5.84 1.445 6.385 1.45 ;
 RECT 6.03 1.45 6.385 1.545 ;
 RECT 1.175 0.655 1.275 1.515 ;
 RECT 1.175 1.745 1.275 2.465 ;
 RECT 1.055 1.515 1.275 1.745 ;
 RECT 4.565 0.635 4.665 1.59 ;
 RECT 4.565 1.59 4.885 1.82 ;
 RECT 4.565 1.82 4.665 2.49 ;
 RECT 3.805 1.33 3.925 1.475 ;
 RECT 3.805 1.71 3.905 2.475 ;
 RECT 3.69 1.475 3.925 1.71 ;
 RECT 3.825 0.65 3.925 1.33 ;
 RECT 5.26 0.875 5.59 1.105 ;
 RECT 5.49 1.105 5.59 1.64 ;
 RECT 5.49 1.64 5.725 1.87 ;
 RECT 3.31 1.675 3.41 2.495 ;
 RECT 2.785 1.49 3.03 1.575 ;
 RECT 2.785 1.675 3.03 1.735 ;
 RECT 2.785 1.575 3.41 1.675 ;
 RECT 7.1 1.64 7.2 2.69 ;
 RECT 5.88 2.47 6.1 2.69 ;
 RECT 5.88 2.69 7.2 2.79 ;
 RECT 2.28 1.49 2.59 1.62 ;
 RECT 2.425 1.735 2.525 2.685 ;
 RECT 2.49 1.255 2.59 1.49 ;
 RECT 3.355 0.47 3.645 0.705 ;
 RECT 3.355 0.705 3.455 1.155 ;
 RECT 4.125 1.78 4.225 2.685 ;
 RECT 2.49 0.685 2.59 1.155 ;
 RECT 2.28 1.62 2.525 1.735 ;
 RECT 2.425 2.685 4.225 2.785 ;
 RECT 2.49 1.155 3.455 1.255 ;
 RECT 1.65 0.655 1.75 1.48 ;
 RECT 1.455 1.48 1.75 1.72 ;
 RECT 1.65 1.72 1.75 2.37 ;
 RECT 6.78 0.645 6.88 1.24 ;
 RECT 6.78 1.45 6.88 2.255 ;
 RECT 6.76 1.24 6.995 1.45 ;
 RECT 6.31 0.685 6.41 1.255 ;
 RECT 6.235 0.455 6.465 0.685 ;
 RECT 7.59 0.65 7.69 1.48 ;
 RECT 7.59 1.72 7.69 2.56 ;
 RECT 7.495 1.48 7.725 1.72 ;
 RECT 10.34 0.2 10.44 1.225 ;
 RECT 9.87 1.325 9.97 2.79 ;
 RECT 10.34 1.325 10.44 2.79 ;
 RECT 9.76 1.225 10.44 1.27 ;
 RECT 9.76 1.035 9.97 1.225 ;
 RECT 9.87 1.27 10.44 1.325 ;
 RECT 9.87 0.2 9.97 1.035 ;
 RECT 2.81 0.185 4.225 0.285 ;
 RECT 2.81 0.285 2.91 0.525 ;
 RECT 4.125 0.285 4.225 1.26 ;
 RECT 2.77 0.525 3 0.76 ;
 RECT 8.115 1.12 8.95 1.225 ;
 RECT 8.115 1.325 8.95 1.35 ;
 RECT 9.395 0.2 9.495 1.225 ;
 RECT 9.395 1.325 9.495 2.79 ;
 RECT 8.115 1.225 9.495 1.325 ;
 RECT 8.85 0.195 8.95 1.12 ;
 LAYER CO ;
 RECT 2.71 0.905 2.84 1.035 ;
 RECT 1.505 1.535 1.635 1.665 ;
 RECT 1.92 1.995 2.05 2.125 ;
 RECT 2 0.875 2.13 1.005 ;
 RECT 1.395 2.05 1.525 2.18 ;
 RECT 9.145 1.85 9.275 1.98 ;
 RECT 2.645 1.825 2.775 1.955 ;
 RECT 8.585 0.42 8.715 0.55 ;
 RECT 8.6 1.59 8.73 1.72 ;
 RECT 0.925 0.875 1.055 1.005 ;
 RECT 0.925 2.05 1.055 2.18 ;
 RECT 8.6 1.85 8.73 1.98 ;
 RECT 8.6 2.115 8.73 2.245 ;
 RECT 10.56 2.375 10.69 2.505 ;
 RECT 10.09 1.85 10.22 1.98 ;
 RECT 10.09 2.115 10.22 2.245 ;
 RECT 10.09 2.375 10.22 2.505 ;
 RECT 10.09 1.59 10.22 1.72 ;
 RECT 10.09 0.77 10.22 0.9 ;
 RECT 9.62 0.165 9.75 0.295 ;
 RECT 9.145 2.375 9.275 2.505 ;
 RECT 9.145 0.77 9.275 0.9 ;
 RECT 3.555 2.07 3.685 2.2 ;
 RECT 1.105 1.565 1.235 1.695 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 10.56 0.505 10.69 0.635 ;
 RECT 7.81 0.87 7.94 1 ;
 RECT 7.32 2.01 7.45 2.14 ;
 RECT 7.88 2.13 8.01 2.26 ;
 RECT 3.465 0.525 3.595 0.655 ;
 RECT 5.075 0.51 5.205 0.64 ;
 RECT 7.55 1.535 7.68 1.665 ;
 RECT 4.455 2.64 4.585 2.77 ;
 RECT 9.62 2.115 9.75 2.245 ;
 RECT 9.62 2.375 9.75 2.505 ;
 RECT 5.545 1.69 5.675 1.82 ;
 RECT 5.33 0.915 5.46 1.045 ;
 RECT 7.395 0.4 7.525 0.53 ;
 RECT 4.345 0.38 4.475 0.51 ;
 RECT 6.53 1.9 6.66 2.03 ;
 RECT 6.53 0.87 6.66 1 ;
 RECT 6.06 0.87 6.19 1 ;
 RECT 6.285 0.505 6.415 0.635 ;
 RECT 8.6 2.375 8.73 2.505 ;
 RECT 9.145 1.59 9.275 1.72 ;
 RECT 5.93 2.525 6.06 2.655 ;
 RECT 6.035 1.815 6.165 1.945 ;
 RECT 9.8 1.085 9.93 1.215 ;
 RECT 8.165 1.17 8.295 1.3 ;
 RECT 9.145 2.115 9.275 2.245 ;
 RECT 2.115 2.385 2.245 2.515 ;
 RECT 2.82 0.58 2.95 0.71 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 10.56 1.59 10.69 1.72 ;
 RECT 10.56 1.85 10.69 1.98 ;
 RECT 10.56 2.115 10.69 2.245 ;
 RECT 4.7 1.63 4.83 1.76 ;
 RECT 3.74 1.525 3.87 1.655 ;
 RECT 4.99 0.88 5.12 1.01 ;
 RECT 4.985 2.015 5.115 2.145 ;
 RECT 2.14 0.255 2.27 0.385 ;
 RECT 9.62 1.59 9.75 1.72 ;
 RECT 9.62 1.85 9.75 1.98 ;
 RECT 3.575 0.88 3.705 1.01 ;
 RECT 3.06 2.105 3.19 2.235 ;
 RECT 3.105 0.88 3.235 1.01 ;
 RECT 2.84 1.535 2.97 1.665 ;
 RECT 1.395 0.875 1.525 1.005 ;
 RECT 6.81 1.28 6.94 1.41 ;
 RECT 2.335 1.535 2.465 1.665 ;
 LAYER M1 ;
 RECT 4.98 1.05 5.12 1.185 ;
 RECT 4.98 1.325 5.12 2.215 ;
 RECT 4.195 1.185 5.12 1.325 ;
 RECT 3.675 1.52 4.335 1.66 ;
 RECT 4.98 1.015 5.53 1.05 ;
 RECT 4.195 1.325 4.335 1.52 ;
 RECT 4.92 0.875 5.53 1.015 ;
 RECT 3.39 0.52 4.2 0.66 ;
 RECT 4.06 0.66 4.2 0.79 ;
 RECT 4.62 0.505 5.275 0.645 ;
 RECT 4.06 0.79 4.76 0.93 ;
 RECT 4.62 0.645 4.76 0.79 ;
 RECT 2.575 1.82 2.895 1.96 ;
 RECT 2.755 1.96 2.895 2.51 ;
 RECT 2.755 2.51 3.97 2.65 ;
 RECT 2.705 1.715 2.895 1.82 ;
 RECT 3.83 2.495 3.97 2.51 ;
 RECT 2.815 0.5 2.955 0.84 ;
 RECT 2.705 0.84 2.955 1.035 ;
 RECT 2.705 1.035 2.845 1.485 ;
 RECT 2.705 1.485 2.975 1.715 ;
 RECT 5.26 1.21 5.84 1.35 ;
 RECT 5.26 1.35 5.4 2.1 ;
 RECT 5.26 2.1 6 2.24 ;
 RECT 5.26 2.24 5.4 2.355 ;
 RECT 5.86 2.24 6 2.52 ;
 RECT 3.83 2.355 5.4 2.495 ;
 RECT 5.98 0.5 6.49 0.58 ;
 RECT 5.7 0.58 6.49 0.64 ;
 RECT 5.7 0.64 6.16 0.72 ;
 RECT 5.86 2.52 6.13 2.66 ;
 RECT 5.7 0.72 5.84 1.21 ;
 RECT 0.67 1.01 0.81 1.195 ;
 RECT 0.67 1.335 0.81 2.045 ;
 RECT 0.67 0.87 1.125 1.01 ;
 RECT 0.67 2.045 1.125 2.185 ;
 RECT 0.67 1.195 1.81 1.335 ;
 RECT 1.67 0.67 1.81 1.195 ;
 RECT 1.67 0.53 2.62 0.67 ;
 RECT 3.1 0.36 3.24 0.8 ;
 RECT 2.48 0.36 2.62 0.53 ;
 RECT 2.48 0.22 3.24 0.36 ;
 RECT 3.1 0.8 3.255 1.095 ;
 RECT 3.115 1.095 3.255 2.035 ;
 RECT 3.055 2.035 3.255 2.305 ;
 RECT 8.86 0.58 9 0.84 ;
 RECT 7.805 0.84 9 0.98 ;
 RECT 6.805 1.245 8.015 1.385 ;
 RECT 7.875 1.105 8.015 1.245 ;
 RECT 7.875 1.385 8.015 2.33 ;
 RECT 7.805 0.76 7.945 0.84 ;
 RECT 7.805 0.98 8.015 1.105 ;
 RECT 6.805 1.21 6.945 1.245 ;
 RECT 6.805 1.385 6.945 1.465 ;
 RECT 9.795 0.58 9.935 1.29 ;
 RECT 8.86 0.44 9.935 0.58 ;
 RECT 6.525 1.815 6.735 1.895 ;
 RECT 6.525 0.805 6.665 1.675 ;
 RECT 6.455 1.895 6.735 2.035 ;
 RECT 6.525 1.675 7.385 1.815 ;
 RECT 7.245 1.67 7.385 1.675 ;
 RECT 8.16 1.12 8.3 2.505 ;
 RECT 7.245 1.53 7.735 1.67 ;
 RECT 7.595 2.505 8.3 2.645 ;
 RECT 7.595 1.67 7.735 2.505 ;
 RECT 5.54 1.685 6.195 1.81 ;
 RECT 6.055 1.005 6.195 1.685 ;
 RECT 5.54 1.81 6.235 1.825 ;
 RECT 5.54 1.825 5.68 1.89 ;
 RECT 5.54 1.62 5.68 1.685 ;
 RECT 5.965 1.825 6.235 1.95 ;
 RECT 5.985 0.865 6.265 1.005 ;
 RECT 3.48 1.96 3.76 2.215 ;
 RECT 3.57 1.015 3.71 1.22 ;
 RECT 3.395 1.22 3.71 1.36 ;
 RECT 3.395 1.82 4.835 1.96 ;
 RECT 4.695 1.56 4.835 1.82 ;
 RECT 3.5 0.875 3.78 1.015 ;
 RECT 3.395 1.36 3.535 1.82 ;
 RECT 1.995 1.045 2.305 1.185 ;
 RECT 2.165 1.185 2.305 1.53 ;
 RECT 1.995 0.81 2.135 1.045 ;
 RECT 2.295 1.67 2.435 1.99 ;
 RECT 1.85 1.99 2.435 2.13 ;
 RECT 2.165 1.53 2.535 1.67 ;
 END
END DFFX2

MACRO FADDX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.24 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.24 2.96 ;
 RECT 4.455 2.14 4.725 2.28 ;
 RECT 3.575 2.075 3.715 2.8 ;
 RECT 8.275 1.9 8.415 2.8 ;
 RECT 9.855 1.9 9.995 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.26 2.095 1.4 2.8 ;
 RECT 4.52 2.28 4.66 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.24 0.08 ;
 RECT 8.475 0.08 8.615 0.34 ;
 RECT 4.44 0.08 4.745 0.245 ;
 RECT 3.485 0.08 3.8 0.28 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 9.855 0.08 9.995 0.795 ;
 RECT 1.26 0.08 1.4 0.41 ;
 END
 END VSS

 PIN A
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.75 2.415 6.34 2.66 ;
 END
 ANTENNAGATEAREA 0.476 ;
 END A

 PIN B
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.015 0.365 2.155 0.965 ;
 RECT 2.015 0.225 3.085 0.365 ;
 RECT 5.34 0.36 5.48 0.665 ;
 RECT 7.88 0.82 8.41 0.96 ;
 RECT 7.295 1.615 8.41 1.755 ;
 RECT 7.28 1.05 7.435 1.195 ;
 RECT 1.27 0.965 2.155 1.105 ;
 RECT 1.27 1.105 1.715 1.505 ;
 RECT 1.27 0.93 1.715 0.965 ;
 RECT 7.88 0.36 8.02 0.82 ;
 RECT 5.34 0.22 8.02 0.36 ;
 RECT 8.27 0.96 8.41 1.615 ;
 RECT 7.295 1.195 7.435 1.615 ;
 RECT 7.295 0.985 7.435 1.05 ;
 RECT 2.945 0.85 3.195 1.02 ;
 RECT 2.945 0.365 3.085 0.665 ;
 RECT 2.945 0.665 5.48 0.85 ;
 END
 ANTENNAGATEAREA 0.476 ;
 END B

 PIN CI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.4 3.55 1.435 ;
 RECT 3.195 1.16 3.55 1.26 ;
 RECT 2.585 1.035 2.725 1.26 ;
 RECT 5.625 1.85 6.815 1.99 ;
 RECT 6.645 1.095 6.815 1.4 ;
 RECT 4.665 1.175 5.765 1.26 ;
 RECT 2.585 1.315 4.945 1.4 ;
 RECT 2.585 1.26 5.765 1.315 ;
 RECT 4.735 1.105 4.875 1.175 ;
 RECT 5.625 1.315 5.765 1.85 ;
 RECT 6.675 1.4 6.815 1.85 ;
 END
 ANTENNAGATEAREA 0.357 ;
 END CI

 PIN CO
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.385 1.43 9.525 2.085 ;
 RECT 9.385 1.155 9.95 1.43 ;
 RECT 9.385 0.595 9.525 1.155 ;
 END
 ANTENNADIFFAREA 0.464 ;
 END CO

 PIN S
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.56 2.035 9.175 2.405 ;
 RECT 9.035 0.595 9.175 2.035 ;
 END
 ANTENNADIFFAREA 0.477 ;
 END S

 OBS
 LAYER PO ;
 RECT 4.775 0.095 4.875 1.135 ;
 RECT 4.775 1.345 4.875 2.51 ;
 RECT 4.69 1.135 4.92 1.345 ;
 RECT 1.515 0.285 1.615 0.93 ;
 RECT 1.515 1.14 1.615 2.51 ;
 RECT 1.485 0.93 1.715 1.14 ;
 RECT 2.105 0.285 2.205 1.065 ;
 RECT 2.105 1.275 2.205 2.51 ;
 RECT 2.105 1.065 2.77 1.275 ;
 RECT 8.815 0.215 8.915 1.135 ;
 RECT 7.935 1.135 8.915 1.345 ;
 RECT 8.815 1.345 8.915 2.79 ;
 RECT 7.02 0.375 7.12 1.02 ;
 RECT 7.02 1.23 7.12 2.51 ;
 RECT 7.02 1.02 7.475 1.23 ;
 RECT 4.305 0.09 4.405 0.67 ;
 RECT 4.135 0.67 4.405 0.88 ;
 RECT 4.305 0.88 4.405 2.51 ;
 RECT 1.045 0.285 1.145 2.69 ;
 RECT 5.855 2.4 6.085 2.69 ;
 RECT 3.83 0.105 3.93 2.69 ;
 RECT 7.655 0.375 7.755 2.69 ;
 RECT 3.36 0.285 3.46 2.69 ;
 RECT 1.045 2.69 7.755 2.79 ;
 RECT 5.25 0.195 5.35 0.97 ;
 RECT 5.25 1.07 5.35 2.51 ;
 RECT 6.185 0.94 6.415 0.97 ;
 RECT 6.185 1.07 6.415 1.15 ;
 RECT 5.25 0.095 8.355 0.195 ;
 RECT 8.11 0.195 8.355 0.5 ;
 RECT 5.25 0.97 6.415 1.07 ;
 RECT 9.64 0.4 9.74 2.79 ;
 RECT 9.275 0.14 9.74 0.4 ;
 RECT 6.715 0.375 6.815 1.115 ;
 RECT 6.715 1.345 6.815 2.51 ;
 RECT 6.595 1.115 6.84 1.345 ;
 RECT 2.99 0.285 3.09 0.845 ;
 RECT 2.99 1.055 3.09 2.51 ;
 RECT 2.95 0.845 3.18 1.055 ;
 LAYER CO ;
 RECT 9.86 1.97 9.99 2.1 ;
 RECT 9.39 1.885 9.52 2.015 ;
 RECT 9.39 0.665 9.52 0.795 ;
 RECT 9.04 1.885 9.17 2.015 ;
 RECT 9.04 0.665 9.17 0.795 ;
 RECT 5.91 0.58 6.04 0.71 ;
 RECT 5.91 1.495 6.04 1.625 ;
 RECT 6.235 0.98 6.365 1.11 ;
 RECT 2.59 1.105 2.72 1.235 ;
 RECT 4.74 1.175 4.87 1.305 ;
 RECT 5 0.39 5.13 0.52 ;
 RECT 5 1.845 5.13 1.975 ;
 RECT 4.525 0.11 4.655 0.24 ;
 RECT 4.525 2.145 4.655 2.275 ;
 RECT 3.58 2.145 3.71 2.275 ;
 RECT 2.67 0.595 2.8 0.725 ;
 RECT 2.67 1.845 2.8 1.975 ;
 RECT 1.74 0.57 1.87 0.7 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 1.535 0.97 1.665 1.1 ;
 RECT 8.165 0.325 8.295 0.455 ;
 RECT 8.28 2.23 8.41 2.36 ;
 RECT 3 0.885 3.13 1.015 ;
 RECT 9.86 0.595 9.99 0.725 ;
 RECT 8.28 1.97 8.41 2.1 ;
 RECT 7.985 1.175 8.115 1.305 ;
 RECT 7.295 1.06 7.425 1.19 ;
 RECT 6.65 1.175 6.78 1.305 ;
 RECT 3.58 0.145 3.71 0.275 ;
 RECT 4.185 0.71 4.315 0.84 ;
 RECT 4.055 0.39 4.185 0.52 ;
 RECT 4.055 1.845 4.185 1.975 ;
 RECT 1.74 1.82 1.87 1.95 ;
 RECT 1.265 0.205 1.395 0.335 ;
 RECT 1.265 2.145 1.395 2.275 ;
 RECT 0.795 0.57 0.925 0.7 ;
 RECT 0.795 1.82 0.925 1.95 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 5.91 2.45 6.04 2.58 ;
 RECT 9.33 0.225 9.46 0.355 ;
 RECT 8.48 0.135 8.61 0.265 ;
 LAYER M1 ;
 RECT 3.985 0.385 5.2 0.525 ;
 RECT 0.79 1.745 0.93 1.815 ;
 RECT 0.79 1.955 0.93 2.02 ;
 RECT 0.79 1.815 1.94 1.955 ;
 RECT 3.985 1.84 5.2 1.98 ;
 RECT 8.16 0.255 8.3 0.54 ;
 RECT 8.755 0.36 8.895 0.54 ;
 RECT 8.16 0.54 8.895 0.68 ;
 RECT 8.755 0.22 9.53 0.36 ;
 RECT 0.79 0.705 0.93 0.775 ;
 RECT 1.735 0.705 1.875 0.77 ;
 RECT 1.735 0.5 1.875 0.565 ;
 RECT 0.79 0.5 0.93 0.565 ;
 RECT 0.79 0.565 1.875 0.705 ;
 RECT 2.3 1.705 3.835 1.845 ;
 RECT 3.695 1.68 3.835 1.705 ;
 RECT 2.3 1.845 2.805 1.915 ;
 RECT 2.665 0.525 2.805 0.66 ;
 RECT 2.3 0.66 2.805 0.8 ;
 RECT 2.665 1.915 2.805 2.045 ;
 RECT 2.3 0.8 2.44 1.705 ;
 RECT 6.23 1.15 6.37 1.18 ;
 RECT 6.185 0.95 6.415 1.15 ;
 RECT 5.34 1.68 5.485 1.97 ;
 RECT 5.34 1.97 5.48 2.135 ;
 RECT 3.695 1.54 5.485 1.68 ;
 RECT 6.185 0.94 7.14 0.95 ;
 RECT 6.23 0.81 7.14 0.94 ;
 RECT 5.34 2.135 7.14 2.275 ;
 RECT 7 0.95 7.14 2.135 ;
 RECT 5.905 0.65 6.045 1.685 ;
 RECT 7.59 0.65 7.73 1.17 ;
 RECT 5.905 0.51 7.73 0.65 ;
 RECT 7.975 1.1 8.12 1.17 ;
 RECT 7.59 1.17 8.12 1.31 ;
 RECT 7.975 1.31 8.12 1.41 ;
 END
END FADDX1

MACRO FADDX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.88 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.88 2.96 ;
 RECT 4.455 2.14 4.725 2.28 ;
 RECT 3.575 2.075 3.715 2.8 ;
 RECT 8.275 1.9 8.415 2.8 ;
 RECT 1.26 2.095 1.4 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 9.505 1.9 9.645 2.8 ;
 RECT 10.445 1.9 10.585 2.8 ;
 RECT 4.52 2.28 4.66 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.88 0.08 ;
 RECT 9.505 0.5 10.295 0.64 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 10.155 0.08 10.295 0.5 ;
 RECT 8.475 0.08 8.615 0.34 ;
 RECT 1.26 0.08 1.4 0.41 ;
 RECT 4.44 0.08 4.745 0.245 ;
 RECT 3.485 0.08 3.8 0.28 ;
 RECT 10.445 0.08 10.585 0.795 ;
 RECT 9.505 0.64 9.645 0.795 ;
 END
 END VSS

 PIN A
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.75 2.415 6.34 2.66 ;
 END
 ANTENNAGATEAREA 0.476 ;
 END A

 PIN B
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.015 0.365 2.155 0.965 ;
 RECT 2.015 0.225 3.085 0.365 ;
 RECT 5.34 0.36 5.48 0.665 ;
 RECT 7.88 0.82 8.41 0.96 ;
 RECT 7.295 1.615 8.41 1.755 ;
 RECT 7.28 1.05 7.435 1.195 ;
 RECT 1.27 0.965 2.155 1.105 ;
 RECT 1.27 1.105 1.715 1.505 ;
 RECT 1.27 0.93 1.715 0.965 ;
 RECT 2.945 0.365 3.085 0.665 ;
 RECT 7.88 0.36 8.02 0.82 ;
 RECT 5.34 0.22 8.02 0.36 ;
 RECT 8.27 0.96 8.41 1.615 ;
 RECT 7.295 1.195 7.435 1.615 ;
 RECT 7.295 0.985 7.435 1.05 ;
 RECT 2.945 0.85 3.195 1.02 ;
 RECT 2.945 0.665 5.48 0.85 ;
 END
 ANTENNAGATEAREA 0.476 ;
 END B

 PIN CI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.585 1.035 2.725 1.26 ;
 RECT 5.625 1.85 6.815 1.99 ;
 RECT 6.645 1.095 6.815 1.4 ;
 RECT 4.665 1.175 5.765 1.26 ;
 RECT 2.585 1.26 5.765 1.315 ;
 RECT 3.195 1.4 3.55 1.435 ;
 RECT 3.195 1.16 3.55 1.26 ;
 RECT 2.585 1.315 4.945 1.4 ;
 RECT 5.625 1.315 5.765 1.85 ;
 RECT 6.675 1.4 6.815 1.85 ;
 RECT 4.735 1.105 4.875 1.175 ;
 END
 ANTENNAGATEAREA 0.357 ;
 END CI

 PIN CO
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.905 0.78 10.18 0.92 ;
 RECT 9.975 1.43 10.115 2.495 ;
 RECT 9.575 1.155 10.115 1.43 ;
 RECT 9.975 0.92 10.115 1.155 ;
 END
 ANTENNADIFFAREA 0.592 ;
 END CO

 PIN S
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.56 2.035 9.175 2.405 ;
 RECT 9.035 0.595 9.175 2.035 ;
 END
 ANTENNADIFFAREA 0.608 ;
 END S

 OBS
 LAYER PO ;
 RECT 4.305 0.09 4.405 0.67 ;
 RECT 4.135 0.67 4.405 0.88 ;
 RECT 4.305 0.88 4.405 2.51 ;
 RECT 1.515 0.285 1.615 0.93 ;
 RECT 1.515 1.14 1.615 2.51 ;
 RECT 1.485 0.93 1.715 1.14 ;
 RECT 7.02 0.375 7.12 1.02 ;
 RECT 7.02 1.23 7.12 2.51 ;
 RECT 7.02 1.02 7.475 1.23 ;
 RECT 6.715 0.375 6.815 1.115 ;
 RECT 6.715 1.345 6.815 2.51 ;
 RECT 6.595 1.115 6.84 1.345 ;
 RECT 5.25 0.195 5.35 0.97 ;
 RECT 5.25 1.07 5.35 2.51 ;
 RECT 6.185 0.94 6.415 0.97 ;
 RECT 6.185 1.07 6.415 1.15 ;
 RECT 5.25 0.095 8.355 0.195 ;
 RECT 8.11 0.195 8.355 0.5 ;
 RECT 5.25 0.97 6.415 1.07 ;
 RECT 2.105 0.285 2.205 1.065 ;
 RECT 2.105 1.065 2.77 1.275 ;
 RECT 2.105 1.275 2.205 2.51 ;
 RECT 4.775 0.095 4.875 1.135 ;
 RECT 4.775 1.345 4.875 2.51 ;
 RECT 4.69 1.135 4.92 1.345 ;
 RECT 9.76 0.4 9.86 1.11 ;
 RECT 9.76 1.11 10.33 1.21 ;
 RECT 9.76 1.21 9.86 2.79 ;
 RECT 10.23 0.29 10.33 1.11 ;
 RECT 10.23 1.21 10.33 2.79 ;
 RECT 9.57 0.14 10.02 0.4 ;
 RECT 1.045 0.285 1.145 2.69 ;
 RECT 3.83 0.105 3.93 2.69 ;
 RECT 7.655 0.375 7.755 2.69 ;
 RECT 3.36 0.285 3.46 2.69 ;
 RECT 5.855 2.4 6.085 2.69 ;
 RECT 1.045 2.69 7.755 2.79 ;
 RECT 2.99 0.285 3.09 0.845 ;
 RECT 2.99 1.055 3.09 2.51 ;
 RECT 2.95 0.845 3.18 1.055 ;
 RECT 8.815 0.215 8.915 1.135 ;
 RECT 8.815 1.345 8.915 2.79 ;
 RECT 9.29 0.215 9.39 1.135 ;
 RECT 7.935 1.135 9.39 1.345 ;
 RECT 9.29 1.345 9.39 2.79 ;
 LAYER CO ;
 RECT 9.51 0.595 9.64 0.725 ;
 RECT 10.45 1.97 10.58 2.1 ;
 RECT 9.98 2.29 10.11 2.42 ;
 RECT 7.985 1.175 8.115 1.305 ;
 RECT 7.295 1.06 7.425 1.19 ;
 RECT 6.65 1.175 6.78 1.305 ;
 RECT 5.91 0.58 6.04 0.71 ;
 RECT 5.91 1.495 6.04 1.625 ;
 RECT 6.235 0.98 6.365 1.11 ;
 RECT 4.185 0.71 4.315 0.84 ;
 RECT 4.055 0.39 4.185 0.52 ;
 RECT 4.055 1.845 4.185 1.975 ;
 RECT 5 0.39 5.13 0.52 ;
 RECT 5 1.845 5.13 1.975 ;
 RECT 4.525 0.11 4.655 0.24 ;
 RECT 4.525 2.145 4.655 2.275 ;
 RECT 1.265 2.145 1.395 2.275 ;
 RECT 0.795 0.57 0.925 0.7 ;
 RECT 0.795 1.82 0.925 1.95 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 1.535 0.97 1.665 1.1 ;
 RECT 9.51 1.97 9.64 2.1 ;
 RECT 10.45 0.595 10.58 0.725 ;
 RECT 3.58 2.145 3.71 2.275 ;
 RECT 2.67 0.595 2.8 0.725 ;
 RECT 2.67 1.845 2.8 1.975 ;
 RECT 1.74 0.57 1.87 0.7 ;
 RECT 1.74 1.82 1.87 1.95 ;
 RECT 1.265 0.205 1.395 0.335 ;
 RECT 2.59 1.105 2.72 1.235 ;
 RECT 4.74 1.175 4.87 1.305 ;
 RECT 3.58 0.145 3.71 0.275 ;
 RECT 9.755 0.225 9.885 0.355 ;
 RECT 8.48 0.135 8.61 0.265 ;
 RECT 8.165 0.325 8.295 0.455 ;
 RECT 5.91 2.45 6.04 2.58 ;
 RECT 8.28 2.23 8.41 2.36 ;
 RECT 3 0.885 3.13 1.015 ;
 RECT 9.98 0.785 10.11 0.915 ;
 RECT 9.04 1.885 9.17 2.015 ;
 RECT 9.04 0.665 9.17 0.795 ;
 RECT 8.28 1.97 8.41 2.1 ;
 LAYER M1 ;
 RECT 3.985 0.385 5.2 0.525 ;
 RECT 0.79 1.745 0.93 1.815 ;
 RECT 0.79 1.955 0.93 2.02 ;
 RECT 0.79 1.815 1.94 1.955 ;
 RECT 3.985 1.84 5.2 1.98 ;
 RECT 8.755 0.36 8.895 0.54 ;
 RECT 8.16 0.54 8.895 0.68 ;
 RECT 8.16 0.255 8.3 0.54 ;
 RECT 8.755 0.22 9.96 0.36 ;
 RECT 5.905 0.65 6.045 1.685 ;
 RECT 5.905 0.51 7.73 0.65 ;
 RECT 7.59 0.65 7.73 1.17 ;
 RECT 7.975 1.1 8.12 1.17 ;
 RECT 7.975 1.31 8.12 1.41 ;
 RECT 7.59 1.17 8.12 1.31 ;
 RECT 0.79 0.705 0.93 0.775 ;
 RECT 1.735 0.705 1.875 0.77 ;
 RECT 0.79 0.5 0.93 0.565 ;
 RECT 1.735 0.5 1.875 0.565 ;
 RECT 0.79 0.565 1.875 0.705 ;
 RECT 2.3 1.705 3.835 1.845 ;
 RECT 3.695 1.68 3.835 1.705 ;
 RECT 2.3 1.845 2.805 1.915 ;
 RECT 2.665 0.525 2.805 0.66 ;
 RECT 2.3 0.66 2.805 0.8 ;
 RECT 2.665 1.915 2.805 2.045 ;
 RECT 2.3 0.8 2.44 1.705 ;
 RECT 6.23 1.15 6.37 1.18 ;
 RECT 6.185 0.95 6.415 1.15 ;
 RECT 3.695 1.54 5.485 1.68 ;
 RECT 5.34 1.68 5.485 1.97 ;
 RECT 5.34 1.97 5.48 2.135 ;
 RECT 6.185 0.94 7.14 0.95 ;
 RECT 6.23 0.81 7.14 0.94 ;
 RECT 5.34 2.135 7.14 2.275 ;
 RECT 7 0.95 7.14 2.135 ;
 END
END FADDX2

MACRO HADDX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 2.97 2.33 3.245 2.47 ;
 RECT 1.72 2.285 1.86 2.8 ;
 RECT 0.35 1.945 0.49 2.8 ;
 RECT 4.445 1.895 4.585 2.8 ;
 RECT 3.035 2.47 3.175 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 2.215 0.7 2.485 0.84 ;
 RECT 0.35 0.08 0.49 0.765 ;
 RECT 4.445 0.08 4.585 0.905 ;
 RECT 2.28 0.08 2.42 0.7 ;
 END
 END VSS

 PIN B0
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 1.425 1.275 1.725 ;
 END
 ANTENNAGATEAREA 0.151 ;
 END B0

 PIN A0
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.61 1.285 2.65 1.425 ;
 RECT 1.61 1.425 1.88 1.605 ;
 RECT 1.61 1.28 1.88 1.285 ;
 END
 ANTENNAGATEAREA 0.151 ;
 END A0

 PIN C1
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.515 0.8 4.01 1.12 ;
 RECT 3.87 1.12 4.01 2.12 ;
 RECT 3.87 0.635 4.01 0.8 ;
 END
 ANTENNADIFFAREA 0.526 ;
 END C1

 PIN SO
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.73 1.45 5.23 1.77 ;
 RECT 4.92 1.77 5.06 2.47 ;
 RECT 4.92 0.635 5.06 1.45 ;
 END
 ANTENNADIFFAREA 0.46 ;
 END SO

 OBS
 LAYER PO ;
 RECT 4.7 0.36 4.8 1.08 ;
 RECT 4.565 1.08 4.8 1.31 ;
 RECT 4.7 1.31 4.8 2.75 ;
 RECT 4.18 0.465 4.28 2.75 ;
 RECT 4.05 0.235 4.28 0.465 ;
 RECT 1.98 0.955 2.22 1.185 ;
 RECT 1.98 1.185 2.08 2.78 ;
 RECT 2.065 0.465 2.165 0.955 ;
 RECT 2.4 1.24 2.635 1.365 ;
 RECT 2.535 0.465 2.635 1.24 ;
 RECT 2.81 1.465 2.91 2.7 ;
 RECT 2.4 1.465 2.63 1.47 ;
 RECT 2.4 1.365 2.91 1.465 ;
 RECT 1.415 1.715 1.69 1.815 ;
 RECT 1.59 1.535 1.69 1.715 ;
 RECT 1.415 1.815 1.515 2.78 ;
 RECT 1.59 0.48 1.69 1.305 ;
 RECT 1.58 1.305 1.8 1.535 ;
 RECT 3.29 1.09 3.39 2.7 ;
 RECT 2.835 0.285 2.935 0.99 ;
 RECT 1.11 0.285 1.21 1.435 ;
 RECT 1.025 1.665 1.125 2.78 ;
 RECT 2.835 0.99 3.39 1.09 ;
 RECT 1.11 0.185 2.935 0.285 ;
 RECT 1.005 1.435 1.235 1.665 ;
 LAYER CO ;
 RECT 4.615 1.13 4.745 1.26 ;
 RECT 4.1 0.285 4.23 0.415 ;
 RECT 4.925 0.705 5.055 0.835 ;
 RECT 4.45 0.705 4.58 0.835 ;
 RECT 3.875 0.705 4.005 0.835 ;
 RECT 4.925 2.27 5.055 2.4 ;
 RECT 4.925 1.97 5.055 2.1 ;
 RECT 4.45 2.27 4.58 2.4 ;
 RECT 4.45 1.97 4.58 2.1 ;
 RECT 3.875 1.92 4.005 2.05 ;
 RECT 3.875 1.63 4.005 1.76 ;
 RECT 2.04 1.005 2.17 1.135 ;
 RECT 2.45 1.29 2.58 1.42 ;
 RECT 3.055 0.705 3.185 0.835 ;
 RECT 3.515 1.72 3.645 1.85 ;
 RECT 3.04 2.335 3.17 2.465 ;
 RECT 2.56 1.72 2.69 1.85 ;
 RECT 2.205 2.27 2.335 2.4 ;
 RECT 2.285 0.705 2.415 0.835 ;
 RECT 0.355 0.305 0.485 0.435 ;
 RECT 0.355 0.565 0.485 0.695 ;
 RECT 0.355 2.015 0.485 2.145 ;
 RECT 0.355 2.275 0.485 2.405 ;
 RECT 1.62 1.355 1.75 1.485 ;
 RECT 1.055 1.485 1.185 1.615 ;
 RECT 1.815 0.705 1.945 0.835 ;
 RECT 1.335 0.705 1.465 0.835 ;
 RECT 0.86 0.705 0.99 0.835 ;
 RECT 1.725 2.375 1.855 2.505 ;
 RECT 0.765 1.965 0.895 2.095 ;
 RECT 0.765 2.27 0.895 2.4 ;
 LAYER M1 ;
 RECT 3.51 1.725 3.65 1.9 ;
 RECT 2.555 1.585 3.65 1.725 ;
 RECT 3.05 0.42 3.19 1 ;
 RECT 3.05 1.14 3.19 1.585 ;
 RECT 2.555 1.725 2.695 1.9 ;
 RECT 1.99 1 3.19 1.14 ;
 RECT 3.05 0.28 4.305 0.42 ;
 RECT 0.76 2.095 3.685 2.145 ;
 RECT 2.2 2.145 3.685 2.19 ;
 RECT 3.545 2.19 3.685 2.49 ;
 RECT 1.435 2.05 3.685 2.095 ;
 RECT 4.165 1.26 4.305 2.49 ;
 RECT 3.545 2.49 4.305 2.63 ;
 RECT 1.435 2.005 2.34 2.05 ;
 RECT 2.2 2.19 2.34 2.47 ;
 RECT 0.76 2.015 0.9 2.095 ;
 RECT 0.76 2.235 0.9 2.47 ;
 RECT 0.715 1.235 0.855 1.875 ;
 RECT 0.715 1.875 0.9 2.015 ;
 RECT 1.33 0.84 1.47 1.095 ;
 RECT 1.435 2 1.575 2.005 ;
 RECT 0.76 2.145 1.575 2.235 ;
 RECT 0.715 1.095 1.47 1.235 ;
 RECT 1.265 0.7 1.535 0.84 ;
 RECT 4.615 1.06 4.755 1.12 ;
 RECT 4.165 1.12 4.755 1.26 ;
 RECT 4.615 1.26 4.755 1.31 ;
 RECT 1.81 0.56 1.95 0.7 ;
 RECT 0.855 0.56 0.995 0.7 ;
 RECT 0.855 0.42 1.95 0.56 ;
 RECT 1.745 0.7 2.01 0.84 ;
 RECT 0.81 0.7 1.06 0.84 ;
 END
END HADDX1

MACRO HADDX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.4 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.4 2.96 ;
 RECT 2.97 2.33 3.245 2.47 ;
 RECT 3.805 2.235 4.075 2.375 ;
 RECT 1.72 2.285 1.86 2.8 ;
 RECT 0.35 1.945 0.49 2.8 ;
 RECT 4.935 1.895 5.075 2.8 ;
 RECT 5.88 1.925 6.02 2.8 ;
 RECT 3.035 2.47 3.175 2.8 ;
 RECT 3.87 2.375 4.01 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.4 0.08 ;
 RECT 2.215 0.7 2.485 0.84 ;
 RECT 0.35 0.08 0.49 0.765 ;
 RECT 4.935 0.08 5.075 0.855 ;
 RECT 3.795 0.08 3.935 0.865 ;
 RECT 5.88 0.08 6.02 0.855 ;
 RECT 2.28 0.08 2.42 0.7 ;
 END
 END VSS

 PIN B0
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.99 1.425 1.275 1.725 ;
 END
 ANTENNAGATEAREA 0.151 ;
 END B0

 PIN A0
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.61 1.285 2.65 1.425 ;
 RECT 1.61 1.425 1.88 1.605 ;
 RECT 1.61 1.28 1.88 1.285 ;
 END
 ANTENNAGATEAREA 0.151 ;
 END A0

 PIN C1
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.005 1.47 4.5 1.79 ;
 RECT 4.36 0.585 4.5 1.47 ;
 END
 ANTENNADIFFAREA 0.654 ;
 END C1

 PIN SO
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.41 1.77 5.55 2.47 ;
 RECT 5.41 1.45 5.92 1.77 ;
 RECT 5.41 0.585 5.55 1.45 ;
 END
 ANTENNADIFFAREA 0.57 ;
 END SO

 OBS
 LAYER PO ;
 RECT 5.055 1.08 5.29 1.175 ;
 RECT 5.055 1.175 5.765 1.275 ;
 RECT 5.055 1.275 5.29 1.31 ;
 RECT 5.665 0.355 5.765 1.175 ;
 RECT 5.665 1.275 5.765 2.75 ;
 RECT 5.19 0.345 5.29 1.08 ;
 RECT 5.19 1.31 5.29 2.75 ;
 RECT 4.67 0.44 4.77 1.165 ;
 RECT 4.67 1.265 4.77 2.75 ;
 RECT 4.14 1.165 4.77 1.265 ;
 RECT 4.14 0.35 4.24 1.165 ;
 RECT 4.14 1.265 4.24 2.75 ;
 RECT 4.54 0.21 4.77 0.44 ;
 RECT 1.98 0.955 2.215 1.185 ;
 RECT 1.98 1.185 2.08 2.73 ;
 RECT 2.065 0.465 2.165 0.955 ;
 RECT 2.4 1.24 2.635 1.365 ;
 RECT 2.535 0.465 2.635 1.24 ;
 RECT 2.81 1.465 2.91 2.7 ;
 RECT 2.4 1.465 2.63 1.47 ;
 RECT 2.4 1.365 2.91 1.465 ;
 RECT 1.415 1.655 1.68 1.755 ;
 RECT 1.58 1.535 1.68 1.655 ;
 RECT 1.415 1.755 1.515 2.725 ;
 RECT 1.59 0.465 1.69 1.305 ;
 RECT 1.58 1.305 1.8 1.535 ;
 RECT 3.29 1.09 3.39 2.7 ;
 RECT 2.835 0.285 2.935 0.99 ;
 RECT 1.11 0.285 1.21 1.435 ;
 RECT 1.025 1.665 1.125 2.725 ;
 RECT 2.835 0.99 3.39 1.09 ;
 RECT 1.11 0.185 2.935 0.285 ;
 RECT 1.005 1.435 1.235 1.665 ;
 LAYER CO ;
 RECT 5.885 1.99 6.015 2.12 ;
 RECT 5.885 0.655 6.015 0.785 ;
 RECT 5.885 2.27 6.015 2.4 ;
 RECT 3.875 2.24 4.005 2.37 ;
 RECT 3.8 0.665 3.93 0.795 ;
 RECT 5.105 1.13 5.235 1.26 ;
 RECT 4.59 0.26 4.72 0.39 ;
 RECT 5.415 0.655 5.545 0.785 ;
 RECT 4.94 0.655 5.07 0.785 ;
 RECT 4.365 0.655 4.495 0.785 ;
 RECT 5.415 2.27 5.545 2.4 ;
 RECT 5.415 1.97 5.545 2.1 ;
 RECT 4.94 2.27 5.07 2.4 ;
 RECT 4.94 1.97 5.07 2.1 ;
 RECT 4.365 1.58 4.495 1.71 ;
 RECT 2.035 1.005 2.165 1.135 ;
 RECT 2.45 1.29 2.58 1.42 ;
 RECT 3.055 0.705 3.185 0.835 ;
 RECT 3.515 1.59 3.645 1.72 ;
 RECT 3.04 2.335 3.17 2.465 ;
 RECT 2.56 1.655 2.69 1.785 ;
 RECT 2.205 2.27 2.335 2.4 ;
 RECT 2.285 0.705 2.415 0.835 ;
 RECT 0.355 0.305 0.485 0.435 ;
 RECT 0.355 0.565 0.485 0.695 ;
 RECT 0.355 2.015 0.485 2.145 ;
 RECT 0.355 2.275 0.485 2.405 ;
 RECT 1.62 1.355 1.75 1.485 ;
 RECT 1.055 1.485 1.185 1.615 ;
 RECT 1.815 0.705 1.945 0.835 ;
 RECT 1.335 0.705 1.465 0.835 ;
 RECT 0.86 0.705 0.99 0.835 ;
 RECT 1.725 2.335 1.855 2.465 ;
 RECT 0.765 1.965 0.895 2.095 ;
 RECT 0.765 2.27 0.895 2.4 ;
 LAYER M1 ;
 RECT 0.855 0.56 0.995 0.7 ;
 RECT 1.81 0.56 1.95 0.7 ;
 RECT 0.855 0.42 1.95 0.56 ;
 RECT 1.745 0.7 2.01 0.84 ;
 RECT 0.81 0.7 1.06 0.84 ;
 RECT 3.05 0.635 3.19 1 ;
 RECT 3.05 1.195 3.19 1.585 ;
 RECT 1.985 1 3.19 1.055 ;
 RECT 2.555 1.725 2.695 1.86 ;
 RECT 2.555 1.585 3.705 1.725 ;
 RECT 4.08 0.395 4.22 1.055 ;
 RECT 1.985 1.055 4.22 1.14 ;
 RECT 3.025 1.14 4.22 1.195 ;
 RECT 4.08 0.255 4.79 0.395 ;
 RECT 1.435 2.025 4.795 2.095 ;
 RECT 4.655 1.26 4.795 1.955 ;
 RECT 3.045 1.955 4.795 2.025 ;
 RECT 0.76 2.095 3.185 2.145 ;
 RECT 2.2 2.145 3.185 2.165 ;
 RECT 1.435 2.005 2.34 2.025 ;
 RECT 2.2 2.165 2.34 2.47 ;
 RECT 0.76 2.015 0.9 2.095 ;
 RECT 0.76 2.235 0.9 2.47 ;
 RECT 0.71 1.235 0.85 1.875 ;
 RECT 0.71 1.875 0.9 2.015 ;
 RECT 1.33 0.84 1.47 1.095 ;
 RECT 1.435 2 1.575 2.005 ;
 RECT 0.76 2.145 1.575 2.235 ;
 RECT 0.71 1.095 1.47 1.235 ;
 RECT 1.265 0.7 1.535 0.84 ;
 RECT 5.105 1.06 5.245 1.12 ;
 RECT 4.655 1.12 5.245 1.26 ;
 RECT 5.105 1.26 5.245 1.31 ;
 END
END HADDX2

MACRO LARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.96 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.975 1.16 1.275 1.425 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.965 1.155 2.315 1.45 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.32 2.045 7.705 2.335 ;
 RECT 7.435 2.335 7.575 2.555 ;
 RECT 7.435 0.86 7.575 2.045 ;
 RECT 7.38 0.72 7.61 0.86 ;
 END
 ANTENNADIFFAREA 0.505 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.96 2.96 ;
 RECT 7.915 1.455 8.055 2.8 ;
 RECT 7.03 1.905 7.17 2.8 ;
 RECT 5.715 1.9 5.855 2.8 ;
 RECT 2.66 2.605 2.89 2.8 ;
 RECT 1.84 2.63 2.07 2.8 ;
 RECT 0.93 1.88 1.07 2.8 ;
 RECT 0.425 1.755 0.565 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.96 0.08 ;
 RECT 3.32 0.08 3.46 0.83 ;
 RECT 0.34 0.08 0.48 0.81 ;
 RECT 0.93 0.08 1.07 1.015 ;
 RECT 2.07 0.08 2.21 1.015 ;
 RECT 5.19 0.08 5.42 0.29 ;
 RECT 6.715 0.08 6.855 0.74 ;
 RECT 7.86 0.08 8.09 0.275 ;
 RECT 3.32 0.83 3.575 0.97 ;
 RECT 6.51 0.74 6.855 0.88 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.26 2.065 8.695 2.4 ;
 RECT 8.385 2.4 8.525 2.57 ;
 RECT 8.385 0.415 8.525 2.065 ;
 END
 ANTENNADIFFAREA 0.472 ;
 END QN

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.66 0.46 5.875 0.6 ;
 RECT 5.56 0.345 5.875 0.46 ;
 RECT 3.66 0.235 3.8 0.46 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 OBS
 LAYER PO ;
 RECT 1.185 0.615 1.285 1.175 ;
 RECT 1.03 1.175 1.285 1.405 ;
 RECT 1.185 1.405 1.285 2.37 ;
 RECT 2.33 0.595 2.43 1.18 ;
 RECT 2.01 1.18 2.43 1.41 ;
 RECT 2.125 1.41 2.225 2.375 ;
 RECT 5.97 0.615 6.07 1.14 ;
 RECT 5.97 1.14 6.47 1.37 ;
 RECT 5.97 1.37 6.07 2.385 ;
 RECT 6.815 0.525 6.915 2.585 ;
 RECT 5.035 2.455 5.265 2.585 ;
 RECT 5.035 2.585 6.915 2.685 ;
 RECT 5.5 0.335 5.79 0.565 ;
 RECT 5.5 0.565 5.6 2.385 ;
 RECT 3.175 0.595 3.275 1.095 ;
 RECT 2.97 1.195 3.07 1.58 ;
 RECT 2.97 1.095 3.275 1.195 ;
 RECT 4.5 0.61 4.6 1.55 ;
 RECT 3.815 1.55 4.6 1.65 ;
 RECT 2.8 1.58 3.07 1.81 ;
 RECT 3.815 1.65 3.915 2.485 ;
 RECT 2.97 1.81 3.07 2.485 ;
 RECT 2.97 2.485 3.915 2.585 ;
 RECT 8.17 0.245 8.27 1.02 ;
 RECT 8.005 1.02 8.27 1.255 ;
 RECT 8.17 1.255 8.27 2.755 ;
 RECT 3.615 0.235 3.845 0.315 ;
 RECT 3.615 0.415 3.845 0.465 ;
 RECT 1.485 0.315 3.845 0.415 ;
 RECT 1.655 1.405 1.755 2.365 ;
 RECT 1.485 1.305 1.755 1.405 ;
 RECT 1.485 0.415 1.585 1.305 ;
 RECT 3.535 1.22 3.755 1.37 ;
 RECT 3.535 1.12 4.13 1.22 ;
 RECT 4.03 0.43 4.13 1.12 ;
 RECT 4.03 0.33 5.07 0.43 ;
 RECT 4.97 0.43 5.07 1.835 ;
 RECT 4.285 1.835 5.07 1.935 ;
 RECT 4.285 1.935 4.385 2.48 ;
 RECT 6.285 0.255 6.515 0.42 ;
 RECT 7.69 0.255 7.79 2.755 ;
 RECT 6.285 0.155 7.79 0.255 ;
 LAYER CO ;
 RECT 1.705 0.835 1.835 0.965 ;
 RECT 7.035 0.745 7.165 0.875 ;
 RECT 3.665 0.285 3.795 0.415 ;
 RECT 5.085 2.505 5.215 2.635 ;
 RECT 3.395 0.835 3.525 0.965 ;
 RECT 6.335 0.24 6.465 0.37 ;
 RECT 6.56 0.745 6.69 0.875 ;
 RECT 7.91 0.11 8.04 0.24 ;
 RECT 8.39 0.465 8.52 0.595 ;
 RECT 8.055 1.07 8.185 1.2 ;
 RECT 8.39 0.725 8.52 0.855 ;
 RECT 7.92 2.115 8.05 2.245 ;
 RECT 8.39 1.595 8.52 1.725 ;
 RECT 7.92 2.375 8.05 2.505 ;
 RECT 8.39 1.855 8.52 1.985 ;
 RECT 8.39 2.115 8.52 2.245 ;
 RECT 7.92 1.855 8.05 1.985 ;
 RECT 8.39 2.375 8.52 2.505 ;
 RECT 7.92 2.115 8.05 2.245 ;
 RECT 7.92 2.375 8.05 2.505 ;
 RECT 7.43 0.725 7.56 0.855 ;
 RECT 2.075 0.835 2.205 0.965 ;
 RECT 3.575 1.19 3.705 1.32 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 4.72 0.835 4.85 0.965 ;
 RECT 4.505 2.125 4.635 2.255 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 3.78 0.835 3.91 0.965 ;
 RECT 3.565 2.105 3.695 2.235 ;
 RECT 4.035 2.125 4.165 2.255 ;
 RECT 2.71 2.61 2.84 2.74 ;
 RECT 1.89 2.64 2.02 2.77 ;
 RECT 2.06 1.23 2.19 1.36 ;
 RECT 2.86 1.63 2.99 1.76 ;
 RECT 2.92 0.835 3.05 0.965 ;
 RECT 3.19 2.035 3.32 2.165 ;
 RECT 2.55 0.835 2.68 0.965 ;
 RECT 2.345 2.005 2.475 2.135 ;
 RECT 1.405 1.995 1.535 2.125 ;
 RECT 0.935 0.835 1.065 0.965 ;
 RECT 0.935 1.995 1.065 2.125 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 1.08 1.225 1.21 1.355 ;
 RECT 6.29 1.19 6.42 1.32 ;
 RECT 7.92 1.595 8.05 1.725 ;
 RECT 7.44 1.595 7.57 1.725 ;
 RECT 7.44 1.855 7.57 1.985 ;
 RECT 7.44 2.115 7.57 2.245 ;
 RECT 7.44 2.375 7.57 2.505 ;
 RECT 7.44 1.595 7.57 1.725 ;
 RECT 7.44 1.855 7.57 1.985 ;
 RECT 7.44 2.115 7.57 2.245 ;
 RECT 7.44 2.375 7.57 2.505 ;
 RECT 6.565 1.99 6.695 2.12 ;
 RECT 7.035 1.975 7.165 2.105 ;
 RECT 6.19 1.99 6.32 2.12 ;
 RECT 5.25 1.99 5.38 2.12 ;
 RECT 5.615 0.385 5.745 0.515 ;
 RECT 5.72 1.99 5.85 2.12 ;
 RECT 6.19 0.835 6.32 0.965 ;
 RECT 5.24 0.125 5.37 0.255 ;
 LAYER M1 ;
 RECT 4.22 0.77 4.39 1.02 ;
 RECT 4.22 1.02 4.36 1.775 ;
 RECT 4.03 1.775 4.36 1.915 ;
 RECT 4.03 1.915 4.17 2.5 ;
 RECT 4.03 2.5 5.265 2.64 ;
 RECT 2.915 0.775 3.055 1.185 ;
 RECT 3.185 1.325 3.325 2.03 ;
 RECT 3.185 2.17 3.325 2.185 ;
 RECT 3.1 2.03 3.37 2.17 ;
 RECT 2.915 1.185 3.755 1.325 ;
 RECT 2.545 0.785 2.685 1.625 ;
 RECT 2.34 1.625 3.045 1.765 ;
 RECT 2.34 1.765 2.48 2 ;
 RECT 2.295 2 2.525 2.14 ;
 RECT 2.34 2.14 2.48 2.175 ;
 RECT 1.555 0.97 1.695 1.99 ;
 RECT 1.4 2.13 1.54 2.325 ;
 RECT 1.555 0.83 1.905 0.97 ;
 RECT 1.31 1.99 1.695 2.13 ;
 RECT 3.73 0.83 4.08 0.97 ;
 RECT 3.94 0.97 4.08 1.465 ;
 RECT 3.56 1.465 4.08 1.605 ;
 RECT 3.56 1.605 3.7 2.325 ;
 RECT 1.4 2.325 3.7 2.465 ;
 RECT 6.56 1.325 6.7 1.985 ;
 RECT 7.03 0.575 7.17 1.185 ;
 RECT 6.19 1.185 7.17 1.325 ;
 RECT 6.515 1.985 6.745 2.125 ;
 RECT 7.03 0.435 8.025 0.575 ;
 RECT 7.885 0.575 8.025 1.065 ;
 RECT 7.885 1.065 8.235 1.205 ;
 RECT 5.2 1.985 5.43 2.125 ;
 RECT 5.245 1.69 5.385 1.985 ;
 RECT 6.23 0.375 6.37 0.83 ;
 RECT 6.14 1.985 6.37 2.125 ;
 RECT 6.185 1.69 6.325 1.985 ;
 RECT 5.24 1.55 6.325 1.69 ;
 RECT 5.715 1.3 5.855 1.55 ;
 RECT 4.5 1.16 5.855 1.3 ;
 RECT 5.715 0.97 5.855 1.16 ;
 RECT 5.715 0.83 6.37 0.97 ;
 RECT 4.41 2.12 4.695 2.26 ;
 RECT 4.715 0.78 4.855 1.16 ;
 RECT 4.5 1.3 4.64 2.12 ;
 RECT 6.23 0.235 6.515 0.375 ;
 END
END LARX1

MACRO LARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.24 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.995 1.17 1.275 1.425 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.095 1.16 2.36 1.45 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.32 2.08 7.705 2.37 ;
 RECT 7.435 2.37 7.575 2.61 ;
 RECT 7.38 0.72 7.61 0.86 ;
 RECT 7.435 1.215 8.525 1.355 ;
 RECT 8.3 0.72 8.59 0.86 ;
 RECT 7.435 1.355 7.575 2.08 ;
 RECT 7.435 0.86 7.575 1.215 ;
 RECT 8.385 1.355 8.525 2.58 ;
 RECT 8.385 0.86 8.525 1.215 ;
 END
 ANTENNADIFFAREA 0.952 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.24 2.96 ;
 RECT 7.915 1.555 8.055 2.8 ;
 RECT 7.03 1.905 7.17 2.8 ;
 RECT 5.715 1.9 5.855 2.8 ;
 RECT 2.66 2.605 2.89 2.8 ;
 RECT 1.84 2.63 2.07 2.8 ;
 RECT 0.93 1.88 1.07 2.8 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 9.265 1.555 9.405 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.24 0.08 ;
 RECT 0.34 0.08 0.48 0.81 ;
 RECT 0.93 0.08 1.07 1.015 ;
 RECT 2.07 0.08 2.21 1.015 ;
 RECT 3.32 0.08 3.46 0.83 ;
 RECT 5.19 0.08 5.42 0.29 ;
 RECT 6.715 0.08 6.855 0.74 ;
 RECT 7.86 0.08 8.09 0.275 ;
 RECT 3.32 0.83 3.575 0.97 ;
 RECT 6.51 0.74 6.855 0.88 ;
 RECT 9.195 0.08 9.465 0.265 ;
 END
 END VSS

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.66 0.46 5.795 0.6 ;
 RECT 5.56 0.345 5.795 0.46 ;
 RECT 3.66 0.235 3.8 0.46 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.64 2.055 10 2.39 ;
 RECT 9.735 2.39 9.875 2.635 ;
 RECT 8.785 1.265 9.875 1.405 ;
 RECT 8.73 0.72 8.985 0.86 ;
 RECT 9.735 1.405 9.875 2.055 ;
 RECT 9.735 0.335 9.875 1.265 ;
 RECT 8.785 1.405 8.925 2.61 ;
 RECT 8.785 0.86 8.925 1.265 ;
 END
 ANTENNADIFFAREA 0.957 ;
 END QN

 OBS
 LAYER PO ;
 RECT 1.185 0.615 1.285 1.175 ;
 RECT 1.03 1.175 1.285 1.405 ;
 RECT 1.185 1.405 1.285 2.37 ;
 RECT 2.33 0.595 2.43 1.18 ;
 RECT 2.095 1.18 2.43 1.41 ;
 RECT 2.125 1.41 2.225 2.375 ;
 RECT 5.97 0.615 6.07 1.14 ;
 RECT 5.97 1.14 6.47 1.37 ;
 RECT 5.97 1.37 6.07 2.385 ;
 RECT 6.815 0.525 6.915 2.585 ;
 RECT 5.035 2.455 5.265 2.585 ;
 RECT 5.035 2.585 6.915 2.685 ;
 RECT 3.175 0.595 3.275 1.095 ;
 RECT 2.97 1.195 3.07 1.58 ;
 RECT 2.97 1.095 3.275 1.195 ;
 RECT 4.5 0.61 4.6 1.55 ;
 RECT 3.815 1.55 4.6 1.65 ;
 RECT 2.8 1.58 3.07 1.81 ;
 RECT 3.815 1.65 3.915 2.485 ;
 RECT 2.97 1.81 3.07 2.485 ;
 RECT 2.97 2.485 3.915 2.585 ;
 RECT 3.615 0.235 3.845 0.315 ;
 RECT 3.615 0.415 3.845 0.465 ;
 RECT 1.485 0.315 3.845 0.415 ;
 RECT 1.655 1.405 1.755 2.365 ;
 RECT 1.485 1.305 1.755 1.405 ;
 RECT 1.485 0.415 1.585 1.305 ;
 RECT 3.535 1.22 3.755 1.37 ;
 RECT 3.535 1.12 4.13 1.22 ;
 RECT 4.03 0.43 4.13 1.12 ;
 RECT 4.03 0.33 5.07 0.43 ;
 RECT 4.97 0.43 5.07 1.835 ;
 RECT 4.285 1.835 5.07 1.935 ;
 RECT 4.285 1.935 4.385 2.48 ;
 RECT 9.04 0.22 9.14 1.055 ;
 RECT 8.54 0.22 8.77 0.405 ;
 RECT 9.04 1.155 9.14 2.765 ;
 RECT 9.52 0.245 9.62 1.055 ;
 RECT 9.52 1.155 9.62 2.765 ;
 RECT 8.54 0.12 9.14 0.22 ;
 RECT 9.04 1.055 9.62 1.155 ;
 RECT 8.17 0.14 8.27 1.025 ;
 RECT 8.17 1.125 8.27 2.765 ;
 RECT 7.69 0.255 7.79 1.025 ;
 RECT 7.69 1.125 7.79 2.765 ;
 RECT 6.285 0.255 6.515 0.42 ;
 RECT 7.69 1.025 8.27 1.125 ;
 RECT 6.285 0.155 7.79 0.255 ;
 RECT 5.5 0.375 5.79 0.585 ;
 RECT 5.5 0.585 5.6 2.385 ;
 LAYER CO ;
 RECT 7.91 0.11 8.04 0.24 ;
 RECT 8.39 0.725 8.52 0.855 ;
 RECT 9.74 2.385 9.87 2.515 ;
 RECT 8.79 2.385 8.92 2.515 ;
 RECT 9.27 1.605 9.4 1.735 ;
 RECT 9.74 0.725 9.87 0.855 ;
 RECT 8.39 1.865 8.52 1.995 ;
 RECT 8.39 2.125 8.52 2.255 ;
 RECT 7.92 1.865 8.05 1.995 ;
 RECT 8.39 2.385 8.52 2.515 ;
 RECT 7.92 2.125 8.05 2.255 ;
 RECT 7.92 2.385 8.05 2.515 ;
 RECT 7.43 0.725 7.56 0.855 ;
 RECT 2.075 0.835 2.205 0.965 ;
 RECT 3.575 1.19 3.705 1.32 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 4.72 0.835 4.85 0.965 ;
 RECT 4.505 2.125 4.635 2.255 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 3.78 0.835 3.91 0.965 ;
 RECT 3.565 2.105 3.695 2.235 ;
 RECT 4.035 2.125 4.165 2.255 ;
 RECT 2.71 2.61 2.84 2.74 ;
 RECT 1.89 2.64 2.02 2.77 ;
 RECT 2.145 1.23 2.275 1.36 ;
 RECT 2.86 1.63 2.99 1.76 ;
 RECT 2.92 0.835 3.05 0.965 ;
 RECT 3.19 2.035 3.32 2.165 ;
 RECT 2.55 0.835 2.68 0.965 ;
 RECT 2.345 2.005 2.475 2.135 ;
 RECT 1.405 1.995 1.535 2.125 ;
 RECT 0.935 0.835 1.065 0.965 ;
 RECT 5.61 0.415 5.74 0.545 ;
 RECT 7.92 2.125 8.05 2.255 ;
 RECT 9.27 2.125 9.4 2.255 ;
 RECT 9.27 2.385 9.4 2.515 ;
 RECT 8.79 0.725 8.92 0.855 ;
 RECT 9.74 1.605 9.87 1.735 ;
 RECT 9.74 1.865 9.87 1.995 ;
 RECT 9.74 2.125 9.87 2.255 ;
 RECT 9.27 1.865 9.4 1.995 ;
 RECT 7.035 0.745 7.165 0.875 ;
 RECT 3.665 0.285 3.795 0.415 ;
 RECT 5.085 2.505 5.215 2.635 ;
 RECT 3.395 0.835 3.525 0.965 ;
 RECT 6.335 0.24 6.465 0.37 ;
 RECT 0.935 1.995 1.065 2.125 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 8.39 1.605 8.52 1.735 ;
 RECT 7.92 2.385 8.05 2.515 ;
 RECT 7.92 1.605 8.05 1.735 ;
 RECT 7.44 1.865 7.57 1.995 ;
 RECT 1.08 1.225 1.21 1.355 ;
 RECT 6.29 1.19 6.42 1.32 ;
 RECT 7.44 1.605 7.57 1.735 ;
 RECT 7.44 1.865 7.57 1.995 ;
 RECT 7.44 1.605 7.57 1.735 ;
 RECT 6.565 1.99 6.695 2.12 ;
 RECT 7.035 1.975 7.165 2.105 ;
 RECT 6.19 1.99 6.32 2.12 ;
 RECT 5.25 1.99 5.38 2.12 ;
 RECT 5.72 1.99 5.85 2.12 ;
 RECT 6.19 0.835 6.32 0.965 ;
 RECT 5.24 0.125 5.37 0.255 ;
 RECT 1.705 0.835 1.835 0.965 ;
 RECT 9.74 0.465 9.87 0.595 ;
 RECT 8.59 0.225 8.72 0.355 ;
 RECT 9.26 0.11 9.39 0.24 ;
 RECT 7.44 1.605 7.57 1.735 ;
 RECT 7.44 1.865 7.57 1.995 ;
 RECT 7.44 2.125 7.57 2.255 ;
 RECT 8.39 1.605 8.52 1.735 ;
 RECT 8.39 1.865 8.52 1.995 ;
 RECT 8.39 2.125 8.52 2.255 ;
 RECT 7.92 1.865 8.05 1.995 ;
 RECT 8.79 1.605 8.92 1.735 ;
 RECT 8.79 1.865 8.92 1.995 ;
 RECT 8.79 2.125 8.92 2.255 ;
 RECT 7.44 2.125 7.57 2.255 ;
 RECT 7.44 2.385 7.57 2.515 ;
 RECT 7.44 2.125 7.57 2.255 ;
 RECT 7.44 2.385 7.57 2.515 ;
 RECT 8.39 2.385 8.52 2.515 ;
 RECT 7.44 2.385 7.57 2.515 ;
 RECT 7.92 2.125 8.05 2.255 ;
 RECT 7.92 1.605 8.05 1.735 ;
 RECT 8.39 0.725 8.52 0.855 ;
 RECT 7.92 2.385 8.05 2.515 ;
 RECT 7.43 0.725 7.56 0.855 ;
 RECT 6.56 0.745 6.69 0.875 ;
 LAYER M1 ;
 RECT 4.22 0.77 4.39 1.02 ;
 RECT 4.22 1.02 4.36 1.775 ;
 RECT 4.03 1.775 4.36 1.915 ;
 RECT 4.03 1.915 4.17 2.5 ;
 RECT 4.03 2.5 5.265 2.64 ;
 RECT 2.915 0.775 3.055 1.185 ;
 RECT 3.185 1.325 3.325 2.03 ;
 RECT 3.185 2.17 3.325 2.185 ;
 RECT 3.1 2.03 3.37 2.17 ;
 RECT 2.915 1.185 3.755 1.325 ;
 RECT 2.545 0.785 2.685 1.625 ;
 RECT 2.34 1.625 3.045 1.765 ;
 RECT 2.34 1.765 2.48 2 ;
 RECT 2.295 2 2.525 2.14 ;
 RECT 2.34 2.14 2.48 2.175 ;
 RECT 1.7 0.785 1.84 1.99 ;
 RECT 1.4 2.13 1.54 2.325 ;
 RECT 1.31 1.99 1.84 2.13 ;
 RECT 3.73 0.83 4.08 0.97 ;
 RECT 3.94 0.97 4.08 1.465 ;
 RECT 3.56 1.465 4.08 1.605 ;
 RECT 3.56 1.605 3.7 2.325 ;
 RECT 1.4 2.325 3.7 2.465 ;
 RECT 7.03 0.575 7.17 1.185 ;
 RECT 6.19 1.185 7.17 1.325 ;
 RECT 6.515 1.985 6.745 2.125 ;
 RECT 6.56 1.325 6.7 1.985 ;
 RECT 8.465 0.36 8.605 0.435 ;
 RECT 7.03 0.435 8.605 0.575 ;
 RECT 8.465 0.22 8.88 0.36 ;
 RECT 5.2 1.985 5.43 2.125 ;
 RECT 5.245 1.69 5.385 1.985 ;
 RECT 6.23 0.375 6.37 0.83 ;
 RECT 6.14 1.985 6.37 2.125 ;
 RECT 6.185 1.69 6.325 1.985 ;
 RECT 5.24 1.55 6.325 1.69 ;
 RECT 5.715 1.3 5.855 1.55 ;
 RECT 4.5 1.16 5.855 1.3 ;
 RECT 5.715 0.97 5.855 1.16 ;
 RECT 5.715 0.83 6.37 0.97 ;
 RECT 4.41 2.12 4.695 2.26 ;
 RECT 4.715 0.78 4.855 1.16 ;
 RECT 4.5 1.3 4.64 2.12 ;
 RECT 6.23 0.235 6.515 0.375 ;
 END
END LARX2

MACRO LASRNX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.96 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.97 1.155 1.275 1.425 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.09 1.155 2.395 1.465 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.005 1.105 7.35 1.44 ;
 END
 ANTENNAGATEAREA 0.06 ;
 END SETB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.96 2.96 ;
 RECT 1.84 2.63 2.07 2.8 ;
 RECT 2.66 2.605 2.89 2.8 ;
 RECT 7.03 1.905 7.17 2.8 ;
 RECT 5.715 1.9 5.855 2.8 ;
 RECT 0.93 1.88 1.07 2.8 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 7.88 1.495 8.02 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.96 0.08 ;
 RECT 3.32 0.08 3.46 0.83 ;
 RECT 0.34 0.08 0.48 0.825 ;
 RECT 0.93 0.08 1.07 1.015 ;
 RECT 2.07 0.08 2.21 1.015 ;
 RECT 5.19 0.08 5.42 0.305 ;
 RECT 6.715 0.08 6.855 0.735 ;
 RECT 7.88 0.08 8.02 0.92 ;
 RECT 3.32 0.83 3.575 0.97 ;
 RECT 6.51 0.735 6.855 0.88 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.31 2.105 8.635 2.395 ;
 RECT 8.35 2.395 8.49 2.61 ;
 RECT 8.35 0.4 8.49 2.105 ;
 END
 ANTENNADIFFAREA 0.472 ;
 END QN

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.66 0.235 3.8 0.46 ;
 RECT 3.66 0.46 5.92 0.6 ;
 RECT 5.56 0.6 5.92 0.64 ;
 RECT 5.56 0.325 5.92 0.46 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 OBS
 LAYER PO ;
 RECT 1.185 0.615 1.285 1.175 ;
 RECT 1.03 1.175 1.285 1.405 ;
 RECT 1.185 1.405 1.285 2.37 ;
 RECT 2.33 0.595 2.43 1.18 ;
 RECT 2.125 1.18 2.43 1.41 ;
 RECT 2.125 1.41 2.225 2.375 ;
 RECT 5.97 0.615 6.07 1.14 ;
 RECT 5.97 1.14 6.47 1.37 ;
 RECT 5.97 1.37 6.07 2.385 ;
 RECT 6.815 0.505 6.915 2.585 ;
 RECT 5.035 2.455 5.265 2.585 ;
 RECT 5.035 2.585 6.915 2.685 ;
 RECT 7.285 0.51 7.385 1.155 ;
 RECT 7.095 1.155 7.385 1.385 ;
 RECT 7.285 1.385 7.385 2.35 ;
 RECT 8.135 0.14 8.235 1.02 ;
 RECT 7.97 1.02 8.235 1.255 ;
 RECT 8.135 1.255 8.235 2.79 ;
 RECT 3.535 1.22 3.755 1.37 ;
 RECT 3.535 1.12 4.13 1.22 ;
 RECT 4.03 0.43 4.13 1.12 ;
 RECT 4.03 0.33 5.07 0.43 ;
 RECT 4.97 0.43 5.07 1.835 ;
 RECT 4.285 1.835 5.07 1.935 ;
 RECT 4.285 1.935 4.385 2.48 ;
 RECT 3.615 0.235 3.845 0.315 ;
 RECT 3.615 0.415 3.845 0.465 ;
 RECT 1.485 0.315 3.845 0.415 ;
 RECT 1.485 0.415 1.585 1.305 ;
 RECT 1.485 1.305 1.755 1.405 ;
 RECT 1.655 1.405 1.755 2.365 ;
 RECT 3.175 0.595 3.275 1.095 ;
 RECT 2.97 1.095 3.275 1.195 ;
 RECT 4.5 0.61 4.6 1.55 ;
 RECT 2.97 1.195 3.07 1.58 ;
 RECT 3.815 1.55 4.6 1.65 ;
 RECT 2.8 1.58 3.07 1.81 ;
 RECT 3.815 1.65 3.915 2.485 ;
 RECT 2.97 1.81 3.07 2.485 ;
 RECT 2.97 2.485 3.915 2.585 ;
 RECT 5.5 0.355 5.79 0.565 ;
 RECT 5.5 0.565 5.6 2.385 ;
 LAYER CO ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 1.08 1.225 1.21 1.355 ;
 RECT 6.29 1.19 6.42 1.32 ;
 RECT 7.885 1.625 8.015 1.755 ;
 RECT 7.145 1.205 7.275 1.335 ;
 RECT 7.505 1.99 7.635 2.12 ;
 RECT 6.565 1.99 6.695 2.12 ;
 RECT 7.035 1.975 7.165 2.105 ;
 RECT 7.505 0.74 7.635 0.87 ;
 RECT 6.19 1.99 6.32 2.12 ;
 RECT 5.25 1.99 5.38 2.12 ;
 RECT 5.72 1.99 5.85 2.12 ;
 RECT 6.19 0.835 6.32 0.965 ;
 RECT 5.24 0.125 5.37 0.255 ;
 RECT 1.705 0.835 1.835 0.965 ;
 RECT 7.885 0.48 8.015 0.61 ;
 RECT 7.885 0.74 8.015 0.87 ;
 RECT 3.665 0.285 3.795 0.415 ;
 RECT 5.085 2.495 5.215 2.625 ;
 RECT 3.395 0.835 3.525 0.965 ;
 RECT 6.56 0.74 6.69 0.87 ;
 RECT 8.355 0.465 8.485 0.595 ;
 RECT 8.02 1.07 8.15 1.2 ;
 RECT 8.355 0.725 8.485 0.855 ;
 RECT 7.885 2.145 8.015 2.275 ;
 RECT 8.355 1.625 8.485 1.755 ;
 RECT 7.885 2.405 8.015 2.535 ;
 RECT 8.355 1.885 8.485 2.015 ;
 RECT 8.355 2.145 8.485 2.275 ;
 RECT 7.885 1.885 8.015 2.015 ;
 RECT 8.355 2.405 8.485 2.535 ;
 RECT 7.885 2.145 8.015 2.275 ;
 RECT 7.885 2.405 8.015 2.535 ;
 RECT 2.075 0.835 2.205 0.965 ;
 RECT 3.575 1.19 3.705 1.32 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 4.72 0.835 4.85 0.965 ;
 RECT 4.505 2.125 4.635 2.255 ;
 RECT 5.61 0.395 5.74 0.525 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 3.78 0.835 3.91 0.965 ;
 RECT 3.565 1.995 3.695 2.125 ;
 RECT 4.035 2.125 4.165 2.255 ;
 RECT 2.71 2.61 2.84 2.74 ;
 RECT 1.89 2.64 2.02 2.77 ;
 RECT 2.205 1.23 2.335 1.36 ;
 RECT 2.86 1.63 2.99 1.76 ;
 RECT 2.92 0.835 3.05 0.965 ;
 RECT 3.19 2.035 3.32 2.165 ;
 RECT 2.55 0.835 2.68 0.965 ;
 RECT 2.345 2.005 2.475 2.135 ;
 RECT 1.405 1.995 1.535 2.125 ;
 RECT 0.935 0.835 1.065 0.965 ;
 RECT 0.935 1.995 1.065 2.125 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 LAYER M1 ;
 RECT 4.22 0.76 4.39 1.02 ;
 RECT 4.22 1.02 4.36 1.765 ;
 RECT 4.03 1.765 4.36 1.905 ;
 RECT 4.03 1.905 4.17 2.49 ;
 RECT 4.03 2.49 5.265 2.63 ;
 RECT 2.545 0.785 2.685 1.625 ;
 RECT 2.34 1.625 3.045 1.765 ;
 RECT 2.34 1.765 2.48 2 ;
 RECT 2.295 2 2.525 2.14 ;
 RECT 2.34 2.14 2.48 2.175 ;
 RECT 7.5 0.67 7.64 1.06 ;
 RECT 7.455 1.985 7.685 2.125 ;
 RECT 7.5 1.205 7.64 1.6 ;
 RECT 7.5 1.74 7.64 1.985 ;
 RECT 6.56 1.6 7.64 1.74 ;
 RECT 6.515 1.985 6.745 2.125 ;
 RECT 6.19 1.185 6.7 1.325 ;
 RECT 6.56 1.325 6.7 1.6 ;
 RECT 6.56 1.74 6.7 1.985 ;
 RECT 7.5 1.06 8.21 1.205 ;
 RECT 2.915 0.775 3.055 1.185 ;
 RECT 2.915 1.185 3.755 1.325 ;
 RECT 3.185 1.325 3.325 2.03 ;
 RECT 3.1 2.03 3.37 2.17 ;
 RECT 3.185 2.17 3.325 2.185 ;
 RECT 1.7 0.785 1.84 1.99 ;
 RECT 1.31 1.99 1.84 2.13 ;
 RECT 1.4 2.13 1.54 2.325 ;
 RECT 3.73 0.83 4.08 0.97 ;
 RECT 3.94 0.97 4.08 1.465 ;
 RECT 3.56 1.465 4.08 1.605 ;
 RECT 3.56 1.605 3.7 2.325 ;
 RECT 1.4 2.325 3.7 2.465 ;
 RECT 5.2 1.985 5.43 2.125 ;
 RECT 5.245 1.69 5.385 1.985 ;
 RECT 4.715 0.78 4.855 1.16 ;
 RECT 4.5 1.3 4.64 2.12 ;
 RECT 4.41 2.12 4.695 2.26 ;
 RECT 6.14 1.985 6.37 2.125 ;
 RECT 6.185 1.69 6.325 1.985 ;
 RECT 5.715 0.83 6.37 0.97 ;
 RECT 5.245 1.55 6.325 1.69 ;
 RECT 5.715 0.97 5.855 1.16 ;
 RECT 5.715 1.3 5.855 1.55 ;
 RECT 4.5 1.16 5.855 1.3 ;
 END
END LASRNX1

MACRO LASRNX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.6 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.96 1.28 1.275 1.6 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.98 1.16 2.34 1.485 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.015 1.11 7.35 1.435 ;
 END
 ANTENNAGATEAREA 0.06 ;
 END SETB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.6 2.96 ;
 RECT 1.84 2.63 2.07 2.8 ;
 RECT 2.66 2.605 2.89 2.8 ;
 RECT 7.03 1.905 7.17 2.8 ;
 RECT 5.715 1.9 5.855 2.8 ;
 RECT 0.93 1.88 1.07 2.8 ;
 RECT 8.375 1.775 8.515 2.8 ;
 RECT 0.425 1.755 0.565 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.6 0.08 ;
 RECT 3.32 0.08 3.46 0.825 ;
 RECT 0.34 0.08 0.48 0.81 ;
 RECT 0.93 0.08 1.07 1.025 ;
 RECT 2.07 0.08 2.21 1.02 ;
 RECT 5.19 0.08 5.42 0.29 ;
 RECT 6.715 0.08 6.855 0.78 ;
 RECT 8.32 0.08 8.55 0.295 ;
 RECT 3.32 0.825 3.575 0.97 ;
 RECT 6.51 0.78 6.855 0.94 ;
 END
 END VSS

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.6 0.32 5.92 0.39 ;
 RECT 3.66 0.235 3.8 0.46 ;
 RECT 5.6 0.6 5.92 0.64 ;
 RECT 3.66 0.46 5.92 0.6 ;
 RECT 5.56 0.39 5.92 0.46 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.845 2.075 9.28 2.405 ;
 RECT 8.845 2.405 8.985 2.65 ;
 RECT 8.845 1.615 8.985 2.075 ;
 RECT 7.895 1.475 8.985 1.615 ;
 RECT 7.895 1.615 8.035 2.66 ;
 RECT 7.895 0.905 8.035 1.475 ;
 RECT 8.845 0.4 8.985 1.475 ;
 RECT 7.835 0.765 8.085 0.905 ;
 END
 ANTENNADIFFAREA 0.977 ;
 END QN

 OBS
 LAYER PO ;
 RECT 2.33 0.595 2.43 1.18 ;
 RECT 2.01 1.18 2.43 1.41 ;
 RECT 2.125 1.41 2.225 2.375 ;
 RECT 5.97 0.61 6.07 1.14 ;
 RECT 5.97 1.14 6.47 1.37 ;
 RECT 5.97 1.37 6.07 2.385 ;
 RECT 7.285 0.545 7.385 1.155 ;
 RECT 7.095 1.155 7.385 1.385 ;
 RECT 7.285 1.385 7.385 2.35 ;
 RECT 3.535 1.22 3.755 1.37 ;
 RECT 3.535 1.12 4.13 1.22 ;
 RECT 4.03 0.43 4.13 1.12 ;
 RECT 4.03 0.33 5.07 0.43 ;
 RECT 4.97 0.43 5.07 1.835 ;
 RECT 4.285 1.835 5.07 1.935 ;
 RECT 4.285 1.935 4.385 2.48 ;
 RECT 3.175 0.595 3.275 1.095 ;
 RECT 2.97 1.095 3.275 1.195 ;
 RECT 4.5 0.61 4.6 1.55 ;
 RECT 2.97 1.195 3.07 1.58 ;
 RECT 3.815 1.55 4.6 1.65 ;
 RECT 2.8 1.58 3.07 1.81 ;
 RECT 3.815 1.65 3.915 2.485 ;
 RECT 2.97 1.81 3.07 2.485 ;
 RECT 2.97 2.485 3.915 2.585 ;
 RECT 3.615 0.235 3.845 0.315 ;
 RECT 3.615 0.415 3.845 0.465 ;
 RECT 1.485 0.315 3.845 0.415 ;
 RECT 1.485 0.415 1.585 1.305 ;
 RECT 1.485 1.305 1.755 1.405 ;
 RECT 1.655 1.405 1.755 2.365 ;
 RECT 5.035 2.455 5.265 2.585 ;
 RECT 6.815 0.56 6.915 2.585 ;
 RECT 5.035 2.585 6.915 2.685 ;
 RECT 8.63 1.345 8.73 2.685 ;
 RECT 8.15 0.185 8.25 2.685 ;
 RECT 8.63 0.14 8.73 1.115 ;
 RECT 8.435 1.115 8.73 1.345 ;
 RECT 8.15 2.685 8.73 2.785 ;
 RECT 5.5 0.39 5.79 0.6 ;
 RECT 5.5 0.6 5.6 2.385 ;
 RECT 1.185 0.615 1.285 1.355 ;
 RECT 1 1.355 1.285 1.565 ;
 RECT 1.185 1.565 1.285 2.37 ;
 LAYER CO ;
 RECT 3.575 1.19 3.705 1.32 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 4.72 0.835 4.85 0.965 ;
 RECT 4.505 2.125 4.635 2.255 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 3.78 0.835 3.91 0.965 ;
 RECT 3.565 1.995 3.695 2.125 ;
 RECT 4.035 2.125 4.165 2.255 ;
 RECT 2.71 2.61 2.84 2.74 ;
 RECT 1.89 2.64 2.02 2.77 ;
 RECT 2.06 1.23 2.19 1.36 ;
 RECT 2.86 1.63 2.99 1.76 ;
 RECT 2.92 0.835 3.05 0.965 ;
 RECT 3.19 2.035 3.32 2.165 ;
 RECT 2.55 0.835 2.68 0.965 ;
 RECT 2.345 2.005 2.475 2.135 ;
 RECT 1.405 1.995 1.535 2.125 ;
 RECT 0.935 0.835 1.065 0.965 ;
 RECT 0.935 1.995 1.065 2.125 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 8.485 1.165 8.615 1.295 ;
 RECT 7.9 1.625 8.03 1.755 ;
 RECT 7.9 1.885 8.03 2.015 ;
 RECT 8.85 0.51 8.98 0.64 ;
 RECT 8.85 2.405 8.98 2.535 ;
 RECT 7.9 2.145 8.03 2.275 ;
 RECT 8.38 2.145 8.51 2.275 ;
 RECT 6.29 1.19 6.42 1.32 ;
 RECT 7.145 1.205 7.275 1.335 ;
 RECT 7.505 1.99 7.635 2.12 ;
 RECT 6.565 1.99 6.695 2.12 ;
 RECT 5.61 0.43 5.74 0.56 ;
 RECT 1.05 1.395 1.18 1.525 ;
 RECT 7.035 1.975 7.165 2.105 ;
 RECT 7.505 0.79 7.635 0.92 ;
 RECT 6.19 1.99 6.32 2.12 ;
 RECT 5.25 1.99 5.38 2.12 ;
 RECT 5.72 1.99 5.85 2.12 ;
 RECT 6.19 0.835 6.32 0.965 ;
 RECT 5.24 0.125 5.37 0.255 ;
 RECT 1.705 0.835 1.835 0.965 ;
 RECT 7.9 2.405 8.03 2.535 ;
 RECT 8.85 0.77 8.98 0.9 ;
 RECT 8.38 2.405 8.51 2.535 ;
 RECT 7.9 1.625 8.03 1.755 ;
 RECT 8.38 2.145 8.51 2.275 ;
 RECT 7.9 0.77 8.03 0.9 ;
 RECT 7.9 1.885 8.03 2.015 ;
 RECT 8.85 1.625 8.98 1.755 ;
 RECT 7.9 2.145 8.03 2.275 ;
 RECT 8.38 2.405 8.51 2.535 ;
 RECT 8.85 1.885 8.98 2.015 ;
 RECT 8.85 2.145 8.98 2.275 ;
 RECT 8.37 0.115 8.5 0.245 ;
 RECT 8.38 1.885 8.51 2.015 ;
 RECT 7.9 2.405 8.03 2.535 ;
 RECT 3.665 0.285 3.795 0.415 ;
 RECT 5.085 2.505 5.215 2.635 ;
 RECT 3.395 0.835 3.525 0.965 ;
 RECT 6.56 0.79 6.69 0.92 ;
 RECT 2.075 0.835 2.205 0.965 ;
 LAYER M1 ;
 RECT 4.22 0.77 4.39 1.02 ;
 RECT 4.22 1.02 4.36 1.775 ;
 RECT 4.03 1.775 4.36 1.915 ;
 RECT 4.03 1.915 4.17 2.5 ;
 RECT 4.03 2.5 5.265 2.64 ;
 RECT 2.545 0.785 2.685 1.625 ;
 RECT 2.34 1.625 3.045 1.765 ;
 RECT 2.34 1.765 2.48 2 ;
 RECT 2.295 2 2.525 2.14 ;
 RECT 2.34 2.14 2.48 2.175 ;
 RECT 2.915 0.775 3.055 1.185 ;
 RECT 2.915 1.185 3.755 1.325 ;
 RECT 3.185 1.325 3.325 2.03 ;
 RECT 3.1 2.03 3.37 2.17 ;
 RECT 3.185 2.17 3.325 2.185 ;
 RECT 6.19 1.185 6.7 1.325 ;
 RECT 6.56 1.325 6.7 1.58 ;
 RECT 6.56 1.72 6.7 1.985 ;
 RECT 7.455 1.985 7.685 2.125 ;
 RECT 7.5 0.575 7.64 1.58 ;
 RECT 7.5 1.72 7.64 1.985 ;
 RECT 6.56 1.58 7.64 1.72 ;
 RECT 6.515 1.985 6.745 2.125 ;
 RECT 8.415 1.16 8.7 1.3 ;
 RECT 8.415 0.575 8.555 1.16 ;
 RECT 7.5 0.435 8.555 0.575 ;
 RECT 1.7 0.785 1.84 1.99 ;
 RECT 1.31 1.99 1.84 2.13 ;
 RECT 1.4 2.13 1.54 2.325 ;
 RECT 3.73 0.83 4.08 0.97 ;
 RECT 3.94 0.97 4.08 1.465 ;
 RECT 3.56 1.465 4.08 1.605 ;
 RECT 3.56 1.605 3.7 2.325 ;
 RECT 1.4 2.325 3.7 2.465 ;
 RECT 5.2 1.985 5.43 2.125 ;
 RECT 5.245 1.69 5.385 1.985 ;
 RECT 4.715 0.78 4.855 1.16 ;
 RECT 4.5 1.3 4.64 2.12 ;
 RECT 4.41 2.12 4.695 2.26 ;
 RECT 6.14 1.985 6.37 2.125 ;
 RECT 6.185 1.69 6.325 1.985 ;
 RECT 5.715 0.83 6.37 0.97 ;
 RECT 5.24 1.55 6.325 1.69 ;
 RECT 5.715 0.97 5.855 1.16 ;
 RECT 5.715 1.3 5.855 1.55 ;
 RECT 4.5 1.16 5.855 1.3 ;
 END
END LASRNX2

MACRO LASRQX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.96 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.94 1.155 1.275 1.45 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.12 1.16 2.385 1.45 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.045 1.1 7.35 1.41 ;
 END
 ANTENNAGATEAREA 0.06 ;
 END SETB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.96 2.96 ;
 RECT 1.84 2.63 2.07 2.8 ;
 RECT 2.66 2.605 2.89 2.8 ;
 RECT 7.03 1.905 7.17 2.8 ;
 RECT 5.715 1.9 5.855 2.8 ;
 RECT 0.93 1.88 1.07 2.8 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 7.88 1.485 8.02 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.96 0.08 ;
 RECT 3.32 0.08 3.46 0.83 ;
 RECT 0.34 0.08 0.48 0.825 ;
 RECT 0.93 0.08 1.07 1.015 ;
 RECT 2.07 0.08 2.21 1.015 ;
 RECT 5.19 0.08 5.42 0.305 ;
 RECT 6.715 0.08 6.855 0.735 ;
 RECT 7.88 0.08 8.02 0.92 ;
 RECT 3.32 0.83 3.575 0.97 ;
 RECT 6.51 0.735 6.855 0.875 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.31 2.105 8.635 2.395 ;
 RECT 8.35 2.395 8.49 2.61 ;
 RECT 8.35 0.4 8.49 2.105 ;
 END
 ANTENNADIFFAREA 0.472 ;
 END Q

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.66 0.46 5.895 0.6 ;
 RECT 5.56 0.345 5.895 0.46 ;
 RECT 3.66 0.235 3.8 0.46 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 OBS
 LAYER PO ;
 RECT 1.185 0.615 1.285 1.175 ;
 RECT 1.03 1.175 1.285 1.405 ;
 RECT 1.185 1.405 1.285 2.37 ;
 RECT 2.33 0.595 2.43 1.18 ;
 RECT 2.125 1.18 2.43 1.41 ;
 RECT 2.125 1.41 2.225 2.375 ;
 RECT 5.97 0.615 6.07 1.14 ;
 RECT 5.97 1.14 6.47 1.37 ;
 RECT 5.97 1.37 6.07 2.385 ;
 RECT 6.815 0.52 6.915 2.585 ;
 RECT 5.035 2.455 5.265 2.585 ;
 RECT 5.035 2.585 6.915 2.685 ;
 RECT 7.285 0.52 7.385 1.155 ;
 RECT 7.095 1.155 7.385 1.385 ;
 RECT 7.285 1.385 7.385 2.35 ;
 RECT 3.535 1.22 3.755 1.37 ;
 RECT 3.535 1.12 4.13 1.22 ;
 RECT 4.03 0.43 4.13 1.12 ;
 RECT 4.03 0.33 5.07 0.43 ;
 RECT 4.97 0.43 5.07 1.835 ;
 RECT 4.285 1.835 5.07 1.935 ;
 RECT 4.285 1.935 4.385 2.48 ;
 RECT 8.135 0.34 8.235 2.785 ;
 RECT 6.27 0.24 8.235 0.34 ;
 RECT 6.27 0.34 6.5 0.47 ;
 RECT 3.175 0.595 3.275 1.095 ;
 RECT 2.97 1.095 3.275 1.195 ;
 RECT 4.5 0.61 4.6 1.55 ;
 RECT 2.97 1.195 3.07 1.58 ;
 RECT 3.815 1.55 4.6 1.65 ;
 RECT 2.8 1.58 3.07 1.81 ;
 RECT 3.815 1.65 3.915 2.485 ;
 RECT 2.97 1.81 3.07 2.485 ;
 RECT 2.97 2.485 3.915 2.585 ;
 RECT 3.615 0.235 3.845 0.315 ;
 RECT 3.615 0.415 3.845 0.465 ;
 RECT 1.485 0.315 3.845 0.415 ;
 RECT 1.485 0.415 1.585 1.305 ;
 RECT 1.485 1.305 1.755 1.405 ;
 RECT 1.655 1.405 1.755 2.365 ;
 RECT 5.5 0.35 5.79 0.56 ;
 RECT 5.5 0.56 5.6 2.385 ;
 LAYER CO ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 1.08 1.225 1.21 1.355 ;
 RECT 6.29 1.19 6.42 1.32 ;
 RECT 7.885 1.625 8.015 1.755 ;
 RECT 7.145 1.205 7.275 1.335 ;
 RECT 7.505 1.99 7.635 2.12 ;
 RECT 6.565 1.99 6.695 2.12 ;
 RECT 7.035 1.975 7.165 2.105 ;
 RECT 7.505 0.74 7.635 0.87 ;
 RECT 6.19 1.99 6.32 2.12 ;
 RECT 5.25 1.99 5.38 2.12 ;
 RECT 5.72 1.99 5.85 2.12 ;
 RECT 6.19 0.835 6.32 0.965 ;
 RECT 5.24 0.125 5.37 0.255 ;
 RECT 1.705 0.835 1.835 0.965 ;
 RECT 6.32 0.29 6.45 0.42 ;
 RECT 7.885 0.48 8.015 0.61 ;
 RECT 7.885 0.74 8.015 0.87 ;
 RECT 3.665 0.285 3.795 0.415 ;
 RECT 5.085 2.495 5.215 2.625 ;
 RECT 3.395 0.835 3.525 0.965 ;
 RECT 6.56 0.74 6.69 0.87 ;
 RECT 8.355 0.465 8.485 0.595 ;
 RECT 8.355 0.725 8.485 0.855 ;
 RECT 7.885 2.145 8.015 2.275 ;
 RECT 8.355 1.625 8.485 1.755 ;
 RECT 7.885 2.405 8.015 2.535 ;
 RECT 8.355 1.885 8.485 2.015 ;
 RECT 8.355 2.145 8.485 2.275 ;
 RECT 7.885 1.885 8.015 2.015 ;
 RECT 8.355 2.405 8.485 2.535 ;
 RECT 7.885 2.145 8.015 2.275 ;
 RECT 7.885 2.405 8.015 2.535 ;
 RECT 2.075 0.835 2.205 0.965 ;
 RECT 3.575 1.19 3.705 1.32 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 4.72 0.835 4.85 0.965 ;
 RECT 4.505 2.125 4.635 2.255 ;
 RECT 5.61 0.39 5.74 0.52 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 3.78 0.835 3.91 0.965 ;
 RECT 3.565 1.995 3.695 2.125 ;
 RECT 4.035 2.125 4.165 2.255 ;
 RECT 2.71 2.61 2.84 2.74 ;
 RECT 1.89 2.64 2.02 2.77 ;
 RECT 2.205 1.23 2.335 1.36 ;
 RECT 2.86 1.63 2.99 1.76 ;
 RECT 2.92 0.835 3.05 0.965 ;
 RECT 3.19 2.035 3.32 2.165 ;
 RECT 2.55 0.835 2.68 0.965 ;
 RECT 2.345 2.005 2.475 2.135 ;
 RECT 1.405 1.995 1.535 2.125 ;
 RECT 0.935 0.835 1.065 0.965 ;
 RECT 0.935 1.995 1.065 2.125 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 LAYER M1 ;
 RECT 4.22 0.76 4.39 1.02 ;
 RECT 4.22 1.02 4.36 1.765 ;
 RECT 4.03 1.765 4.36 1.905 ;
 RECT 4.03 1.905 4.17 2.49 ;
 RECT 4.03 2.49 5.265 2.63 ;
 RECT 2.545 0.785 2.685 1.625 ;
 RECT 2.34 1.625 3.045 1.765 ;
 RECT 2.34 1.765 2.48 2 ;
 RECT 2.295 2 2.525 2.14 ;
 RECT 2.34 2.14 2.48 2.175 ;
 RECT 4.715 0.78 4.855 1.16 ;
 RECT 4.5 1.3 4.64 2.12 ;
 RECT 4.41 2.12 4.695 2.26 ;
 RECT 5.2 1.985 5.43 2.125 ;
 RECT 5.245 1.69 5.385 1.985 ;
 RECT 6.23 0.24 6.5 0.47 ;
 RECT 6.14 1.985 6.37 2.125 ;
 RECT 6.23 0.47 6.37 0.83 ;
 RECT 6.185 1.69 6.325 1.985 ;
 RECT 5.715 0.83 6.37 0.97 ;
 RECT 5.245 1.55 6.325 1.69 ;
 RECT 5.715 0.97 5.855 1.16 ;
 RECT 5.715 1.3 5.855 1.55 ;
 RECT 4.5 1.16 5.855 1.3 ;
 RECT 2.915 0.775 3.055 1.185 ;
 RECT 2.915 1.185 3.755 1.325 ;
 RECT 3.185 1.325 3.325 2.03 ;
 RECT 3.1 2.03 3.37 2.17 ;
 RECT 3.185 2.17 3.325 2.185 ;
 RECT 1.7 0.785 1.84 1.99 ;
 RECT 1.31 1.99 1.84 2.13 ;
 RECT 1.4 2.13 1.54 2.325 ;
 RECT 3.73 0.83 4.08 0.97 ;
 RECT 3.94 0.97 4.08 1.465 ;
 RECT 3.56 1.465 4.08 1.605 ;
 RECT 3.56 1.605 3.7 2.325 ;
 RECT 1.4 2.325 3.7 2.465 ;
 RECT 6.19 1.185 6.7 1.325 ;
 RECT 6.56 1.325 6.7 1.58 ;
 RECT 6.56 1.72 6.7 1.985 ;
 RECT 6.515 1.985 6.745 2.125 ;
 RECT 7.455 1.985 7.685 2.125 ;
 RECT 7.5 0.685 7.64 1.58 ;
 RECT 7.5 1.72 7.64 1.985 ;
 RECT 6.56 1.58 7.64 1.72 ;
 END
END LASRQX1

MACRO LASRQX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.28 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.95 1.16 1.275 1.475 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.085 1.16 2.39 1.45 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.01 1.125 7.35 1.43 ;
 END
 ANTENNAGATEAREA 0.06 ;
 END SETB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.28 2.96 ;
 RECT 1.84 2.63 2.07 2.8 ;
 RECT 2.66 2.605 2.89 2.8 ;
 RECT 7.03 1.905 7.17 2.8 ;
 RECT 5.715 1.9 5.855 2.8 ;
 RECT 0.93 1.88 1.07 2.8 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 8.365 1.495 8.505 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.28 0.08 ;
 RECT 6.715 0.08 6.855 0.83 ;
 RECT 0.34 0.08 0.48 0.81 ;
 RECT 0.93 0.08 1.07 1.015 ;
 RECT 2.07 0.08 2.21 1.02 ;
 RECT 3.32 0.08 3.46 0.825 ;
 RECT 5.19 0.08 5.42 0.29 ;
 RECT 8.365 0.08 8.505 0.94 ;
 RECT 6.51 0.83 6.855 0.97 ;
 RECT 3.32 0.825 3.575 0.97 ;
 END
 END VSS

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.66 0.46 5.91 0.6 ;
 RECT 5.56 0.33 5.91 0.46 ;
 RECT 3.66 0.235 3.8 0.46 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.825 2.095 8.15 2.375 ;
 RECT 7.885 1.31 8.025 2.095 ;
 RECT 7.885 1.17 8.975 1.31 ;
 RECT 8.835 1.31 8.975 2.64 ;
 RECT 8.835 0.41 8.975 1.17 ;
 RECT 7.885 0.395 8.025 1.17 ;
 END
 ANTENNADIFFAREA 0.904 ;
 END Q

 OBS
 LAYER PO ;
 RECT 1.185 0.615 1.285 1.175 ;
 RECT 1.03 1.175 1.285 1.405 ;
 RECT 1.185 1.405 1.285 2.37 ;
 RECT 2.33 0.595 2.43 1.18 ;
 RECT 2.125 1.18 2.43 1.41 ;
 RECT 2.125 1.41 2.225 2.375 ;
 RECT 5.97 0.615 6.07 1.14 ;
 RECT 5.97 1.14 6.47 1.37 ;
 RECT 5.97 1.37 6.07 2.385 ;
 RECT 7.285 0.61 7.385 1.155 ;
 RECT 7.095 1.155 7.385 1.385 ;
 RECT 7.285 1.385 7.385 2.35 ;
 RECT 3.535 1.22 3.755 1.37 ;
 RECT 3.535 1.12 4.13 1.22 ;
 RECT 4.03 0.43 4.13 1.12 ;
 RECT 4.03 0.33 5.07 0.43 ;
 RECT 4.97 0.43 5.07 1.835 ;
 RECT 4.285 1.835 5.07 1.935 ;
 RECT 4.285 1.935 4.385 2.48 ;
 RECT 6.815 0.615 6.915 2.585 ;
 RECT 5.035 2.455 5.265 2.585 ;
 RECT 5.035 2.585 6.915 2.685 ;
 RECT 6.285 0.255 6.515 0.42 ;
 RECT 6.28 0.155 8.24 0.255 ;
 RECT 8.62 0.14 8.72 1.02 ;
 RECT 8.14 0.255 8.24 1.02 ;
 RECT 8.62 1.255 8.72 2.685 ;
 RECT 8.14 1.02 8.72 1.255 ;
 RECT 8.14 1.255 8.24 2.68 ;
 RECT 3.175 0.595 3.275 1.095 ;
 RECT 2.97 1.095 3.275 1.195 ;
 RECT 4.5 0.61 4.6 1.55 ;
 RECT 2.97 1.195 3.07 1.58 ;
 RECT 3.815 1.55 4.6 1.65 ;
 RECT 2.8 1.58 3.07 1.81 ;
 RECT 3.815 1.65 3.915 2.485 ;
 RECT 2.97 1.81 3.07 2.485 ;
 RECT 2.97 2.485 3.915 2.585 ;
 RECT 3.615 0.235 3.845 0.315 ;
 RECT 3.615 0.415 3.845 0.465 ;
 RECT 1.485 0.315 3.845 0.415 ;
 RECT 1.485 0.415 1.585 1.305 ;
 RECT 1.485 1.305 1.755 1.405 ;
 RECT 1.655 1.405 1.755 2.365 ;
 RECT 5.5 0.39 5.79 0.6 ;
 RECT 5.5 0.6 5.6 2.385 ;
 LAYER CO ;
 RECT 7.89 0.725 8.02 0.855 ;
 RECT 8.84 1.635 8.97 1.765 ;
 RECT 8.84 1.895 8.97 2.025 ;
 RECT 8.84 2.155 8.97 2.285 ;
 RECT 8.37 1.895 8.5 2.025 ;
 RECT 3.665 0.285 3.795 0.415 ;
 RECT 5.085 2.505 5.215 2.635 ;
 RECT 3.395 0.835 3.525 0.965 ;
 RECT 6.335 0.24 6.465 0.37 ;
 RECT 6.56 0.835 6.69 0.965 ;
 RECT 2.075 0.835 2.205 0.965 ;
 RECT 3.575 1.19 3.705 1.32 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 4.72 0.835 4.85 0.965 ;
 RECT 4.505 2.125 4.635 2.255 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 3.78 0.835 3.91 0.965 ;
 RECT 3.565 1.995 3.695 2.125 ;
 RECT 4.035 2.125 4.165 2.255 ;
 RECT 2.71 2.61 2.84 2.74 ;
 RECT 1.89 2.64 2.02 2.77 ;
 RECT 2.235 1.23 2.365 1.36 ;
 RECT 2.86 1.63 2.99 1.76 ;
 RECT 2.92 0.835 3.05 0.965 ;
 RECT 3.19 2.035 3.32 2.165 ;
 RECT 2.55 0.835 2.68 0.965 ;
 RECT 2.345 2.005 2.475 2.135 ;
 RECT 1.405 1.995 1.535 2.125 ;
 RECT 0.935 0.835 1.065 0.965 ;
 RECT 0.935 1.995 1.065 2.125 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 5.61 0.43 5.74 0.56 ;
 RECT 1.08 1.225 1.21 1.355 ;
 RECT 6.29 1.19 6.42 1.32 ;
 RECT 7.145 1.205 7.275 1.335 ;
 RECT 7.505 1.99 7.635 2.12 ;
 RECT 6.565 1.99 6.695 2.12 ;
 RECT 7.035 1.975 7.165 2.105 ;
 RECT 7.505 0.835 7.635 0.965 ;
 RECT 6.19 1.99 6.32 2.12 ;
 RECT 5.25 1.99 5.38 2.12 ;
 RECT 5.72 1.99 5.85 2.12 ;
 RECT 6.19 0.835 6.32 0.965 ;
 RECT 5.24 0.125 5.37 0.255 ;
 RECT 1.705 0.835 1.835 0.965 ;
 RECT 8.84 0.465 8.97 0.595 ;
 RECT 8.37 0.485 8.5 0.615 ;
 RECT 8.37 0.745 8.5 0.875 ;
 RECT 7.89 0.465 8.02 0.595 ;
 RECT 8.37 1.635 8.5 1.765 ;
 RECT 7.89 1.635 8.02 1.765 ;
 RECT 7.89 1.895 8.02 2.025 ;
 RECT 7.89 2.155 8.02 2.285 ;
 RECT 8.37 2.155 8.5 2.285 ;
 RECT 8.84 0.725 8.97 0.855 ;
 RECT 8.37 2.155 8.5 2.285 ;
 LAYER M1 ;
 RECT 4.22 0.77 4.39 1.02 ;
 RECT 4.22 1.02 4.36 1.775 ;
 RECT 4.03 1.775 4.36 1.915 ;
 RECT 4.03 1.915 4.17 2.5 ;
 RECT 4.03 2.5 5.265 2.64 ;
 RECT 2.545 0.785 2.685 1.625 ;
 RECT 2.34 1.625 3.045 1.765 ;
 RECT 2.34 1.765 2.48 2 ;
 RECT 2.295 2 2.525 2.14 ;
 RECT 2.34 2.14 2.48 2.175 ;
 RECT 5.2 1.985 5.43 2.125 ;
 RECT 5.245 1.69 5.385 1.985 ;
 RECT 6.14 1.985 6.37 2.125 ;
 RECT 6.23 0.375 6.37 0.83 ;
 RECT 6.185 1.69 6.325 1.985 ;
 RECT 5.715 0.83 6.37 0.97 ;
 RECT 5.24 1.55 6.325 1.69 ;
 RECT 5.715 0.97 5.855 1.16 ;
 RECT 5.715 1.3 5.855 1.55 ;
 RECT 4.5 1.16 5.855 1.3 ;
 RECT 4.715 0.78 4.855 1.16 ;
 RECT 4.5 1.3 4.64 2.12 ;
 RECT 4.41 2.12 4.695 2.26 ;
 RECT 6.23 0.235 6.515 0.375 ;
 RECT 2.915 0.775 3.055 1.185 ;
 RECT 2.915 1.185 3.755 1.325 ;
 RECT 3.185 1.325 3.325 2.03 ;
 RECT 3.1 2.03 3.37 2.17 ;
 RECT 3.185 2.17 3.325 2.185 ;
 RECT 1.7 0.785 1.84 1.99 ;
 RECT 1.31 1.99 1.84 2.13 ;
 RECT 1.4 2.13 1.54 2.325 ;
 RECT 3.73 0.83 4.08 0.97 ;
 RECT 3.94 0.97 4.08 1.465 ;
 RECT 3.56 1.465 4.08 1.605 ;
 RECT 3.56 1.605 3.7 2.325 ;
 RECT 1.4 2.325 3.7 2.465 ;
 RECT 6.19 1.185 6.7 1.325 ;
 RECT 6.56 1.325 6.7 1.57 ;
 RECT 6.56 1.71 6.7 1.985 ;
 RECT 6.515 1.985 6.745 2.125 ;
 RECT 7.455 1.985 7.685 2.125 ;
 RECT 7.5 0.765 7.64 1.57 ;
 RECT 7.5 1.71 7.64 1.985 ;
 RECT 6.56 1.57 7.64 1.71 ;
 END
END LASRQX2

MACRO LASRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.28 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.9 1.305 1.275 1.64 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.125 1.16 2.365 1.47 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.835 2.43 8.12 2.66 ;
 RECT 7.895 0.86 8.035 2.43 ;
 RECT 7.84 0.72 8.07 0.86 ;
 END
 ANTENNADIFFAREA 0.505 ;
 END Q

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.055 1.13 7.35 1.405 ;
 END
 ANTENNAGATEAREA 0.06 ;
 END SETB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.28 2.96 ;
 RECT 1.84 2.54 2.07 2.8 ;
 RECT 2.66 2.51 2.89 2.8 ;
 RECT 7.03 1.905 7.17 2.8 ;
 RECT 5.715 1.9 5.855 2.8 ;
 RECT 0.93 1.88 1.07 2.8 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 8.375 1.495 8.515 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.28 0.08 ;
 RECT 3.32 0.08 3.46 0.825 ;
 RECT 0.34 0.08 0.48 0.81 ;
 RECT 0.93 0.08 1.07 1.025 ;
 RECT 2.07 0.08 2.21 1.02 ;
 RECT 5.19 0.08 5.42 0.29 ;
 RECT 6.715 0.08 6.855 0.74 ;
 RECT 8.32 0.08 8.55 0.275 ;
 RECT 3.32 0.825 3.575 0.97 ;
 RECT 6.51 0.74 6.855 0.88 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.655 2.28 9.035 2.545 ;
 RECT 8.845 0.4 8.985 2.28 ;
 END
 ANTENNADIFFAREA 0.472 ;
 END QN

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.66 0.46 5.88 0.6 ;
 RECT 5.56 0.36 5.88 0.46 ;
 RECT 3.66 0.235 3.8 0.46 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 OBS
 LAYER PO ;
 RECT 5.97 0.615 6.07 1.14 ;
 RECT 5.97 1.14 6.47 1.37 ;
 RECT 5.97 1.37 6.07 2.385 ;
 RECT 6.815 0.515 6.915 2.585 ;
 RECT 5.035 2.455 5.265 2.585 ;
 RECT 5.035 2.585 6.915 2.685 ;
 RECT 7.285 0.515 7.385 1.155 ;
 RECT 7.095 1.155 7.385 1.385 ;
 RECT 7.285 1.385 7.385 2.35 ;
 RECT 8.63 0.14 8.73 1.02 ;
 RECT 8.465 1.02 8.73 1.255 ;
 RECT 8.63 1.255 8.73 2.79 ;
 RECT 3.535 1.22 3.755 1.37 ;
 RECT 3.535 1.12 4.13 1.22 ;
 RECT 4.03 0.43 4.13 1.12 ;
 RECT 4.03 0.33 5.07 0.43 ;
 RECT 4.97 0.43 5.07 1.835 ;
 RECT 4.285 1.835 5.07 1.935 ;
 RECT 4.285 1.935 4.385 2.48 ;
 RECT 8.15 0.255 8.25 2.79 ;
 RECT 6.285 0.155 8.25 0.255 ;
 RECT 6.285 0.255 6.515 0.42 ;
 RECT 3.175 0.595 3.275 1.095 ;
 RECT 2.97 1.095 3.275 1.195 ;
 RECT 4.5 0.61 4.6 1.55 ;
 RECT 2.97 1.195 3.07 1.58 ;
 RECT 3.815 1.55 4.6 1.65 ;
 RECT 2.8 1.58 3.07 1.81 ;
 RECT 3.815 1.65 3.915 2.385 ;
 RECT 2.97 1.81 3.07 2.385 ;
 RECT 2.97 2.385 3.915 2.485 ;
 RECT 3.615 0.235 3.845 0.315 ;
 RECT 3.615 0.415 3.845 0.465 ;
 RECT 1.485 0.315 3.845 0.415 ;
 RECT 1.485 0.415 1.585 1.305 ;
 RECT 1.485 1.305 1.755 1.405 ;
 RECT 1.655 1.405 1.755 2.365 ;
 RECT 5.5 0.375 5.79 0.585 ;
 RECT 5.5 0.585 5.6 2.385 ;
 RECT 2.33 0.595 2.43 1.18 ;
 RECT 2.125 1.41 2.225 2.255 ;
 RECT 2.125 1.18 2.43 1.41 ;
 RECT 1.185 0.615 1.285 1.365 ;
 RECT 1 1.365 1.285 1.575 ;
 RECT 1.185 1.575 1.285 2.37 ;
 LAYER CO ;
 RECT 7.9 1.625 8.03 1.755 ;
 RECT 7.9 1.885 8.03 2.015 ;
 RECT 7.9 2.145 8.03 2.275 ;
 RECT 7.9 2.405 8.03 2.535 ;
 RECT 7.9 1.625 8.03 1.755 ;
 RECT 7.9 1.885 8.03 2.015 ;
 RECT 7.9 2.145 8.03 2.275 ;
 RECT 7.9 2.405 8.03 2.535 ;
 RECT 7.145 1.205 7.275 1.335 ;
 RECT 7.505 1.99 7.635 2.12 ;
 RECT 6.565 1.99 6.695 2.12 ;
 RECT 7.035 1.975 7.165 2.105 ;
 RECT 7.505 0.745 7.635 0.875 ;
 RECT 6.19 1.99 6.32 2.12 ;
 RECT 5.25 1.99 5.38 2.12 ;
 RECT 5.72 1.99 5.85 2.12 ;
 RECT 6.19 0.835 6.32 0.965 ;
 RECT 5.24 0.125 5.37 0.255 ;
 RECT 1.705 0.835 1.835 0.965 ;
 RECT 3.665 0.285 3.795 0.415 ;
 RECT 5.085 2.505 5.215 2.635 ;
 RECT 3.395 0.835 3.525 0.965 ;
 RECT 6.335 0.24 6.465 0.37 ;
 RECT 6.56 0.745 6.69 0.875 ;
 RECT 8.37 0.11 8.5 0.24 ;
 RECT 8.85 0.465 8.98 0.595 ;
 RECT 8.515 1.07 8.645 1.2 ;
 RECT 8.85 0.725 8.98 0.855 ;
 RECT 8.38 2.145 8.51 2.275 ;
 RECT 8.85 1.625 8.98 1.755 ;
 RECT 8.38 2.405 8.51 2.535 ;
 RECT 8.85 1.885 8.98 2.015 ;
 RECT 5.61 0.415 5.74 0.545 ;
 RECT 2.185 1.23 2.315 1.36 ;
 RECT 1.05 1.405 1.18 1.535 ;
 RECT 8.85 2.145 8.98 2.275 ;
 RECT 8.38 1.885 8.51 2.015 ;
 RECT 8.85 2.405 8.98 2.535 ;
 RECT 8.38 2.145 8.51 2.275 ;
 RECT 8.38 2.405 8.51 2.535 ;
 RECT 7.89 0.725 8.02 0.855 ;
 RECT 2.075 0.835 2.205 0.965 ;
 RECT 3.575 1.19 3.705 1.32 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 4.72 0.835 4.85 0.965 ;
 RECT 4.505 2.125 4.635 2.255 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 3.78 0.835 3.91 0.965 ;
 RECT 3.565 1.995 3.695 2.125 ;
 RECT 4.035 2.125 4.165 2.255 ;
 RECT 2.71 2.515 2.84 2.645 ;
 RECT 1.89 2.545 2.02 2.675 ;
 RECT 2.86 1.63 2.99 1.76 ;
 RECT 2.92 0.835 3.05 0.965 ;
 RECT 3.19 1.935 3.32 2.065 ;
 RECT 2.55 0.835 2.68 0.965 ;
 RECT 2.345 1.885 2.475 2.015 ;
 RECT 1.405 1.995 1.535 2.125 ;
 RECT 0.935 0.835 1.065 0.965 ;
 RECT 0.935 1.995 1.065 2.125 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 6.29 1.19 6.42 1.32 ;
 RECT 8.38 1.625 8.51 1.755 ;
 LAYER M1 ;
 RECT 6.19 1.185 6.7 1.325 ;
 RECT 6.56 1.325 6.7 1.57 ;
 RECT 6.56 1.71 6.7 1.985 ;
 RECT 7.455 1.985 7.685 2.125 ;
 RECT 7.5 0.575 7.64 1.57 ;
 RECT 7.5 1.71 7.64 1.985 ;
 RECT 6.56 1.57 7.64 1.71 ;
 RECT 6.515 1.985 6.745 2.125 ;
 RECT 8.345 1.065 8.695 1.205 ;
 RECT 8.345 0.575 8.485 1.065 ;
 RECT 7.5 0.435 8.485 0.575 ;
 RECT 4.22 0.77 4.39 1.02 ;
 RECT 4.22 1.02 4.36 1.775 ;
 RECT 4.03 1.775 4.36 1.915 ;
 RECT 4.03 1.915 4.17 2.5 ;
 RECT 4.03 2.5 5.265 2.64 ;
 RECT 2.545 0.785 2.685 1.625 ;
 RECT 2.34 1.625 3.045 1.765 ;
 RECT 2.34 1.765 2.525 1.88 ;
 RECT 2.295 1.88 2.525 2.02 ;
 RECT 5.2 1.985 5.43 2.125 ;
 RECT 5.245 1.69 5.385 1.985 ;
 RECT 6.14 1.985 6.37 2.125 ;
 RECT 6.23 0.375 6.37 0.83 ;
 RECT 6.185 1.69 6.325 1.985 ;
 RECT 5.715 0.83 6.37 0.97 ;
 RECT 5.24 1.55 6.325 1.69 ;
 RECT 5.715 0.97 5.855 1.16 ;
 RECT 5.715 1.3 5.855 1.55 ;
 RECT 4.5 1.16 5.855 1.3 ;
 RECT 4.715 0.78 4.855 1.16 ;
 RECT 4.5 1.3 4.64 2.12 ;
 RECT 4.41 2.12 4.695 2.26 ;
 RECT 6.23 0.235 6.515 0.375 ;
 RECT 2.915 0.775 3.055 1.185 ;
 RECT 2.915 1.185 3.755 1.325 ;
 RECT 3.185 1.325 3.325 1.93 ;
 RECT 3.1 1.93 3.37 2.07 ;
 RECT 3.185 2.07 3.325 2.085 ;
 RECT 1.7 0.785 1.84 1.99 ;
 RECT 1.31 1.99 1.84 2.13 ;
 RECT 1.7 2.13 1.84 2.23 ;
 RECT 3.73 0.83 4.08 0.97 ;
 RECT 3.94 0.97 4.08 1.465 ;
 RECT 3.56 1.465 4.08 1.605 ;
 RECT 3.56 1.605 3.7 2.23 ;
 RECT 1.7 2.23 3.7 2.37 ;
 END
END LASRX1

MACRO LASRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.88 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.98 1.32 1.275 1.63 ;
 END
 ANTENNAGATEAREA 0.057 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.09 1.16 2.37 1.45 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.04 1.095 7.35 1.425 ;
 END
 ANTENNAGATEAREA 0.06 ;
 END SETB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.88 2.96 ;
 RECT 1.84 2.63 2.07 2.8 ;
 RECT 2.66 2.605 2.89 2.8 ;
 RECT 7.03 1.905 7.17 2.8 ;
 RECT 5.715 1.9 5.855 2.8 ;
 RECT 0.93 1.88 1.07 2.8 ;
 RECT 9.735 1.76 9.875 2.8 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 8.365 1.47 8.505 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.88 0.08 ;
 RECT 3.32 0.08 3.46 0.825 ;
 RECT 0.34 0.08 0.48 0.81 ;
 RECT 0.93 0.08 1.07 1.025 ;
 RECT 2.07 0.08 2.21 1.02 ;
 RECT 5.19 0.08 5.42 0.29 ;
 RECT 6.715 0.08 6.855 0.735 ;
 RECT 8.305 0.08 8.55 0.275 ;
 RECT 9.68 0.08 9.91 0.295 ;
 RECT 3.32 0.825 3.575 0.97 ;
 RECT 6.51 0.735 6.855 0.885 ;
 END
 END VSS

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.66 0.46 5.91 0.6 ;
 RECT 5.56 0.32 5.91 0.46 ;
 RECT 3.66 0.235 3.8 0.46 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END RSTB

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.845 2.27 8.12 2.62 ;
 RECT 7.885 1.31 8.025 2.27 ;
 RECT 7.885 1.17 8.975 1.31 ;
 RECT 8.835 1.31 8.975 2.615 ;
 RECT 7.885 0.86 8.025 1.17 ;
 RECT 7.83 0.72 8.06 0.86 ;
 RECT 8.78 0.72 9.03 0.86 ;
 RECT 8.835 0.86 8.975 1.17 ;
 END
 ANTENNADIFFAREA 1.02 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.205 2.26 10.53 2.59 ;
 RECT 10.205 1.6 10.345 2.26 ;
 RECT 9.255 1.46 10.345 1.6 ;
 RECT 9.255 1.6 9.395 2.605 ;
 RECT 10.205 0.445 10.345 1.46 ;
 RECT 9.195 0.765 9.445 0.905 ;
 RECT 9.255 0.905 9.395 1.46 ;
 END
 ANTENNADIFFAREA 0.977 ;
 END QN

 OBS
 LAYER PO ;
 RECT 6.815 0.525 6.915 2.585 ;
 RECT 5.035 2.455 5.265 2.585 ;
 RECT 5.035 2.585 6.915 2.685 ;
 RECT 3.175 0.595 3.275 1.095 ;
 RECT 2.97 1.095 3.275 1.195 ;
 RECT 4.5 0.61 4.6 1.55 ;
 RECT 2.97 1.195 3.07 1.58 ;
 RECT 3.815 1.55 4.6 1.65 ;
 RECT 2.8 1.58 3.07 1.81 ;
 RECT 3.815 1.65 3.915 2.485 ;
 RECT 2.97 1.81 3.07 2.485 ;
 RECT 2.97 2.485 3.915 2.585 ;
 RECT 3.615 0.235 3.845 0.315 ;
 RECT 3.615 0.415 3.845 0.465 ;
 RECT 1.485 0.315 3.845 0.415 ;
 RECT 1.485 0.415 1.585 1.305 ;
 RECT 1.485 1.305 1.755 1.405 ;
 RECT 1.655 1.405 1.755 2.39 ;
 RECT 3.535 1.22 3.755 1.37 ;
 RECT 3.535 1.12 4.13 1.22 ;
 RECT 4.03 0.43 4.13 1.12 ;
 RECT 4.03 0.33 5.07 0.43 ;
 RECT 4.97 0.43 5.07 1.835 ;
 RECT 4.285 1.835 5.07 1.935 ;
 RECT 4.285 1.935 4.385 2.48 ;
 RECT 9.99 0.29 10.09 1.115 ;
 RECT 9.795 1.115 10.09 1.345 ;
 RECT 9.51 0.255 9.61 2.67 ;
 RECT 9.99 1.345 10.09 2.67 ;
 RECT 9.51 2.67 10.09 2.77 ;
 RECT 6.28 0.255 6.515 0.42 ;
 RECT 6.28 0.155 8.24 0.255 ;
 RECT 8.62 0.195 8.72 1.02 ;
 RECT 8.14 0.255 8.24 1.02 ;
 RECT 8.62 1.255 8.72 2.775 ;
 RECT 8.14 1.02 8.72 1.255 ;
 RECT 8.14 1.255 8.24 2.775 ;
 RECT 1.185 0.615 1.285 1.33 ;
 RECT 1.03 1.33 1.285 1.575 ;
 RECT 1.185 1.575 1.285 2.39 ;
 RECT 2.33 0.595 2.43 1.18 ;
 RECT 2.125 1.18 2.43 1.41 ;
 RECT 2.125 1.41 2.225 2.375 ;
 RECT 5.97 0.615 6.07 1.14 ;
 RECT 5.97 1.14 6.47 1.37 ;
 RECT 5.97 1.37 6.07 2.385 ;
 RECT 7.285 0.52 7.385 1.155 ;
 RECT 7.095 1.155 7.385 1.385 ;
 RECT 7.285 1.385 7.385 2.35 ;
 RECT 5.5 0.365 5.79 0.6 ;
 RECT 5.575 0.355 5.79 0.365 ;
 RECT 5.5 0.6 5.6 2.385 ;
 LAYER CO ;
 RECT 8.84 0.725 8.97 0.855 ;
 RECT 8.37 2.39 8.5 2.52 ;
 RECT 9.26 2.39 9.39 2.52 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 4.505 2.125 4.635 2.255 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 3.78 0.835 3.91 0.965 ;
 RECT 3.565 1.995 3.695 2.125 ;
 RECT 4.035 2.125 4.165 2.255 ;
 RECT 2.71 2.61 2.84 2.74 ;
 RECT 1.89 2.64 2.02 2.77 ;
 RECT 2.22 1.23 2.35 1.36 ;
 RECT 2.86 1.63 2.99 1.76 ;
 RECT 2.92 0.835 3.05 0.965 ;
 RECT 3.19 2.035 3.32 2.165 ;
 RECT 2.55 0.835 2.68 0.965 ;
 RECT 2.345 2.005 2.475 2.135 ;
 RECT 1.405 1.995 1.535 2.125 ;
 RECT 0.935 0.835 1.065 0.965 ;
 RECT 0.935 1.995 1.065 2.125 ;
 RECT 7.89 1.87 8.02 2 ;
 RECT 8.84 1.61 8.97 1.74 ;
 RECT 10.21 0.77 10.34 0.9 ;
 RECT 1.705 0.835 1.835 0.965 ;
 RECT 9.845 1.165 9.975 1.295 ;
 RECT 9.26 1.61 9.39 1.74 ;
 RECT 9.26 1.87 9.39 2 ;
 RECT 10.21 0.51 10.34 0.64 ;
 RECT 10.21 2.39 10.34 2.52 ;
 RECT 9.26 2.13 9.39 2.26 ;
 RECT 9.74 2.13 9.87 2.26 ;
 RECT 1.08 1.385 1.21 1.515 ;
 RECT 6.29 1.19 6.42 1.32 ;
 RECT 7.89 1.61 8.02 1.74 ;
 RECT 8.37 2.13 8.5 2.26 ;
 RECT 7.88 0.725 8.01 0.855 ;
 RECT 9.74 2.39 9.87 2.52 ;
 RECT 9.26 1.61 9.39 1.74 ;
 RECT 9.74 2.13 9.87 2.26 ;
 RECT 9.26 0.77 9.39 0.9 ;
 RECT 9.26 1.87 9.39 2 ;
 RECT 10.21 1.61 10.34 1.74 ;
 RECT 9.26 2.13 9.39 2.26 ;
 RECT 9.74 2.39 9.87 2.52 ;
 RECT 10.21 1.87 10.34 2 ;
 RECT 10.21 2.13 10.34 2.26 ;
 RECT 9.73 0.115 9.86 0.245 ;
 RECT 9.74 1.87 9.87 2 ;
 RECT 9.26 2.39 9.39 2.52 ;
 RECT 4.25 0.835 4.38 0.965 ;
 RECT 4.72 0.835 4.85 0.965 ;
 RECT 7.505 1.99 7.635 2.12 ;
 RECT 6.565 1.99 6.695 2.12 ;
 RECT 7.035 1.975 7.165 2.105 ;
 RECT 7.505 0.745 7.635 0.875 ;
 RECT 6.19 1.99 6.32 2.12 ;
 RECT 5.25 1.99 5.38 2.12 ;
 RECT 5.61 0.405 5.74 0.535 ;
 RECT 5.72 1.99 5.85 2.12 ;
 RECT 6.19 0.835 6.32 0.965 ;
 RECT 5.24 0.125 5.37 0.255 ;
 RECT 7.89 2.13 8.02 2.26 ;
 RECT 8.37 2.39 8.5 2.52 ;
 RECT 8.84 1.87 8.97 2 ;
 RECT 8.84 2.13 8.97 2.26 ;
 RECT 8.36 0.11 8.49 0.24 ;
 RECT 8.37 1.87 8.5 2 ;
 RECT 7.89 2.39 8.02 2.52 ;
 RECT 3.665 0.285 3.795 0.415 ;
 RECT 5.085 2.505 5.215 2.635 ;
 RECT 3.395 0.835 3.525 0.965 ;
 RECT 6.335 0.24 6.465 0.37 ;
 RECT 6.56 0.745 6.69 0.875 ;
 RECT 2.075 0.835 2.205 0.965 ;
 RECT 3.575 1.19 3.705 1.32 ;
 RECT 7.145 1.205 7.275 1.335 ;
 RECT 8.37 1.61 8.5 1.74 ;
 RECT 7.89 1.61 8.02 1.74 ;
 RECT 7.89 1.87 8.02 2 ;
 RECT 8.84 2.39 8.97 2.52 ;
 RECT 7.89 2.13 8.02 2.26 ;
 RECT 8.37 2.13 8.5 2.26 ;
 RECT 7.89 2.39 8.02 2.52 ;
 LAYER M1 ;
 RECT 6.19 1.185 6.7 1.325 ;
 RECT 6.56 1.325 6.7 1.565 ;
 RECT 6.56 1.705 6.7 1.985 ;
 RECT 6.515 1.985 6.745 2.125 ;
 RECT 7.455 1.985 7.685 2.125 ;
 RECT 7.5 0.575 7.64 1.565 ;
 RECT 7.5 1.705 7.64 1.985 ;
 RECT 6.56 1.565 7.64 1.705 ;
 RECT 9.775 1.16 10.06 1.3 ;
 RECT 9.775 0.575 9.915 1.16 ;
 RECT 7.5 0.435 9.915 0.575 ;
 RECT 5.2 1.985 5.43 2.125 ;
 RECT 5.245 1.69 5.385 1.985 ;
 RECT 4.715 0.78 4.855 1.16 ;
 RECT 4.5 1.3 4.64 2.12 ;
 RECT 4.41 2.12 4.695 2.26 ;
 RECT 6.14 1.985 6.37 2.125 ;
 RECT 6.23 0.375 6.37 0.83 ;
 RECT 6.185 1.69 6.325 1.985 ;
 RECT 5.715 0.83 6.37 0.97 ;
 RECT 5.24 1.55 6.325 1.69 ;
 RECT 5.715 0.97 5.855 1.16 ;
 RECT 5.715 1.3 5.855 1.55 ;
 RECT 4.5 1.16 5.855 1.3 ;
 RECT 6.23 0.235 6.515 0.375 ;
 RECT 4.22 0.77 4.39 1.02 ;
 RECT 4.22 1.02 4.36 1.775 ;
 RECT 4.03 1.775 4.36 1.915 ;
 RECT 4.03 1.915 4.17 2.5 ;
 RECT 4.03 2.5 5.265 2.64 ;
 RECT 2.915 0.775 3.055 1.185 ;
 RECT 3.185 1.325 3.325 2.03 ;
 RECT 3.185 2.17 3.325 2.185 ;
 RECT 3.1 2.03 3.37 2.17 ;
 RECT 2.915 1.185 3.755 1.325 ;
 RECT 2.545 0.785 2.685 1.625 ;
 RECT 2.34 1.625 3.045 1.765 ;
 RECT 2.34 1.765 2.48 2 ;
 RECT 2.295 2 2.525 2.14 ;
 RECT 2.34 2.14 2.48 2.175 ;
 RECT 1.7 0.785 1.84 1.99 ;
 RECT 1.31 1.99 1.84 2.13 ;
 RECT 1.4 2.13 1.54 2.325 ;
 RECT 3.73 0.83 4.08 0.97 ;
 RECT 3.94 0.97 4.08 1.465 ;
 RECT 3.56 1.465 4.08 1.605 ;
 RECT 3.56 1.605 3.7 2.325 ;
 RECT 1.4 2.325 3.7 2.465 ;
 END
END LASRX2

MACRO LASX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.64 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.995 0.24 1.285 0.615 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.52 1.16 1.92 1.45 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.06 2.28 7.335 2.55 ;
 RECT 7.12 0.86 7.26 2.28 ;
 RECT 7.065 0.72 7.295 0.86 ;
 END
 ANTENNADIFFAREA 0.527 ;
 END Q

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.415 2.265 6.705 2.53 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END SETB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.64 2.96 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 6.065 1.97 6.46 2.11 ;
 RECT 7.6 1.495 7.74 2.8 ;
 RECT 4.7 1.9 4.84 2.8 ;
 RECT 2.175 2.605 2.405 2.8 ;
 RECT 1.355 2.63 1.585 2.8 ;
 RECT 6.065 2.11 6.205 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.64 0.08 ;
 RECT 0.34 0.08 0.48 0.81 ;
 RECT 7.545 0.08 7.775 0.275 ;
 RECT 5.78 0.735 6.37 0.875 ;
 RECT 5.125 0.83 5.355 0.97 ;
 RECT 1.49 0.705 1.885 0.845 ;
 RECT 2.905 0.08 3.045 1.03 ;
 RECT 5.78 0.875 5.92 0.93 ;
 RECT 5.78 0.685 5.92 0.735 ;
 RECT 6.23 0.08 6.37 0.735 ;
 RECT 5.17 0.08 5.31 0.83 ;
 RECT 1.49 0.845 1.63 1.015 ;
 RECT 1.745 0.08 1.885 0.705 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.015 2.06 8.29 2.395 ;
 RECT 8.07 0.565 8.21 2.06 ;
 END
 ANTENNADIFFAREA 0.454 ;
 END QN

 OBS
 LAYER PO ;
 RECT 1.845 0.575 1.945 1.18 ;
 RECT 1.525 1.18 1.945 1.41 ;
 RECT 1.64 1.41 1.74 2.405 ;
 RECT 2.69 0.575 2.79 1.095 ;
 RECT 2.485 1.195 2.585 1.58 ;
 RECT 2.485 1.095 2.79 1.195 ;
 RECT 4.015 0.61 4.115 1.55 ;
 RECT 3.33 1.55 4.115 1.65 ;
 RECT 2.315 1.58 2.585 1.81 ;
 RECT 3.33 1.65 3.43 2.485 ;
 RECT 2.485 1.81 2.585 2.485 ;
 RECT 2.485 2.485 3.43 2.585 ;
 RECT 5.51 0.255 5.74 0.42 ;
 RECT 5.51 0.155 7.475 0.255 ;
 RECT 7.375 0.255 7.475 2.77 ;
 RECT 7.855 0.305 7.955 1.02 ;
 RECT 7.69 1.02 7.955 1.255 ;
 RECT 7.855 1.255 7.955 2.775 ;
 RECT 1.005 0.24 1.285 0.47 ;
 RECT 1.185 0.47 1.285 2.485 ;
 RECT 3.05 1.22 3.27 1.37 ;
 RECT 3.05 1.12 3.645 1.22 ;
 RECT 3.545 0.43 3.645 1.12 ;
 RECT 3.545 0.33 4.585 0.43 ;
 RECT 4.485 0.43 4.585 1.835 ;
 RECT 3.8 1.835 4.585 1.935 ;
 RECT 3.8 1.935 3.9 2.48 ;
 RECT 6.51 0.51 6.61 2.27 ;
 RECT 6.415 2.27 6.635 2.5 ;
 RECT 6.04 0.515 6.14 2.685 ;
 RECT 4.275 2.455 4.505 2.685 ;
 RECT 4.275 2.685 6.14 2.785 ;
 RECT 4.955 0.615 5.055 2.335 ;
 RECT 5.45 2.275 5.68 2.335 ;
 RECT 5.45 2.435 5.68 2.505 ;
 RECT 4.955 2.335 5.68 2.435 ;
 LAYER CO ;
 RECT 7.125 1.895 7.255 2.025 ;
 RECT 7.125 2.155 7.255 2.285 ;
 RECT 6.465 2.32 6.595 2.45 ;
 RECT 6.73 1.99 6.86 2.12 ;
 RECT 5.79 1.99 5.92 2.12 ;
 RECT 6.26 1.975 6.39 2.105 ;
 RECT 6.73 0.74 6.86 0.87 ;
 RECT 5.175 1.99 5.305 2.12 ;
 RECT 4.705 1.99 4.835 2.12 ;
 RECT 5.175 0.835 5.305 0.965 ;
 RECT 0.93 0.835 1.06 0.965 ;
 RECT 4.705 0.835 4.835 0.965 ;
 RECT 1.055 0.29 1.185 0.42 ;
 RECT 4.325 2.505 4.455 2.635 ;
 RECT 2.91 0.835 3.04 0.965 ;
 RECT 5.56 0.24 5.69 0.37 ;
 RECT 5.785 0.74 5.915 0.87 ;
 RECT 7.595 0.11 7.725 0.24 ;
 RECT 7.74 1.07 7.87 1.2 ;
 RECT 8.075 0.635 8.205 0.765 ;
 RECT 7.605 2.155 7.735 2.285 ;
 RECT 8.075 1.635 8.205 1.765 ;
 RECT 7.605 2.415 7.735 2.545 ;
 RECT 8.075 1.895 8.205 2.025 ;
 RECT 8.075 2.155 8.205 2.285 ;
 RECT 7.605 1.895 7.735 2.025 ;
 RECT 7.605 2.155 7.735 2.285 ;
 RECT 7.115 0.725 7.245 0.855 ;
 RECT 1.495 0.835 1.625 0.965 ;
 RECT 3.09 1.19 3.22 1.32 ;
 RECT 3.765 0.835 3.895 0.965 ;
 RECT 4.235 0.835 4.365 0.965 ;
 RECT 4.02 2.125 4.15 2.255 ;
 RECT 3.765 0.835 3.895 0.965 ;
 RECT 3.295 0.835 3.425 0.965 ;
 RECT 3.08 1.995 3.21 2.125 ;
 RECT 3.55 2.125 3.68 2.255 ;
 RECT 2.225 2.61 2.355 2.74 ;
 RECT 1.405 2.64 1.535 2.77 ;
 RECT 1.575 1.23 1.705 1.36 ;
 RECT 2.375 1.63 2.505 1.76 ;
 RECT 2.435 0.835 2.565 0.965 ;
 RECT 2.705 2.035 2.835 2.165 ;
 RECT 2.065 0.835 2.195 0.965 ;
 RECT 1.86 2.005 1.99 2.135 ;
 RECT 0.93 2.11 1.06 2.24 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 5.5 2.325 5.63 2.455 ;
 RECT 7.605 1.635 7.735 1.765 ;
 RECT 7.125 1.635 7.255 1.765 ;
 RECT 7.125 1.895 7.255 2.025 ;
 RECT 7.125 2.155 7.255 2.285 ;
 RECT 7.125 1.635 7.255 1.765 ;
 LAYER M1 ;
 RECT 3.735 0.77 3.905 1.02 ;
 RECT 3.735 1.02 3.875 1.775 ;
 RECT 3.545 1.775 3.875 1.915 ;
 RECT 3.545 1.915 3.685 2.5 ;
 RECT 3.545 2.5 4.505 2.64 ;
 RECT 2.7 1.325 2.84 2.03 ;
 RECT 2.7 2.17 2.84 2.185 ;
 RECT 2.43 0.775 2.57 1.185 ;
 RECT 2.615 2.03 2.885 2.17 ;
 RECT 2.43 1.185 3.27 1.325 ;
 RECT 2.06 0.785 2.2 1.625 ;
 RECT 1.855 1.625 2.56 1.765 ;
 RECT 1.855 1.765 1.995 2 ;
 RECT 1.81 2 2.04 2.14 ;
 RECT 1.855 2.14 1.995 2.175 ;
 RECT 0.925 0.775 1.065 2.325 ;
 RECT 0.925 2.325 3.215 2.465 ;
 RECT 3.245 0.83 3.595 0.97 ;
 RECT 3.455 0.97 3.595 1.465 ;
 RECT 3.075 1.465 3.595 1.605 ;
 RECT 3.075 1.605 3.215 2.325 ;
 RECT 5.785 1.675 5.925 2.32 ;
 RECT 5.45 2.32 5.925 2.46 ;
 RECT 6.68 1.985 6.91 2.125 ;
 RECT 6.725 0.575 6.865 1.535 ;
 RECT 6.725 1.675 6.865 1.985 ;
 RECT 5.785 1.535 6.865 1.675 ;
 RECT 7.57 1.065 7.92 1.205 ;
 RECT 7.57 0.575 7.71 1.065 ;
 RECT 6.725 0.435 7.71 0.575 ;
 RECT 4.23 0.78 4.37 1.61 ;
 RECT 4.015 1.75 4.155 2.12 ;
 RECT 3.925 2.12 4.21 2.26 ;
 RECT 4.7 0.78 4.84 1.11 ;
 RECT 4.7 1.25 4.84 1.61 ;
 RECT 5.5 0.235 5.74 0.375 ;
 RECT 5.5 0.375 5.64 1.11 ;
 RECT 5.17 1.75 5.31 2.195 ;
 RECT 4.695 1.11 5.64 1.25 ;
 RECT 4.015 1.61 5.31 1.75 ;
 END
END LASX1

MACRO LASX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.92 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.01 0.225 1.285 0.61 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.38 1.16 1.92 1.45 ;
 END
 ANTENNAGATEAREA 0.05 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.06 2.29 7.33 2.54 ;
 RECT 7.065 0.72 7.295 0.86 ;
 RECT 7.12 1.23 8.21 1.37 ;
 RECT 8.025 0.735 8.255 0.875 ;
 RECT 7.12 1.37 7.26 2.29 ;
 RECT 7.12 0.86 7.26 1.23 ;
 RECT 8.07 1.37 8.21 2.61 ;
 RECT 8.07 0.875 8.21 1.23 ;
 END
 ANTENNADIFFAREA 1.008 ;
 END Q

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.395 2.265 6.705 2.535 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END SETB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.92 2.96 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 6.065 1.97 6.46 2.11 ;
 RECT 8.93 1.78 9.07 2.8 ;
 RECT 4.7 1.9 4.84 2.8 ;
 RECT 2.175 2.605 2.405 2.8 ;
 RECT 1.355 2.63 1.585 2.8 ;
 RECT 7.6 1.74 7.74 2.8 ;
 RECT 6.065 2.11 6.205 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.92 0.08 ;
 RECT 0.34 0.08 0.48 0.81 ;
 RECT 7.545 0.08 7.775 0.275 ;
 RECT 8.875 0.08 9.105 0.27 ;
 RECT 5.78 0.715 6.37 0.855 ;
 RECT 5.125 0.83 5.355 0.97 ;
 RECT 1.49 0.705 1.885 0.845 ;
 RECT 2.905 0.08 3.045 1.03 ;
 RECT 5.78 0.855 5.92 0.91 ;
 RECT 5.78 0.665 5.92 0.715 ;
 RECT 6.23 0.08 6.37 0.715 ;
 RECT 5.17 0.08 5.31 0.83 ;
 RECT 1.49 0.845 1.63 1.015 ;
 RECT 1.745 0.08 1.885 0.705 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.32 2.12 9.56 2.36 ;
 RECT 8.45 1.425 9.54 1.565 ;
 RECT 8.395 0.72 8.625 0.86 ;
 RECT 9.4 1.565 9.54 2.12 ;
 RECT 8.45 1.565 8.59 2.455 ;
 RECT 8.45 0.86 8.59 1.425 ;
 RECT 9.4 0.565 9.54 1.425 ;
 END
 ANTENNADIFFAREA 0.953 ;
 END QN

 OBS
 LAYER PO ;
 RECT 6.51 0.45 6.61 2.26 ;
 RECT 6.45 2.26 6.705 2.49 ;
 RECT 8.705 0.155 8.805 1.1 ;
 RECT 8.705 1.2 8.805 2.74 ;
 RECT 9.02 1.02 9.285 1.1 ;
 RECT 9.02 1.2 9.285 1.255 ;
 RECT 8.705 1.1 9.285 1.2 ;
 RECT 9.185 0.14 9.285 1.02 ;
 RECT 9.185 1.255 9.285 2.74 ;
 RECT 6.04 0.45 6.14 2.685 ;
 RECT 4.275 2.455 4.505 2.685 ;
 RECT 4.275 2.685 6.14 2.785 ;
 RECT 1.185 0.47 1.285 2.51 ;
 RECT 1.02 0.24 1.285 0.47 ;
 RECT 1.845 0.575 1.945 1.18 ;
 RECT 1.525 1.18 1.945 1.41 ;
 RECT 1.64 1.41 1.74 2.405 ;
 RECT 3.05 1.22 3.27 1.37 ;
 RECT 3.05 1.12 3.645 1.22 ;
 RECT 3.545 0.43 3.645 1.12 ;
 RECT 3.545 0.33 4.585 0.43 ;
 RECT 4.485 0.43 4.585 1.835 ;
 RECT 3.8 1.835 4.585 1.935 ;
 RECT 3.8 1.935 3.9 2.48 ;
 RECT 4.955 0.615 5.055 2.335 ;
 RECT 5.45 2.275 5.68 2.335 ;
 RECT 5.45 2.435 5.68 2.505 ;
 RECT 4.955 2.335 5.68 2.435 ;
 RECT 2.69 0.575 2.79 1.095 ;
 RECT 2.485 1.195 2.585 1.58 ;
 RECT 2.485 1.095 2.79 1.195 ;
 RECT 4.015 0.61 4.115 1.55 ;
 RECT 3.33 1.55 4.115 1.65 ;
 RECT 2.315 1.58 2.585 1.81 ;
 RECT 3.33 1.65 3.43 2.485 ;
 RECT 2.485 1.81 2.585 2.485 ;
 RECT 2.485 2.485 3.43 2.585 ;
 RECT 7.855 0.14 7.955 1.025 ;
 RECT 7.855 1.125 7.955 2.725 ;
 RECT 5.51 0.255 5.74 0.42 ;
 RECT 7.375 0.255 7.475 1.025 ;
 RECT 7.375 1.125 7.475 2.725 ;
 RECT 7.375 1.025 7.955 1.125 ;
 RECT 5.51 0.155 7.475 0.255 ;
 LAYER CO ;
 RECT 7.125 2.155 7.255 2.285 ;
 RECT 0.93 2.11 1.06 2.24 ;
 RECT 7.125 1.635 7.255 1.765 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 4.705 1.99 4.835 2.12 ;
 RECT 5.175 0.835 5.305 0.965 ;
 RECT 5.495 2.325 5.625 2.455 ;
 RECT 6.505 2.31 6.635 2.44 ;
 RECT 6.73 1.99 6.86 2.12 ;
 RECT 5.79 1.99 5.92 2.12 ;
 RECT 6.26 1.975 6.39 2.105 ;
 RECT 8.455 2.155 8.585 2.285 ;
 RECT 8.455 1.635 8.585 1.765 ;
 RECT 8.445 0.725 8.575 0.855 ;
 RECT 9.405 1.635 9.535 1.765 ;
 RECT 9.405 0.635 9.535 0.765 ;
 RECT 0.93 0.835 1.06 0.965 ;
 RECT 4.705 0.835 4.835 0.965 ;
 RECT 5.785 0.72 5.915 0.85 ;
 RECT 7.595 0.11 7.725 0.24 ;
 RECT 8.075 0.745 8.205 0.875 ;
 RECT 7.605 2.155 7.735 2.285 ;
 RECT 8.075 1.635 8.205 1.765 ;
 RECT 1.495 0.835 1.625 0.965 ;
 RECT 3.09 1.19 3.22 1.32 ;
 RECT 3.765 0.835 3.895 0.965 ;
 RECT 4.235 0.835 4.365 0.965 ;
 RECT 4.02 2.125 4.15 2.255 ;
 RECT 1.575 1.23 1.705 1.36 ;
 RECT 2.375 1.63 2.505 1.76 ;
 RECT 2.435 0.835 2.565 0.965 ;
 RECT 2.705 2.035 2.835 2.165 ;
 RECT 2.065 0.835 2.195 0.965 ;
 RECT 1.86 2.005 1.99 2.135 ;
 RECT 7.125 1.895 7.255 2.025 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 6.73 0.72 6.86 0.85 ;
 RECT 5.175 1.945 5.305 2.075 ;
 RECT 4.325 2.505 4.455 2.635 ;
 RECT 8.455 1.635 8.585 1.765 ;
 RECT 8.925 0.11 9.055 0.24 ;
 RECT 8.455 2.155 8.585 2.285 ;
 RECT 8.455 1.895 8.585 2.025 ;
 RECT 8.935 2.155 9.065 2.285 ;
 RECT 9.405 2.155 9.535 2.285 ;
 RECT 9.07 1.07 9.2 1.2 ;
 RECT 8.935 2.155 9.065 2.285 ;
 RECT 9.405 1.895 9.535 2.025 ;
 RECT 8.455 1.895 8.585 2.025 ;
 RECT 8.935 1.895 9.065 2.025 ;
 RECT 1.07 0.29 1.2 0.42 ;
 RECT 2.91 0.835 3.04 0.965 ;
 RECT 5.56 0.24 5.69 0.37 ;
 RECT 8.075 1.895 8.205 2.025 ;
 RECT 8.075 2.155 8.205 2.285 ;
 RECT 7.605 1.895 7.735 2.025 ;
 RECT 7.605 2.155 7.735 2.285 ;
 RECT 7.115 0.725 7.245 0.855 ;
 RECT 3.765 0.835 3.895 0.965 ;
 RECT 3.295 0.835 3.425 0.965 ;
 RECT 3.08 1.995 3.21 2.125 ;
 RECT 3.55 2.125 3.68 2.255 ;
 RECT 2.225 2.61 2.355 2.74 ;
 RECT 1.405 2.64 1.535 2.77 ;
 RECT 7.125 2.155 7.255 2.285 ;
 RECT 7.125 1.635 7.255 1.765 ;
 RECT 7.125 1.895 7.255 2.025 ;
 LAYER M1 ;
 RECT 3.735 0.77 3.905 1.02 ;
 RECT 3.735 1.02 3.875 1.775 ;
 RECT 3.545 1.775 3.875 1.915 ;
 RECT 3.545 1.915 3.685 2.5 ;
 RECT 3.545 2.5 4.505 2.64 ;
 RECT 2.7 1.325 2.84 2.03 ;
 RECT 2.7 2.17 2.84 2.185 ;
 RECT 2.43 0.775 2.57 1.185 ;
 RECT 2.615 2.03 2.885 2.17 ;
 RECT 2.43 1.185 3.27 1.325 ;
 RECT 2.06 0.785 2.2 1.625 ;
 RECT 1.855 1.625 2.56 1.765 ;
 RECT 1.855 1.765 1.995 2 ;
 RECT 1.81 2 2.04 2.14 ;
 RECT 1.855 2.14 1.995 2.175 ;
 RECT 0.925 0.775 1.065 2.325 ;
 RECT 0.925 2.325 3.215 2.465 ;
 RECT 3.245 0.83 3.595 0.97 ;
 RECT 3.455 0.97 3.595 1.465 ;
 RECT 3.075 1.465 3.595 1.605 ;
 RECT 3.075 1.605 3.215 2.325 ;
 RECT 5.785 1.675 5.925 2.32 ;
 RECT 5.49 2.32 5.925 2.46 ;
 RECT 5.49 2.255 5.63 2.32 ;
 RECT 5.49 2.46 5.63 2.525 ;
 RECT 6.68 1.985 6.91 2.125 ;
 RECT 6.725 0.575 6.865 1.535 ;
 RECT 6.725 1.675 6.865 1.985 ;
 RECT 5.785 1.535 6.865 1.675 ;
 RECT 9.065 0.575 9.205 1.26 ;
 RECT 6.725 0.435 9.205 0.575 ;
 RECT 4.23 0.78 4.37 1.61 ;
 RECT 4.015 1.75 4.155 2.12 ;
 RECT 3.925 2.12 4.21 2.26 ;
 RECT 4.7 0.78 4.84 1.11 ;
 RECT 4.7 1.25 4.84 1.61 ;
 RECT 5.5 0.235 5.74 0.375 ;
 RECT 5.5 0.375 5.64 1.11 ;
 RECT 5.17 1.75 5.31 2.145 ;
 RECT 4.7 1.11 5.64 1.25 ;
 RECT 4.015 1.61 5.31 1.75 ;
 END
END LASX2

MACRO LATCHX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.68 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.68 2.96 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 6.64 1.495 6.78 2.8 ;
 RECT 5.17 1.9 5.31 2.8 ;
 RECT 2.175 2.605 2.405 2.8 ;
 RECT 1.355 2.63 1.585 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.68 0.08 ;
 RECT 0.345 0.08 0.485 0.81 ;
 RECT 6.585 0.08 6.815 0.275 ;
 RECT 1.49 0.705 1.885 0.845 ;
 RECT 5.175 0.08 5.315 0.955 ;
 RECT 2.905 0.08 3.045 1.03 ;
 RECT 1.49 0.845 1.63 1.015 ;
 RECT 1.745 0.08 1.885 0.705 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 0.36 1.285 0.63 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.52 1.16 1.92 1.45 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.1 2.32 6.36 2.56 ;
 RECT 6.16 0.86 6.3 2.32 ;
 RECT 6.105 0.72 6.335 0.86 ;
 END
 ANTENNADIFFAREA 0.517 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.055 2.06 7.41 2.395 ;
 RECT 7.11 0.565 7.25 2.06 ;
 END
 ANTENNADIFFAREA 0.533 ;
 END QN

 OBS
 LAYER PO ;
 RECT 1.845 0.575 1.945 1.18 ;
 RECT 1.525 1.18 1.945 1.41 ;
 RECT 1.64 1.41 1.74 2.405 ;
 RECT 2.69 0.575 2.79 1.095 ;
 RECT 2.485 1.195 2.585 1.58 ;
 RECT 2.485 1.095 2.79 1.195 ;
 RECT 4.015 0.61 4.115 1.55 ;
 RECT 3.33 1.55 4.115 1.65 ;
 RECT 2.315 1.58 2.585 1.81 ;
 RECT 3.33 1.65 3.43 2.485 ;
 RECT 2.485 1.81 2.585 2.485 ;
 RECT 2.485 2.485 3.43 2.585 ;
 RECT 6.895 0.115 6.995 1.02 ;
 RECT 6.73 1.02 6.995 1.255 ;
 RECT 6.895 1.255 6.995 2.745 ;
 RECT 4.955 0.5 5.055 1.24 ;
 RECT 4.955 1.24 5.18 1.47 ;
 RECT 4.955 1.47 5.055 2.385 ;
 RECT 3.05 1.22 3.27 1.37 ;
 RECT 3.05 1.12 3.645 1.22 ;
 RECT 3.545 0.43 3.645 1.12 ;
 RECT 3.545 0.33 4.585 0.43 ;
 RECT 4.485 0.43 4.585 1.835 ;
 RECT 3.8 1.835 4.585 1.935 ;
 RECT 3.8 1.935 3.9 2.48 ;
 RECT 5.43 0.5 5.53 2.685 ;
 RECT 6.415 0.105 6.515 2.685 ;
 RECT 4.275 2.455 4.505 2.685 ;
 RECT 4.275 2.685 6.515 2.785 ;
 RECT 1.025 0.39 1.285 0.6 ;
 RECT 1.185 0.6 1.285 2.655 ;
 LAYER CO ;
 RECT 6.645 1.635 6.775 1.765 ;
 RECT 6.165 1.895 6.295 2.025 ;
 RECT 6.165 2.155 6.295 2.285 ;
 RECT 6.165 1.895 6.295 2.025 ;
 RECT 6.165 2.155 6.295 2.285 ;
 RECT 5.685 2.03 5.815 2.16 ;
 RECT 5.685 0.74 5.815 0.87 ;
 RECT 5.175 1.99 5.305 2.12 ;
 RECT 4.705 2.03 4.835 2.16 ;
 RECT 5.18 0.74 5.31 0.87 ;
 RECT 5 1.29 5.13 1.42 ;
 RECT 0.93 0.835 1.06 0.965 ;
 RECT 4.705 0.74 4.835 0.87 ;
 RECT 4.325 2.505 4.455 2.635 ;
 RECT 2.91 0.835 3.04 0.965 ;
 RECT 6.635 0.11 6.765 0.24 ;
 RECT 6.78 1.07 6.91 1.2 ;
 RECT 7.115 0.635 7.245 0.765 ;
 RECT 6.645 2.155 6.775 2.285 ;
 RECT 7.115 1.635 7.245 1.765 ;
 RECT 7.115 1.895 7.245 2.025 ;
 RECT 7.115 2.155 7.245 2.285 ;
 RECT 6.645 1.895 6.775 2.025 ;
 RECT 6.645 2.155 6.775 2.285 ;
 RECT 6.155 0.725 6.285 0.855 ;
 RECT 1.495 0.835 1.625 0.965 ;
 RECT 3.09 1.19 3.22 1.32 ;
 RECT 3.765 0.835 3.895 0.965 ;
 RECT 4.235 0.835 4.365 0.965 ;
 RECT 4.02 2.125 4.15 2.255 ;
 RECT 3.765 0.835 3.895 0.965 ;
 RECT 3.295 0.835 3.425 0.965 ;
 RECT 3.08 1.995 3.21 2.125 ;
 RECT 3.55 2.125 3.68 2.255 ;
 RECT 2.225 2.61 2.355 2.74 ;
 RECT 1.405 2.64 1.535 2.77 ;
 RECT 1.575 1.23 1.705 1.36 ;
 RECT 2.375 1.63 2.505 1.76 ;
 RECT 2.435 0.835 2.565 0.965 ;
 RECT 2.705 2.035 2.835 2.165 ;
 RECT 2.065 0.835 2.195 0.965 ;
 RECT 1.86 2 1.99 2.13 ;
 RECT 0.93 2.11 1.06 2.24 ;
 RECT 0.35 0.605 0.48 0.735 ;
 RECT 0.35 0.345 0.48 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 1.075 0.43 1.205 0.56 ;
 LAYER M1 ;
 RECT 4.7 0.67 4.84 1.61 ;
 RECT 4.7 1.75 4.84 2.23 ;
 RECT 4.23 0.78 4.37 1.61 ;
 RECT 4.015 1.75 4.155 2.12 ;
 RECT 4.015 1.61 4.84 1.75 ;
 RECT 3.925 2.12 4.21 2.26 ;
 RECT 3.735 0.77 3.905 1.02 ;
 RECT 3.735 1.02 3.875 1.775 ;
 RECT 3.545 1.775 3.875 1.915 ;
 RECT 3.545 1.915 3.685 2.5 ;
 RECT 3.545 2.5 4.505 2.64 ;
 RECT 2.7 1.325 2.84 2.03 ;
 RECT 2.7 2.17 2.84 2.185 ;
 RECT 2.43 0.775 2.57 1.185 ;
 RECT 2.615 2.03 2.885 2.17 ;
 RECT 2.43 1.185 3.27 1.325 ;
 RECT 4.995 1.22 5.135 1.285 ;
 RECT 4.995 1.425 5.135 1.49 ;
 RECT 5.68 0.575 5.82 1.285 ;
 RECT 4.995 1.285 5.82 1.425 ;
 RECT 5.68 1.425 5.82 2.025 ;
 RECT 5.635 2.025 5.865 2.165 ;
 RECT 6.61 1.065 6.96 1.205 ;
 RECT 6.61 0.575 6.75 1.065 ;
 RECT 5.68 0.435 6.75 0.575 ;
 RECT 2.06 0.785 2.2 1.625 ;
 RECT 1.855 1.625 2.56 1.765 ;
 RECT 1.855 1.765 1.995 1.995 ;
 RECT 1.81 1.995 2.04 2.135 ;
 RECT 1.855 2.135 1.995 2.17 ;
 RECT 0.925 0.775 1.065 2.325 ;
 RECT 0.925 2.325 3.215 2.465 ;
 RECT 3.245 0.83 3.595 0.97 ;
 RECT 3.455 0.97 3.595 1.465 ;
 RECT 3.075 1.465 3.595 1.605 ;
 RECT 3.075 1.605 3.215 2.325 ;
 END
END LATCHX1

MACRO LATCHX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.96 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.96 2.96 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 6.64 1.76 6.78 2.8 ;
 RECT 5.17 1.9 5.31 2.8 ;
 RECT 2.175 2.605 2.405 2.8 ;
 RECT 1.355 2.63 1.585 2.8 ;
 RECT 7.99 1.78 8.13 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.96 0.08 ;
 RECT 0.345 0.08 0.485 0.81 ;
 RECT 6.585 0.08 6.815 0.275 ;
 RECT 7.925 0.08 8.185 0.285 ;
 RECT 1.49 0.705 1.885 0.845 ;
 RECT 5.175 0.08 5.315 0.955 ;
 RECT 2.905 0.08 3.045 1.03 ;
 RECT 1.49 0.845 1.63 1.015 ;
 RECT 1.745 0.08 1.885 0.705 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.98 0.24 1.285 0.625 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.52 1.16 1.92 1.45 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.1 2.28 6.36 2.55 ;
 RECT 6.105 0.72 6.335 0.86 ;
 RECT 6.16 1.415 7.25 1.555 ;
 RECT 7.045 0.74 7.315 0.88 ;
 RECT 6.16 1.555 6.3 2.28 ;
 RECT 6.16 0.86 6.3 1.415 ;
 RECT 7.11 1.555 7.25 2.61 ;
 RECT 7.11 0.88 7.25 1.415 ;
 RECT 7.11 0.735 7.25 0.74 ;
 END
 ANTENNADIFFAREA 0.946 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.35 2.06 8.66 2.395 ;
 RECT 7.51 1.47 8.6 1.61 ;
 RECT 7.455 0.72 7.685 0.86 ;
 RECT 8.46 1.61 8.6 2.06 ;
 RECT 7.51 1.61 7.65 2.66 ;
 RECT 7.51 0.86 7.65 1.47 ;
 RECT 8.46 0.565 8.6 1.47 ;
 END
 ANTENNADIFFAREA 0.968 ;
 END QN

 OBS
 LAYER PO ;
 RECT 8.08 1.02 8.345 1.085 ;
 RECT 7.765 1.085 8.345 1.185 ;
 RECT 8.08 1.185 8.345 1.255 ;
 RECT 7.765 0.14 7.865 1.085 ;
 RECT 7.765 1.185 7.865 2.755 ;
 RECT 8.245 0.14 8.345 1.02 ;
 RECT 8.245 1.255 8.345 2.755 ;
 RECT 1.845 0.575 1.945 1.18 ;
 RECT 1.525 1.18 1.945 1.41 ;
 RECT 1.64 1.41 1.74 2.405 ;
 RECT 2.69 0.575 2.79 1.095 ;
 RECT 2.485 1.195 2.585 1.58 ;
 RECT 2.485 1.095 2.79 1.195 ;
 RECT 4.015 0.61 4.115 1.55 ;
 RECT 3.33 1.55 4.115 1.65 ;
 RECT 2.315 1.58 2.585 1.81 ;
 RECT 3.33 1.65 3.43 2.485 ;
 RECT 2.485 1.81 2.585 2.485 ;
 RECT 2.485 2.485 3.43 2.585 ;
 RECT 5.43 0.5 5.53 2.685 ;
 RECT 6.415 0.105 6.515 1.015 ;
 RECT 6.415 1.115 6.515 2.685 ;
 RECT 6.895 0.105 6.995 1.015 ;
 RECT 6.895 1.115 6.995 2.755 ;
 RECT 4.275 2.685 6.515 2.785 ;
 RECT 4.275 2.455 4.505 2.685 ;
 RECT 6.415 1.015 6.995 1.115 ;
 RECT 0.985 0.24 1.285 0.47 ;
 RECT 1.185 0.47 1.285 2.67 ;
 RECT 4.955 0.5 5.055 1.24 ;
 RECT 4.955 1.24 5.18 1.47 ;
 RECT 4.955 1.47 5.055 2.385 ;
 RECT 3.05 1.22 3.27 1.37 ;
 RECT 3.05 1.12 3.645 1.22 ;
 RECT 3.545 0.43 3.645 1.12 ;
 RECT 3.545 0.33 4.585 0.43 ;
 RECT 4.485 0.43 4.585 1.835 ;
 RECT 3.8 1.835 4.585 1.935 ;
 RECT 3.8 1.935 3.9 2.48 ;
 LAYER CO ;
 RECT 5.18 0.74 5.31 0.87 ;
 RECT 7.515 1.61 7.645 1.74 ;
 RECT 7.995 1.895 8.125 2.025 ;
 RECT 7.985 0.11 8.115 0.24 ;
 RECT 7.995 2.155 8.125 2.285 ;
 RECT 7.505 0.725 7.635 0.855 ;
 RECT 7.515 1.895 7.645 2.025 ;
 RECT 7.515 1.895 7.645 2.025 ;
 RECT 8.13 1.07 8.26 1.2 ;
 RECT 8.465 1.635 8.595 1.765 ;
 RECT 7.515 2.155 7.645 2.285 ;
 RECT 7.995 2.155 8.125 2.285 ;
 RECT 8.465 2.155 8.595 2.285 ;
 RECT 7.515 2.155 7.645 2.285 ;
 RECT 8.465 1.895 8.595 2.025 ;
 RECT 8.465 0.635 8.595 0.765 ;
 RECT 5 1.29 5.13 1.42 ;
 RECT 0.93 0.835 1.06 0.965 ;
 RECT 4.705 0.74 4.835 0.87 ;
 RECT 1.035 0.29 1.165 0.42 ;
 RECT 4.325 2.505 4.455 2.635 ;
 RECT 2.91 0.835 3.04 0.965 ;
 RECT 6.635 0.11 6.765 0.24 ;
 RECT 7.115 0.745 7.245 0.875 ;
 RECT 6.645 2.155 6.775 2.285 ;
 RECT 7.115 1.895 7.245 2.025 ;
 RECT 7.115 2.155 7.245 2.285 ;
 RECT 6.645 1.895 6.775 2.025 ;
 RECT 6.645 2.155 6.775 2.285 ;
 RECT 6.155 0.725 6.285 0.855 ;
 RECT 1.495 0.835 1.625 0.965 ;
 RECT 3.09 1.19 3.22 1.32 ;
 RECT 3.765 0.835 3.895 0.965 ;
 RECT 4.235 0.835 4.365 0.965 ;
 RECT 4.02 2.125 4.15 2.255 ;
 RECT 3.765 0.835 3.895 0.965 ;
 RECT 3.295 0.835 3.425 0.965 ;
 RECT 3.08 1.995 3.21 2.125 ;
 RECT 3.55 2.125 3.68 2.255 ;
 RECT 2.225 2.61 2.355 2.74 ;
 RECT 1.405 2.64 1.535 2.77 ;
 RECT 1.575 1.23 1.705 1.36 ;
 RECT 2.375 1.63 2.505 1.76 ;
 RECT 2.435 0.835 2.565 0.965 ;
 RECT 2.705 2.035 2.835 2.165 ;
 RECT 2.065 0.835 2.195 0.965 ;
 RECT 1.86 2 1.99 2.13 ;
 RECT 0.93 2.11 1.06 2.24 ;
 RECT 0.35 0.605 0.48 0.735 ;
 RECT 0.35 0.345 0.48 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 6.165 1.895 6.295 2.025 ;
 RECT 6.165 2.155 6.295 2.285 ;
 RECT 6.165 1.895 6.295 2.025 ;
 RECT 6.165 2.155 6.295 2.285 ;
 RECT 5.685 2.03 5.815 2.16 ;
 RECT 5.685 0.74 5.815 0.87 ;
 RECT 5.175 1.99 5.305 2.12 ;
 RECT 4.705 2.03 4.835 2.16 ;
 LAYER M1 ;
 RECT 4.995 1.22 5.135 1.285 ;
 RECT 4.995 1.425 5.135 1.49 ;
 RECT 5.635 2.025 5.865 2.165 ;
 RECT 5.68 1.425 5.82 2.025 ;
 RECT 4.995 1.285 5.82 1.425 ;
 RECT 5.68 0.575 5.82 1.285 ;
 RECT 8.125 0.575 8.265 1.27 ;
 RECT 5.68 0.435 8.265 0.575 ;
 RECT 4.7 0.67 4.84 1.61 ;
 RECT 4.7 1.75 4.84 2.23 ;
 RECT 4.23 0.78 4.37 1.61 ;
 RECT 4.015 1.75 4.155 2.12 ;
 RECT 4.015 1.61 4.84 1.75 ;
 RECT 3.925 2.12 4.21 2.26 ;
 RECT 3.735 0.77 3.905 1.02 ;
 RECT 3.735 1.02 3.875 1.775 ;
 RECT 3.545 1.775 3.875 1.915 ;
 RECT 3.545 1.915 3.685 2.5 ;
 RECT 3.545 2.5 4.505 2.64 ;
 RECT 2.7 1.325 2.84 2.03 ;
 RECT 2.7 2.17 2.84 2.185 ;
 RECT 2.43 0.775 2.57 1.185 ;
 RECT 2.615 2.03 2.885 2.17 ;
 RECT 2.43 1.185 3.27 1.325 ;
 RECT 2.06 0.785 2.2 1.625 ;
 RECT 1.855 1.625 2.56 1.765 ;
 RECT 1.855 1.765 1.995 1.995 ;
 RECT 1.81 1.995 2.04 2.135 ;
 RECT 1.855 2.135 1.995 2.17 ;
 RECT 0.925 0.775 1.065 2.325 ;
 RECT 0.925 2.325 3.215 2.465 ;
 RECT 3.245 0.83 3.595 0.97 ;
 RECT 3.455 0.97 3.595 1.465 ;
 RECT 3.075 1.465 3.595 1.605 ;
 RECT 3.075 1.605 3.215 2.325 ;
 END
END LATCHX2

MACRO LNANDX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN RIN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 2.195 1.265 2.52 ;
 END
 ANTENNAGATEAREA 0.089 ;
 END RIN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.245 1.435 2.58 1.765 ;
 RECT 2.245 1.765 2.385 2.195 ;
 RECT 2.245 1.295 3.33 1.435 ;
 RECT 2.245 0.42 2.385 1.295 ;
 RECT 3.13 1.98 3.375 2.14 ;
 RECT 2.09 0.28 2.385 0.42 ;
 RECT 3.19 1.435 3.33 1.98 ;
 END
 ANTENNADIFFAREA 0.509 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.93 1.23 2.015 1.37 ;
 RECT 1.58 1.37 2.015 1.44 ;
 RECT 0.93 1.37 1.07 1.925 ;
 RECT 1.58 1.12 2.015 1.23 ;
 RECT 1.875 1.44 2.015 2.35 ;
 RECT 1.875 0.97 2.015 1.12 ;
 RECT 1.875 2.35 2.335 2.49 ;
 RECT 1.83 0.83 2.06 0.97 ;
 END
 ANTENNADIFFAREA 0.509 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 1.585 2.225 1.725 2.8 ;
 RECT 2.525 2.07 2.665 2.8 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 1.405 2.085 1.725 2.225 ;
 RECT 2.525 1.925 2.86 2.07 ;
 RECT 1.405 1.65 1.545 2.085 ;
 RECT 2.72 1.615 2.86 1.925 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 0.34 0.08 0.48 0.81 ;
 RECT 0.93 0.08 1.07 1.015 ;
 RECT 3.19 0.08 3.33 0.91 ;
 END
 END VSS

 PIN SIN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.975 2.28 3.32 2.555 ;
 END
 ANTENNAGATEAREA 0.089 ;
 END SIN

 OBS
 LAYER PO ;
 RECT 2.5 0.365 2.6 2.305 ;
 RECT 2.07 2.305 2.6 2.54 ;
 RECT 1.66 0.235 2.32 0.47 ;
 RECT 1.66 0.47 1.76 2.385 ;
 RECT 1.035 2.24 1.285 2.45 ;
 RECT 1.185 0.44 1.285 2.24 ;
 RECT 2.975 0.365 3.075 2.34 ;
 RECT 2.975 2.34 3.205 2.55 ;
 LAYER CO ;
 RECT 3.195 1.99 3.325 2.12 ;
 RECT 2.25 1.99 2.38 2.12 ;
 RECT 2.14 0.285 2.27 0.415 ;
 RECT 1.41 1.725 1.54 1.855 ;
 RECT 2.725 1.73 2.855 1.86 ;
 RECT 3.195 1.725 3.325 1.855 ;
 RECT 2.25 1.725 2.38 1.855 ;
 RECT 0.935 1.725 1.065 1.855 ;
 RECT 1.88 1.725 2.01 1.855 ;
 RECT 2.25 0.66 2.38 0.79 ;
 RECT 3.195 0.715 3.325 0.845 ;
 RECT 2.12 2.355 2.25 2.485 ;
 RECT 1.88 1.99 2.01 2.12 ;
 RECT 1.41 1.99 1.54 2.12 ;
 RECT 1.88 0.835 2.01 0.965 ;
 RECT 0.935 0.835 1.065 0.965 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 1.085 2.28 1.215 2.41 ;
 RECT 3.025 2.38 3.155 2.51 ;
 END
END LNANDX1

MACRO LNANDX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.4 BY 2.88 ;
 PIN RIN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.965 2.27 1.26 2.64 ;
 END
 ANTENNAGATEAREA 0.178 ;
 END RIN

 PIN SIN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.545 2.27 3.875 2.66 ;
 END
 ANTENNAGATEAREA 0.178 ;
 END SIN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.4 2.96 ;
 RECT 0.425 1.755 0.565 2.8 ;
 RECT 1.4 1.65 1.54 2.8 ;
 RECT 2.345 1.615 2.485 2.8 ;
 RECT 4.975 1.615 5.115 2.8 ;
 RECT 4.03 1.615 4.17 1.65 ;
 RECT 4.035 2.195 4.175 2.8 ;
 RECT 4.03 1.65 4.175 2.195 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.4 0.08 ;
 RECT 1.4 0.08 1.54 0.715 ;
 RECT 0.34 0.08 0.48 0.81 ;
 RECT 4.03 0.08 4.17 0.715 ;
 RECT 1.32 0.715 1.635 0.855 ;
 RECT 3.95 0.715 4.265 0.855 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.82 1.725 3.265 2.16 ;
 RECT 2.82 1.45 2.96 1.725 ;
 RECT 2.82 2.16 2.96 2.18 ;
 RECT 0.93 1.31 2.96 1.45 ;
 RECT 1.875 1.45 2.015 2.185 ;
 RECT 2.82 1.135 2.96 1.31 ;
 RECT 0.885 1.99 1.125 2.13 ;
 RECT 2.245 0.995 3.325 1.135 ;
 RECT 2.245 0.67 2.385 0.995 ;
 RECT 3.185 0.42 3.325 0.995 ;
 RECT 3.18 0.28 3.625 0.42 ;
 RECT 0.93 1.45 1.07 1.99 ;
 END
 ANTENNADIFFAREA 0.907 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.45 1.135 5.79 1.31 ;
 RECT 3.1 1.31 5.79 1.45 ;
 RECT 4.875 0.995 5.955 1.135 ;
 RECT 4.505 1.45 4.645 2.195 ;
 RECT 5.45 1.45 5.59 2.19 ;
 RECT 5.815 0.52 5.955 0.995 ;
 RECT 4.875 0.505 5.015 0.995 ;
 RECT 3.515 1.99 3.755 2.13 ;
 RECT 3.56 1.45 3.7 1.99 ;
 END
 ANTENNAGATEAREA 0.907 ;
 END Q

 OBS
 LAYER PO ;
 RECT 4.76 1.25 4.86 2.355 ;
 RECT 4.76 1.15 5.23 1.25 ;
 RECT 5.13 0.205 5.23 1.15 ;
 RECT 3.345 0.205 3.605 0.47 ;
 RECT 3.345 0.105 5.7 0.205 ;
 RECT 5.6 0.205 5.7 1.47 ;
 RECT 5.23 1.47 5.7 1.57 ;
 RECT 5.23 1.57 5.33 2.36 ;
 RECT 2.97 0.235 3.07 1.265 ;
 RECT 2.5 0.255 2.6 1.15 ;
 RECT 2.97 1.265 3.335 1.47 ;
 RECT 2.12 1.15 2.6 1.25 ;
 RECT 2.6 1.47 3.335 1.57 ;
 RECT 2.13 1.25 2.23 2.42 ;
 RECT 2.6 1.57 2.7 2.42 ;
 RECT 2.13 2.42 2.7 2.52 ;
 RECT 4.285 0.44 4.385 2.44 ;
 RECT 3.815 0.44 3.915 2.44 ;
 RECT 3.64 2.44 4.385 2.675 ;
 RECT 1.185 0.435 1.285 2.43 ;
 RECT 1.03 2.43 1.285 2.44 ;
 RECT 1.03 2.44 1.755 2.64 ;
 RECT 1.655 0.44 1.755 2.44 ;
 LAYER CO ;
 RECT 3.42 0.285 3.55 0.415 ;
 RECT 3.565 1.99 3.695 2.12 ;
 RECT 3.69 2.49 3.82 2.62 ;
 RECT 5.455 1.725 5.585 1.855 ;
 RECT 3.565 1.725 3.695 1.855 ;
 RECT 4.51 1.99 4.64 2.12 ;
 RECT 5.35 0.555 5.48 0.685 ;
 RECT 4.51 1.725 4.64 1.855 ;
 RECT 5.82 0.65 5.95 0.78 ;
 RECT 4.51 1.99 4.64 2.12 ;
 RECT 4.88 0.64 5.01 0.77 ;
 RECT 4.035 0.72 4.165 0.85 ;
 RECT 4.98 1.99 5.11 2.12 ;
 RECT 4.505 0.815 4.635 0.945 ;
 RECT 4.51 1.725 4.64 1.855 ;
 RECT 4.98 1.725 5.11 1.855 ;
 RECT 3.565 0.805 3.695 0.935 ;
 RECT 5.455 1.99 5.585 2.12 ;
 RECT 4.035 1.99 4.165 2.12 ;
 RECT 4.035 1.725 4.165 1.855 ;
 RECT 3.15 1.315 3.28 1.445 ;
 RECT 1.88 1.99 2.01 2.12 ;
 RECT 1.88 1.725 2.01 1.855 ;
 RECT 2.825 1.99 2.955 2.12 ;
 RECT 2.825 1.725 2.955 1.855 ;
 RECT 2.72 0.72 2.85 0.85 ;
 RECT 3.19 0.815 3.32 0.945 ;
 RECT 2.25 0.805 2.38 0.935 ;
 RECT 2.35 1.99 2.48 2.12 ;
 RECT 2.35 1.725 2.48 1.855 ;
 RECT 1.405 1.99 1.535 2.12 ;
 RECT 1.405 1.725 1.535 1.855 ;
 RECT 1.88 1.99 2.01 2.12 ;
 RECT 1.88 1.725 2.01 1.855 ;
 RECT 1.405 0.72 1.535 0.85 ;
 RECT 1.875 0.815 2.005 0.945 ;
 RECT 0.935 1.99 1.065 2.12 ;
 RECT 0.935 1.725 1.065 1.855 ;
 RECT 0.935 0.805 1.065 0.935 ;
 RECT 0.345 0.605 0.475 0.735 ;
 RECT 0.345 0.345 0.475 0.475 ;
 RECT 0.43 2.36 0.56 2.49 ;
 RECT 0.43 2.1 0.56 2.23 ;
 RECT 0.43 1.84 0.56 1.97 ;
 RECT 1.08 2.47 1.21 2.6 ;
 LAYER M1 ;
 RECT 3.56 0.67 3.7 0.995 ;
 RECT 4.5 0.36 4.64 0.995 ;
 RECT 3.56 0.995 4.64 1.135 ;
 RECT 5.34 0.69 5.48 0.855 ;
 RECT 5.265 0.55 5.58 0.69 ;
 RECT 5.34 0.36 5.48 0.55 ;
 RECT 4.5 0.22 5.48 0.36 ;
 RECT 0.93 0.67 1.07 0.995 ;
 RECT 1.87 0.475 2.01 0.995 ;
 RECT 0.93 0.995 2.01 1.135 ;
 RECT 2.635 0.715 2.95 0.855 ;
 RECT 2.71 0.475 2.85 0.715 ;
 RECT 1.87 0.335 2.85 0.475 ;
 END
END LNANDX2

MACRO MUX21X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 2.88 ;
 PIN S
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.95 1.475 1.475 1.75 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END S

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.735 1.13 1.875 1.48 ;
 RECT 1.64 1.63 2.585 1.79 ;
 RECT 1.64 1.48 1.885 1.63 ;
 RECT 2.435 1.79 2.575 1.845 ;
 RECT 2.435 1.57 2.575 1.63 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.1 1.155 2.52 1.415 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END IN1

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.4 0.36 3.65 0.6 ;
 RECT 3.51 0.6 3.65 2.25 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 RECT 1.13 2.005 1.27 2.8 ;
 RECT 0.24 1.545 0.38 2.8 ;
 RECT 3.04 2.03 3.18 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 3.04 0.08 3.18 0.78 ;
 RECT 0.24 0.08 0.38 0.88 ;
 RECT 1.13 0.08 1.27 0.97 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 2.105 1.41 2.205 1.645 ;
 RECT 2.335 0.555 2.435 1.18 ;
 RECT 2.055 1.745 2.155 2.735 ;
 RECT 2.055 1.645 2.205 1.745 ;
 RECT 2.105 1.18 2.435 1.41 ;
 RECT 2.825 0.405 2.925 2.735 ;
 RECT 2.62 0.175 2.925 0.405 ;
 RECT 1.72 0.555 1.82 1.145 ;
 RECT 1.68 1.145 1.925 1.385 ;
 RECT 2.525 1.82 2.625 2.735 ;
 RECT 2.385 1.59 2.625 1.82 ;
 RECT 3.295 0.335 3.395 1.155 ;
 RECT 3.295 1.365 3.395 2.745 ;
 RECT 3.105 1.155 3.395 1.365 ;
 RECT 0.915 1.475 1.485 1.75 ;
 RECT 1.385 0.555 1.485 1.475 ;
 RECT 1.385 1.75 1.485 2.735 ;
 RECT 0.915 0.555 1.015 1.475 ;
 RECT 0.915 1.75 1.015 2.685 ;
 LAYER CO ;
 RECT 3.045 2.35 3.175 2.48 ;
 RECT 3.045 0.585 3.175 0.715 ;
 RECT 2.08 0.775 2.21 0.905 ;
 RECT 2.275 2.115 2.405 2.245 ;
 RECT 1.135 0.775 1.265 0.905 ;
 RECT 0.665 0.775 0.795 0.905 ;
 RECT 1.135 2.055 1.265 2.185 ;
 RECT 0.665 2.055 0.795 2.185 ;
 RECT 3.045 2.09 3.175 2.22 ;
 RECT 1.135 2.315 1.265 2.445 ;
 RECT 3.515 1.79 3.645 1.92 ;
 RECT 3.155 1.195 3.285 1.325 ;
 RECT 3.515 2.05 3.645 2.18 ;
 RECT 3.515 0.775 3.645 0.905 ;
 RECT 2.67 0.225 2.8 0.355 ;
 RECT 2.26 1.23 2.39 1.36 ;
 RECT 1.14 1.55 1.27 1.68 ;
 RECT 0.245 0.69 0.375 0.82 ;
 RECT 0.245 0.43 0.375 0.56 ;
 RECT 0.245 2.12 0.375 2.25 ;
 RECT 0.245 1.86 0.375 1.99 ;
 RECT 0.245 1.6 0.375 1.73 ;
 RECT 2.44 1.64 2.57 1.77 ;
 RECT 1.74 1.195 1.87 1.325 ;
 LAYER M1 ;
 RECT 2.73 0.91 2.87 1.19 ;
 RECT 2.73 1.33 2.87 2.11 ;
 RECT 2.025 0.77 2.87 0.91 ;
 RECT 2.22 2.11 2.87 2.25 ;
 RECT 2.73 1.19 3.29 1.33 ;
 RECT 3.15 1.145 3.29 1.19 ;
 RECT 3.15 1.33 3.29 1.375 ;
 RECT 0.66 0.72 0.8 1.195 ;
 RECT 0.66 1.335 0.8 2.27 ;
 RECT 1.445 0.36 1.585 1.195 ;
 RECT 0.66 1.195 1.585 1.335 ;
 RECT 1.445 0.22 2.87 0.36 ;
 END
END MUX21X1

MACRO AND4X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 0.84 1.055 1.08 ;
 END
 ANTENNAGATEAREA 0.052 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 1.8 1.575 2.125 ;
 END
 ANTENNAGATEAREA 0.052 ;
 END IN2

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.8 0.715 2.215 1.075 ;
 END
 ANTENNAGATEAREA 0.052 ;
 END IN3

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.11 2.36 2.53 2.66 ;
 END
 ANTENNAGATEAREA 0.052 ;
 END IN4

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.08 0.45 3.405 0.825 ;
 RECT 3.22 0.825 3.36 2.26 ;
 RECT 3.22 0.34 3.36 0.45 ;
 END
 ANTENNADIFFAREA 0.449 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.525 2.96 ;
 RECT 2.605 1.56 2.875 1.7 ;
 RECT 1.72 1.51 1.86 2.8 ;
 RECT 0.37 1.495 0.51 2.8 ;
 RECT 0.78 1.51 0.92 2.8 ;
 RECT 2.67 1.7 2.81 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 2.67 0.08 2.81 0.6 ;
 RECT 0.365 0.08 0.505 0.91 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 2.45 0.1 2.55 2.37 ;
 RECT 2.32 2.37 2.55 2.6 ;
 RECT 1.975 0.105 2.075 0.76 ;
 RECT 1.975 0.99 2.075 1.915 ;
 RECT 1.975 0.76 2.205 0.99 ;
 RECT 3 0.105 3.1 1.155 ;
 RECT 3 1.385 3.1 2.76 ;
 RECT 2.73 1.155 3.1 1.385 ;
 RECT 1.035 1.075 1.135 1.92 ;
 RECT 1.035 0.105 1.135 0.845 ;
 RECT 0.825 0.845 1.135 1.075 ;
 RECT 1.505 0.105 1.605 1.89 ;
 RECT 1.375 1.89 1.605 2.12 ;
 LAYER CO ;
 RECT 0.375 2.065 0.505 2.195 ;
 RECT 0.375 1.805 0.505 1.935 ;
 RECT 0.375 1.545 0.505 1.675 ;
 RECT 0.37 0.47 0.5 0.6 ;
 RECT 0.37 0.73 0.5 0.86 ;
 RECT 1.425 1.94 1.555 2.07 ;
 RECT 2.365 2.42 2.495 2.55 ;
 RECT 2.015 0.81 2.145 0.94 ;
 RECT 2.675 0.41 2.805 0.54 ;
 RECT 2.675 1.565 2.805 1.695 ;
 RECT 2.195 1.5 2.325 1.63 ;
 RECT 0.785 0.41 0.915 0.54 ;
 RECT 3.225 0.52 3.355 0.65 ;
 RECT 0.785 1.56 0.915 1.69 ;
 RECT 3.225 1.82 3.355 1.95 ;
 RECT 3.225 2.08 3.355 2.21 ;
 RECT 2.78 1.205 2.91 1.335 ;
 RECT 1.255 1.505 1.385 1.635 ;
 RECT 3.225 1.56 3.355 1.69 ;
 RECT 1.725 1.56 1.855 1.69 ;
 RECT 0.875 0.895 1.005 1.025 ;
 RECT 1.725 1.56 1.855 1.69 ;
 LAYER M1 ;
 RECT 0.78 0.325 0.92 0.51 ;
 RECT 0.78 0.43 0.92 0.615 ;
 RECT 0.905 0.475 1.39 0.615 ;
 RECT 1.185 1.5 1.455 1.64 ;
 RECT 1.25 0.55 1.39 1.345 ;
 RECT 1.25 1.245 1.39 1.64 ;
 RECT 2.19 1.24 2.33 1.7 ;
 RECT 2.73 1.155 2.995 1.385 ;
 RECT 2.73 1.195 2.96 1.345 ;
 RECT 1.25 1.215 2.96 1.355 ;
 END
END AND4X1

MACRO AND4X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.215 1.885 1.58 2.215 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN2

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.985 0.52 2.36 0.845 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 2.67 0.08 2.81 0.505 ;
 RECT 0.365 0.08 0.505 0.91 ;
 RECT 3.725 0.08 3.865 0.505 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 0.37 1.495 0.51 2.8 ;
 RECT 2.67 1.515 2.81 2.8 ;
 RECT 1.72 1.51 1.86 2.8 ;
 RECT 3.73 1.515 3.87 2.8 ;
 RECT 0.78 1.51 0.92 2.8 ;
 END
 END VDD

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.085 2.05 2.53 2.43 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN4

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.8 0.815 1.08 1.095 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN1

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.22 1.16 3.64 1.4 ;
 RECT 3.22 1.4 3.36 2.62 ;
 RECT 3.22 0.27 3.36 1.16 ;
 END
 ANTENNADIFFAREA 0.584 ;
 END Q

 OBS
 LAYER PO ;
 RECT 1.035 0.105 1.135 0.845 ;
 RECT 1.035 1.075 1.135 1.92 ;
 RECT 0.825 0.845 1.135 1.075 ;
 RECT 2.845 1.2 3.59 1.3 ;
 RECT 3.49 0.105 3.59 1.2 ;
 RECT 3 0.105 3.1 1.15 ;
 RECT 2.845 1.15 3.1 1.2 ;
 RECT 2.845 1.3 3.1 1.38 ;
 RECT 3.49 1.3 3.59 2.76 ;
 RECT 3 1.38 3.1 2.76 ;
 RECT 2.45 0.1 2.55 2.055 ;
 RECT 2.32 2.055 2.55 2.285 ;
 RECT 1.505 0.105 1.605 1.885 ;
 RECT 1.375 1.885 1.605 2.115 ;
 RECT 1.975 0.105 2.075 0.615 ;
 RECT 1.975 0.845 2.075 1.915 ;
 RECT 1.975 0.615 2.21 0.845 ;
 LAYER CO ;
 RECT 3.225 2.345 3.355 2.475 ;
 RECT 3.735 1.565 3.865 1.695 ;
 RECT 3.735 1.565 3.865 1.695 ;
 RECT 3.735 2.375 3.865 2.505 ;
 RECT 3.735 2.1 3.865 2.23 ;
 RECT 3.735 1.835 3.865 1.965 ;
 RECT 2.675 2.35 2.805 2.48 ;
 RECT 2.675 2.09 2.805 2.22 ;
 RECT 2.675 1.83 2.805 1.96 ;
 RECT 3.73 0.325 3.86 0.455 ;
 RECT 3.735 1.565 3.865 1.695 ;
 RECT 2.37 2.105 2.5 2.235 ;
 RECT 0.375 1.545 0.505 1.675 ;
 RECT 1.255 1.56 1.385 1.69 ;
 RECT 0.375 1.805 0.505 1.935 ;
 RECT 3.225 0.325 3.355 0.455 ;
 RECT 0.37 0.47 0.5 0.6 ;
 RECT 1.425 1.935 1.555 2.065 ;
 RECT 2.195 1.5 2.325 1.63 ;
 RECT 2.895 1.2 3.025 1.33 ;
 RECT 3.225 2.08 3.355 2.21 ;
 RECT 0.375 2.065 0.505 2.195 ;
 RECT 1.725 1.56 1.855 1.69 ;
 RECT 2.675 1.565 2.805 1.695 ;
 RECT 0.875 0.895 1.005 1.025 ;
 RECT 2.015 0.665 2.145 0.795 ;
 RECT 1.725 1.56 1.855 1.69 ;
 RECT 0.785 1.56 0.915 1.69 ;
 RECT 3.225 1.56 3.355 1.69 ;
 RECT 0.785 0.325 0.915 0.455 ;
 RECT 0.37 0.73 0.5 0.86 ;
 RECT 3.225 1.82 3.355 1.95 ;
 RECT 2.675 0.325 2.805 0.455 ;
 LAYER M1 ;
 RECT 1.66 0.55 1.8 1.345 ;
 RECT 0.905 0.475 1.8 0.615 ;
 RECT 1.25 1.245 1.39 1.74 ;
 RECT 0.78 0.43 0.92 0.615 ;
 RECT 0.78 0.275 0.92 0.46 ;
 RECT 2.19 1.24 2.33 1.69 ;
 RECT 1.25 1.21 2.33 1.35 ;
 RECT 2.845 1.19 3.075 1.34 ;
 RECT 2.195 1.21 3.075 1.35 ;
 END
END AND4X2

MACRO MUX41X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.64 BY 2.88 ;
 PIN S0
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.64 1.155 2.07 1.295 ;
 RECT 1.64 1.295 1.97 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END S0

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.355 1.315 4.605 1.72 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END IN4

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.64 2.96 ;
 RECT 7.915 1.71 8.055 2.8 ;
 RECT 4.21 2.33 4.35 2.8 ;
 RECT 0.31 1.545 0.45 2.8 ;
 RECT 1.705 1.795 1.845 2.8 ;
 RECT 6.15 1.71 6.29 2.8 ;
 RECT 0.765 1.795 0.905 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.64 0.08 ;
 RECT 0.765 0.08 0.905 0.775 ;
 RECT 4.22 0.08 4.36 0.785 ;
 RECT 6.15 0.08 6.29 0.805 ;
 RECT 1.705 0.08 1.845 0.775 ;
 RECT 7.915 0.08 8.055 0.805 ;
 RECT 0.315 0.08 0.455 0.88 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.395 2.265 7.775 2.52 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.43 2.27 6.715 2.52 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 1.14 1.375 1.4 ;
 RECT 1.235 1.4 1.375 1.96 ;
 RECT 1.235 0.735 1.375 1.14 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END Q

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.64 2.28 6.01 2.52 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END IN3

 PIN S1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.195 2.1 8.445 2.43 ;
 END
 ANTENNAGATEAREA 0.233 ;
 END S1

 OBS
 LAYER PO ;
 RECT 7.59 1.53 7.69 2.295 ;
 RECT 7.7 0.4 7.8 1.43 ;
 RECT 7.59 1.43 7.8 1.53 ;
 RECT 7.59 2.295 7.82 2.505 ;
 RECT 5.255 0.87 5.745 0.97 ;
 RECT 5.255 0.4 5.355 0.87 ;
 RECT 5.535 0.97 5.745 1.13 ;
 RECT 6.405 0.4 6.505 2.295 ;
 RECT 6.405 2.295 6.635 2.505 ;
 RECT 1.49 0.35 1.59 1.09 ;
 RECT 1.49 1.19 1.59 2.645 ;
 RECT 1.02 0.35 1.12 1.09 ;
 RECT 1.02 1.19 1.12 2.745 ;
 RECT 2.495 2.34 2.595 2.645 ;
 RECT 1.02 1.09 1.59 1.19 ;
 RECT 1.49 2.645 2.595 2.745 ;
 RECT 2.43 2.13 2.66 2.34 ;
 RECT 4.475 0.385 4.575 1.325 ;
 RECT 4.475 1.535 4.575 2.395 ;
 RECT 4.345 1.325 4.575 1.535 ;
 RECT 7.285 0.4 7.385 1.035 ;
 RECT 4.775 1.435 4.875 2.685 ;
 RECT 6.815 1.25 6.915 2.685 ;
 RECT 6.815 1.15 7.515 1.245 ;
 RECT 7.285 1.035 7.515 1.15 ;
 RECT 6.815 1.245 7.385 1.25 ;
 RECT 4.775 2.685 6.915 2.785 ;
 RECT 1.96 0.57 2.06 1.11 ;
 RECT 1.96 1.34 2.06 1.835 ;
 RECT 1.85 1.15 3.6 1.25 ;
 RECT 1.85 1.11 2.06 1.15 ;
 RECT 1.85 1.25 2.06 1.34 ;
 RECT 3.5 0.4 3.6 1.15 ;
 RECT 3.03 1.25 3.13 2.545 ;
 RECT 3.03 0.43 3.13 0.97 ;
 RECT 3.03 0.22 3.24 0.43 ;
 RECT 3.5 1.485 3.6 2.445 ;
 RECT 3.5 2.445 4.105 2.545 ;
 RECT 4.005 0.22 4.105 2.445 ;
 RECT 3.03 0.12 4.105 0.22 ;
 RECT 8.17 2.21 8.415 2.42 ;
 RECT 5.245 1.25 5.345 2.395 ;
 RECT 4.785 0.22 4.885 1.15 ;
 RECT 6.815 0.22 6.915 0.97 ;
 RECT 7.285 1.435 7.385 2.685 ;
 RECT 4.785 0.12 8.27 0.22 ;
 RECT 8.17 0.22 8.27 2.21 ;
 RECT 8.17 2.42 8.27 2.685 ;
 RECT 4.785 1.15 5.345 1.25 ;
 RECT 7.285 2.685 8.27 2.785 ;
 RECT 5.935 0.4 6.035 2.295 ;
 RECT 5.81 2.295 6.04 2.505 ;
 LAYER CO ;
 RECT 1.24 1.515 1.37 1.645 ;
 RECT 7.92 0.62 8.05 0.75 ;
 RECT 1.71 0.59 1.84 0.72 ;
 RECT 7.035 1.715 7.165 1.845 ;
 RECT 1.89 1.16 2.02 1.29 ;
 RECT 0.77 2.11 0.9 2.24 ;
 RECT 0.77 1.85 0.9 1.98 ;
 RECT 0.77 2.37 0.9 2.5 ;
 RECT 0.77 0.59 0.9 0.72 ;
 RECT 1.24 1.775 1.37 1.905 ;
 RECT 2.48 2.17 2.61 2.3 ;
 RECT 6.455 2.335 6.585 2.465 ;
 RECT 4.995 1.665 5.125 1.795 ;
 RECT 7.335 1.075 7.465 1.205 ;
 RECT 6.155 0.62 6.285 0.75 ;
 RECT 7.035 0.62 7.165 0.75 ;
 RECT 5.005 0.62 5.135 0.75 ;
 RECT 0.315 1.86 0.445 1.99 ;
 RECT 7.64 2.335 7.77 2.465 ;
 RECT 4.215 2.39 4.345 2.52 ;
 RECT 0.32 0.69 0.45 0.82 ;
 RECT 6.155 2.03 6.285 2.16 ;
 RECT 7.92 2.03 8.05 2.16 ;
 RECT 3.72 1.715 3.85 1.845 ;
 RECT 0.315 1.6 0.445 1.73 ;
 RECT 4.395 1.365 4.525 1.495 ;
 RECT 2.78 0.62 2.91 0.75 ;
 RECT 7.92 1.77 8.05 1.9 ;
 RECT 4.225 0.605 4.355 0.735 ;
 RECT 0.32 0.43 0.45 0.56 ;
 RECT 7.035 1.975 7.165 2.105 ;
 RECT 2.78 1.705 2.91 1.835 ;
 RECT 1.24 0.79 1.37 0.92 ;
 RECT 2.18 1.485 2.31 1.615 ;
 RECT 5.575 0.95 5.705 1.08 ;
 RECT 8.39 1.695 8.52 1.825 ;
 RECT 8.39 0.62 8.52 0.75 ;
 RECT 3.72 0.62 3.85 0.75 ;
 RECT 3.25 0.62 3.38 0.75 ;
 RECT 1.71 2.37 1.84 2.5 ;
 RECT 0.315 2.12 0.445 2.25 ;
 RECT 5.86 2.335 5.99 2.465 ;
 RECT 3.07 0.25 3.2 0.38 ;
 RECT 1.71 1.85 1.84 1.98 ;
 RECT 2.225 0.79 2.355 0.92 ;
 RECT 3.25 1.715 3.38 1.845 ;
 RECT 1.71 2.11 1.84 2.24 ;
 RECT 8.235 2.25 8.365 2.38 ;
 RECT 6.155 1.77 6.285 1.9 ;
 LAYER M1 ;
 RECT 6.43 0.41 6.57 0.945 ;
 RECT 7.33 1.205 7.47 1.255 ;
 RECT 5.525 0.945 6.57 1.085 ;
 RECT 6.43 0.27 7.47 0.41 ;
 RECT 7.33 0.41 7.47 1.065 ;
 RECT 8.385 0.565 8.525 1.065 ;
 RECT 8.385 1.205 8.525 1.895 ;
 RECT 7.33 1.065 8.525 1.205 ;
 RECT 3.245 0.56 3.385 2.05 ;
 RECT 2.475 2.19 2.615 2.35 ;
 RECT 2.475 2.05 3.385 2.19 ;
 RECT 2.22 0.385 2.36 1.48 ;
 RECT 2.22 0.245 3.25 0.385 ;
 RECT 2.12 1.48 2.36 1.62 ;
 RECT 3.57 2.045 5.485 2.115 ;
 RECT 3.565 2.115 5.485 2.18 ;
 RECT 5.345 1.365 5.485 2.04 ;
 RECT 3.995 2.04 5.485 2.045 ;
 RECT 3.565 2.185 3.705 2.5 ;
 RECT 3.565 2.18 4.135 2.185 ;
 RECT 2.125 2.5 3.705 2.64 ;
 RECT 2.775 0.56 2.915 1.76 ;
 RECT 2.125 1.9 2.265 2.5 ;
 RECT 2.125 1.76 2.915 1.9 ;
 RECT 7.03 0.56 7.17 1.225 ;
 RECT 7.03 1.365 7.17 2.17 ;
 RECT 5.345 1.225 7.17 1.365 ;
 RECT 3.715 0.56 3.855 0.925 ;
 RECT 3.715 1.065 3.855 1.905 ;
 RECT 3.715 0.925 5.14 1.065 ;
 RECT 5 0.57 5.14 0.925 ;
 RECT 4.99 1.065 5.13 1.87 ;
 END
END MUX41X2

MACRO OA21X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.645 2.12 0.92 2.42 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END IN2

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 1.16 1.36 1.4 ;
 END
 ANTENNAGATEAREA 0.051 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 2.78 0.08 2.92 0.835 ;
 RECT 1.895 0.08 2.035 0.78 ;
 RECT 0.585 0.08 0.725 0.72 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.165 1.16 0.44 1.435 ;
 END
 ANTENNAGATEAREA 0.069 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 2.78 1.645 2.92 2.8 ;
 RECT 1.525 1.83 1.665 2.8 ;
 RECT 1.895 1.555 2.035 2.8 ;
 RECT 0.115 1.775 0.255 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.365 1.4 2.505 2.585 ;
 RECT 2.365 1.16 2.715 1.4 ;
 RECT 2.365 0.695 2.505 1.16 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END Q

 OBS
 LAYER PO ;
 RECT 1.31 0.33 1.41 1.175 ;
 RECT 1.31 1.385 1.41 2.23 ;
 RECT 1.175 1.175 1.41 1.385 ;
 RECT 0.84 0.4 0.94 2.155 ;
 RECT 0.71 2.155 0.94 2.365 ;
 RECT 2.15 0.35 2.25 1.115 ;
 RECT 2.15 1.325 2.25 2.74 ;
 RECT 2.02 1.115 2.25 1.325 ;
 RECT 0.37 1.395 0.47 2.23 ;
 RECT 0.37 0.4 0.47 1.185 ;
 RECT 0.23 1.185 0.47 1.395 ;
 LAYER CO ;
 RECT 1.9 2.39 2.03 2.52 ;
 RECT 1.9 1.87 2.03 2 ;
 RECT 1.9 2.13 2.03 2.26 ;
 RECT 1.9 1.61 2.03 1.74 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 1.06 0.55 1.19 0.68 ;
 RECT 2.37 1.87 2.5 2 ;
 RECT 2.07 1.155 2.2 1.285 ;
 RECT 1.9 0.595 2.03 0.725 ;
 RECT 0.59 0.54 0.72 0.67 ;
 RECT 2.785 0.395 2.915 0.525 ;
 RECT 2.785 1.695 2.915 1.825 ;
 RECT 1.53 1.88 1.66 2.01 ;
 RECT 0.12 0.54 0.25 0.67 ;
 RECT 2.37 2.13 2.5 2.26 ;
 RECT 0.28 1.225 0.41 1.355 ;
 RECT 0.76 2.195 0.89 2.325 ;
 RECT 2.37 2.39 2.5 2.52 ;
 RECT 2.785 2.215 2.915 2.345 ;
 RECT 2.37 0.76 2.5 0.89 ;
 RECT 2.785 0.655 2.915 0.785 ;
 RECT 2.785 1.955 2.915 2.085 ;
 RECT 2.37 1.61 2.5 1.74 ;
 RECT 1.225 1.215 1.355 1.345 ;
 RECT 0.12 1.83 0.25 1.96 ;
 RECT 1.06 1.87 1.19 2 ;
 LAYER M1 ;
 RECT 1.525 0.49 1.665 1.15 ;
 RECT 1.525 1.29 1.665 1.54 ;
 RECT 1.055 1.54 1.665 1.68 ;
 RECT 1.055 1.68 1.195 2.05 ;
 RECT 2.065 1.105 2.205 1.15 ;
 RECT 2.065 1.29 2.205 1.335 ;
 RECT 1.525 1.15 2.205 1.29 ;
 RECT 0.115 0.49 0.255 0.86 ;
 RECT 1.055 0.5 1.195 0.86 ;
 RECT 0.115 0.86 1.195 1 ;
 END
END OA21X1

MACRO OA21X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.365 1.4 2.505 2.585 ;
 RECT 2.365 1.16 2.865 1.4 ;
 RECT 2.365 0.585 2.505 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END Q

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.665 1.16 0.92 1.435 ;
 END
 ANTENNAGATEAREA 0.089 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 3.25 0.08 3.39 0.835 ;
 RECT 1.895 0.08 2.035 0.785 ;
 RECT 0.585 0.08 0.725 0.73 ;
 RECT 2.835 0.08 2.975 0.785 ;
 END
 END VSS

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.365 1.48 1.72 1.72 ;
 END
 ANTENNAGATEAREA 0.051 ;
 END IN3

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 RECT 1.525 1.895 1.665 2.8 ;
 RECT 1.895 2.095 2.035 2.8 ;
 RECT 0.115 1.785 0.255 2.8 ;
 RECT 3.25 1.645 3.39 2.8 ;
 RECT 2.835 2.095 2.975 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.165 1.155 0.44 1.425 ;
 END
 ANTENNAGATEAREA 0.089 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 0.37 1.4 0.47 2.48 ;
 RECT 0.37 0.33 0.47 1.19 ;
 RECT 0.205 1.19 0.47 1.4 ;
 RECT 0.84 0.33 0.94 1.215 ;
 RECT 0.84 1.425 0.94 2.485 ;
 RECT 0.7 1.215 0.94 1.425 ;
 RECT 1.31 1.495 1.55 1.705 ;
 RECT 1.31 1.705 1.41 2.35 ;
 RECT 1.31 0.33 1.41 1.495 ;
 RECT 2.62 1.305 2.72 2.755 ;
 RECT 2.62 0.33 2.72 1.205 ;
 RECT 2.02 1.205 2.72 1.305 ;
 RECT 2.02 1.115 2.25 1.205 ;
 RECT 2.02 1.305 2.25 1.325 ;
 RECT 2.15 0.33 2.25 1.115 ;
 RECT 2.15 1.325 2.25 2.755 ;
 LAYER CO ;
 RECT 1.06 1.69 1.19 1.82 ;
 RECT 0.12 1.845 0.25 1.975 ;
 RECT 2.84 0.6 2.97 0.73 ;
 RECT 2.84 2.145 2.97 2.275 ;
 RECT 2.84 2.405 2.97 2.535 ;
 RECT 3.255 0.655 3.385 0.785 ;
 RECT 1.06 1.95 1.19 2.08 ;
 RECT 0.12 2.105 0.25 2.235 ;
 RECT 1.37 1.535 1.5 1.665 ;
 RECT 2.37 1.625 2.5 1.755 ;
 RECT 3.255 2.215 3.385 2.345 ;
 RECT 2.37 0.64 2.5 0.77 ;
 RECT 1.9 0.6 2.03 0.73 ;
 RECT 1.06 0.55 1.19 0.68 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 3.255 0.395 3.385 0.525 ;
 RECT 2.37 1.885 2.5 2.015 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 2.07 1.155 2.2 1.285 ;
 RECT 3.255 1.695 3.385 1.825 ;
 RECT 1.9 2.405 2.03 2.535 ;
 RECT 1.53 1.95 1.66 2.08 ;
 RECT 0.75 1.255 0.88 1.385 ;
 RECT 0.255 1.23 0.385 1.36 ;
 RECT 2.37 2.145 2.5 2.275 ;
 RECT 2.37 2.405 2.5 2.535 ;
 RECT 0.12 0.55 0.25 0.68 ;
 RECT 3.255 1.955 3.385 2.085 ;
 RECT 1.9 2.145 2.03 2.275 ;
 LAYER M1 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.5 1.195 0.87 ;
 RECT 0.115 0.87 1.195 1.01 ;
 RECT 1.525 0.495 1.665 1.15 ;
 RECT 1.06 1.29 1.2 1.575 ;
 RECT 1.055 1.575 1.2 1.63 ;
 RECT 1.055 1.63 1.195 2.135 ;
 RECT 1.06 1.15 2.205 1.29 ;
 RECT 2.065 1.105 2.205 1.15 ;
 RECT 2.065 1.29 2.205 1.335 ;
 END
END OA21X2

MACRO OA221X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 2.215 0.925 2.52 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN2

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.045 1.16 1.4 1.4 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN4

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 4.09 1.645 4.23 2.8 ;
 RECT 0.115 1.88 0.255 2.8 ;
 RECT 1.995 1.88 2.135 2.8 ;
 RECT 3.205 2.095 3.345 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.675 1.4 3.815 2.585 ;
 RECT 3.675 1.16 3.98 1.4 ;
 RECT 3.675 0.725 3.815 1.16 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END Q

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.28 0.98 2.52 1.33 ;
 END
 ANTENNAGATEAREA 0.055 ;
 END IN5

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.165 1.155 0.44 1.465 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.61 1.155 1.905 1.405 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 4.09 0.08 4.23 0.835 ;
 RECT 3.205 0.08 3.345 0.765 ;
 RECT 0.585 0.08 0.725 0.73 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.37 0.33 0.47 1.165 ;
 RECT 0.205 1.165 0.47 1.375 ;
 RECT 0.37 1.375 0.47 2.335 ;
 RECT 2.62 0.41 2.72 1.01 ;
 RECT 2.25 1.11 2.49 1.225 ;
 RECT 2.25 1.225 2.35 2.035 ;
 RECT 2.25 1.01 2.72 1.11 ;
 RECT 1.78 0.33 1.88 1.17 ;
 RECT 1.78 1.38 1.88 2.335 ;
 RECT 1.635 1.17 1.88 1.38 ;
 RECT 1.31 0.33 1.41 1.175 ;
 RECT 1.31 1.385 1.41 2.335 ;
 RECT 1.18 1.175 1.41 1.385 ;
 RECT 3.46 1.325 3.56 2.755 ;
 RECT 3.46 0.35 3.56 1.115 ;
 RECT 3.33 1.115 3.56 1.325 ;
 RECT 0.84 0.33 0.94 2.245 ;
 RECT 0.71 2.245 0.94 2.455 ;
 LAYER CO ;
 RECT 3.68 0.775 3.81 0.905 ;
 RECT 0.12 1.935 0.25 2.065 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 3.21 2.145 3.34 2.275 ;
 RECT 2.47 1.685 2.6 1.815 ;
 RECT 3.68 2.405 3.81 2.535 ;
 RECT 2.37 0.64 2.5 0.77 ;
 RECT 1.06 0.55 1.19 0.68 ;
 RECT 1.23 1.215 1.36 1.345 ;
 RECT 3.38 1.155 3.51 1.285 ;
 RECT 3.68 1.885 3.81 2.015 ;
 RECT 4.095 1.955 4.225 2.085 ;
 RECT 4.095 1.695 4.225 1.825 ;
 RECT 3.68 2.145 3.81 2.275 ;
 RECT 0.76 2.285 0.89 2.415 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 2.84 0.64 2.97 0.77 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 2 1.935 2.13 2.065 ;
 RECT 1.06 1.71 1.19 1.84 ;
 RECT 3.68 1.625 3.81 1.755 ;
 RECT 4.095 0.655 4.225 0.785 ;
 RECT 3.21 0.58 3.34 0.71 ;
 RECT 0.12 0.55 0.25 0.68 ;
 RECT 4.095 0.395 4.225 0.525 ;
 RECT 2.31 1.055 2.44 1.185 ;
 RECT 1.685 1.21 1.815 1.34 ;
 RECT 4.095 2.215 4.225 2.345 ;
 RECT 0.255 1.205 0.385 1.335 ;
 RECT 3.21 2.405 3.34 2.535 ;
 LAYER M1 ;
 RECT 2.365 0.36 2.505 0.825 ;
 RECT 1.525 0.22 2.505 0.36 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 1.055 1.69 1.195 1.9 ;
 RECT 2.465 1.69 2.605 1.885 ;
 RECT 2.835 0.59 2.975 1.19 ;
 RECT 2.835 1.33 2.975 1.55 ;
 RECT 1.055 1.55 2.975 1.69 ;
 RECT 3.375 1.105 3.515 1.19 ;
 RECT 3.375 1.33 3.515 1.335 ;
 RECT 2.835 1.19 3.515 1.33 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.495 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 END
END OA221X1

MACRO OA221X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.34 1.605 1.72 1.89 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN4

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 4.56 0.08 4.7 0.835 ;
 RECT 3.205 0.08 3.345 0.855 ;
 RECT 0.585 0.08 0.725 0.73 ;
 RECT 4.145 0.08 4.285 0.855 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.13 1.48 0.445 1.755 ;
 END
 ANTENNAGATEAREA 0.078 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 4.56 1.645 4.7 2.8 ;
 RECT 1.995 2.085 2.135 2.8 ;
 RECT 3.205 2.095 3.345 2.8 ;
 RECT 0.115 2.225 0.255 2.8 ;
 RECT 4.145 2.095 4.285 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.675 1.4 3.815 2.585 ;
 RECT 3.675 1.16 4.155 1.4 ;
 RECT 3.675 0.62 3.815 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END Q

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.595 1.3 0.92 1.59 ;
 END
 ANTENNAGATEAREA 0.078 ;
 END IN2

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.86 1.645 2.22 1.89 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN3

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.375 2.275 2.68 2.525 ;
 END
 ANTENNAGATEAREA 0.055 ;
 END IN5

 OBS
 LAYER PO ;
 RECT 0.84 0.33 0.94 1.37 ;
 RECT 0.84 1.58 0.94 2.745 ;
 RECT 0.7 1.37 0.94 1.58 ;
 RECT 1.78 0.33 1.88 1.655 ;
 RECT 1.78 1.655 2.15 1.865 ;
 RECT 1.78 1.865 1.88 2.745 ;
 RECT 1.31 0.33 1.41 1.655 ;
 RECT 1.31 1.865 1.41 2.745 ;
 RECT 1.31 1.655 1.55 1.865 ;
 RECT 3.93 0.32 4.03 1.145 ;
 RECT 3.33 1.145 4.03 1.245 ;
 RECT 3.93 1.245 4.03 2.755 ;
 RECT 3.33 1.115 3.56 1.145 ;
 RECT 3.33 1.245 3.56 1.325 ;
 RECT 3.46 1.325 3.56 2.755 ;
 RECT 3.46 0.32 3.56 1.115 ;
 RECT 2.62 0.33 2.72 1.01 ;
 RECT 2.34 1.01 2.72 1.11 ;
 RECT 2.34 1.11 2.44 2.275 ;
 RECT 2.34 2.275 2.635 2.485 ;
 RECT 0.37 1.745 0.47 2.745 ;
 RECT 0.37 0.33 0.47 1.535 ;
 RECT 0.205 1.535 0.47 1.745 ;
 LAYER CO ;
 RECT 4.15 2.405 4.28 2.535 ;
 RECT 4.15 2.145 4.28 2.275 ;
 RECT 4.15 0.675 4.28 0.805 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 3.21 2.405 3.34 2.535 ;
 RECT 0.12 2.305 0.25 2.435 ;
 RECT 0.255 1.575 0.385 1.705 ;
 RECT 1.06 0.55 1.19 0.68 ;
 RECT 4.565 0.655 4.695 0.785 ;
 RECT 3.68 0.675 3.81 0.805 ;
 RECT 3.68 2.145 3.81 2.275 ;
 RECT 2.56 1.995 2.69 2.125 ;
 RECT 3.68 2.405 3.81 2.535 ;
 RECT 1.97 1.695 2.1 1.825 ;
 RECT 4.565 2.215 4.695 2.345 ;
 RECT 2.37 0.56 2.5 0.69 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 4.565 0.395 4.695 0.525 ;
 RECT 3.38 1.155 3.51 1.285 ;
 RECT 4.565 1.955 4.695 2.085 ;
 RECT 4.565 1.695 4.695 1.825 ;
 RECT 1.06 2.285 1.19 2.415 ;
 RECT 1.37 1.695 1.5 1.825 ;
 RECT 3.68 1.885 3.81 2.015 ;
 RECT 0.12 0.55 0.25 0.68 ;
 RECT 2 2.165 2.13 2.295 ;
 RECT 2.84 0.56 2.97 0.69 ;
 RECT 0.75 1.41 0.88 1.54 ;
 RECT 3.21 0.675 3.34 0.805 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 3.21 2.145 3.34 2.275 ;
 RECT 3.68 1.625 3.81 1.755 ;
 RECT 2.455 2.315 2.585 2.445 ;
 LAYER M1 ;
 RECT 2.365 0.36 2.505 0.745 ;
 RECT 1.525 0.22 2.505 0.36 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 2.835 0.51 2.975 1.15 ;
 RECT 2.835 1.29 2.975 1.99 ;
 RECT 2.5 1.99 2.975 2.13 ;
 RECT 1.055 1.63 1.2 1.7 ;
 RECT 1.055 1.7 1.195 2.535 ;
 RECT 1.06 1.29 1.2 1.63 ;
 RECT 1.06 1.15 3.53 1.29 ;
 RECT 3.375 1.105 3.515 1.15 ;
 RECT 3.375 1.29 3.515 1.335 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.495 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 END
END OA221X2

MACRO OA222X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.405 2.1 0.775 2.47 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 4.64 1.645 4.78 2.8 ;
 RECT 0.115 1.745 0.255 2.8 ;
 RECT 1.995 1.78 2.135 2.8 ;
 RECT 3.675 2.095 3.815 2.8 ;
 END
 END VDD

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.275 2.07 2.545 2.42 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END IN5

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 1.945 1.855 2.305 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END IN3

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.495 1.16 0.885 1.41 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 0.585 0.08 0.725 0.73 ;
 RECT 3.675 0.08 3.815 0.76 ;
 RECT 4.56 0.08 4.7 0.835 ;
 END
 END VSS

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.965 2.285 1.26 2.655 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END IN4

 PIN IN6
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.825 2.09 3.145 2.365 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END IN6

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.145 1.415 4.285 2.585 ;
 RECT 4.145 1.145 4.465 1.415 ;
 RECT 4.145 0.665 4.285 1.145 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END Q

 OBS
 LAYER PO ;
 RECT 3.7 1.115 4.03 1.325 ;
 RECT 3.93 0.325 4.03 1.115 ;
 RECT 3.93 1.325 4.03 2.755 ;
 RECT 2.62 0.54 2.72 1.075 ;
 RECT 2.25 1.175 2.35 2.11 ;
 RECT 2.25 1.075 2.72 1.175 ;
 RECT 2.25 2.11 2.49 2.32 ;
 RECT 1.78 0.33 1.88 2.095 ;
 RECT 1.625 2.095 1.88 2.305 ;
 RECT 1.31 0.33 1.41 2.445 ;
 RECT 0.985 2.445 1.41 2.655 ;
 RECT 0.84 0.33 0.94 1.185 ;
 RECT 0.84 1.395 0.94 2.255 ;
 RECT 0.65 1.185 0.94 1.395 ;
 RECT 0.37 0.33 0.47 2.19 ;
 RECT 0.37 2.19 0.635 2.4 ;
 RECT 3.09 0.54 3.19 1.375 ;
 RECT 2.67 1.475 2.77 2.095 ;
 RECT 2.67 1.375 3.19 1.475 ;
 RECT 2.67 2.095 3.07 2.305 ;
 LAYER CO ;
 RECT 3.75 1.155 3.88 1.285 ;
 RECT 4.565 0.655 4.695 0.785 ;
 RECT 4.565 0.395 4.695 0.525 ;
 RECT 4.15 0.725 4.28 0.855 ;
 RECT 4.15 1.625 4.28 1.755 ;
 RECT 4.15 1.885 4.28 2.015 ;
 RECT 4.15 2.405 4.28 2.535 ;
 RECT 4.15 2.145 4.28 2.275 ;
 RECT 3.68 0.56 3.81 0.69 ;
 RECT 3.68 2.145 3.81 2.275 ;
 RECT 3.68 2.405 3.81 2.535 ;
 RECT 2.31 2.15 2.44 2.28 ;
 RECT 1.675 2.135 1.805 2.265 ;
 RECT 1.055 2.485 1.185 2.615 ;
 RECT 0.7 1.225 0.83 1.355 ;
 RECT 0.455 2.23 0.585 2.36 ;
 RECT 3.31 0.76 3.44 0.89 ;
 RECT 2.84 0.76 2.97 0.89 ;
 RECT 2.37 0.76 2.5 0.89 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 1.06 0.55 1.19 0.68 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 0.12 0.55 0.25 0.68 ;
 RECT 2.89 1.64 3.02 1.77 ;
 RECT 2 1.84 2.13 1.97 ;
 RECT 1.06 1.62 1.19 1.75 ;
 RECT 0.12 1.795 0.25 1.925 ;
 RECT 2.89 2.135 3.02 2.265 ;
 RECT 4.645 1.955 4.775 2.085 ;
 RECT 4.645 1.695 4.775 1.825 ;
 RECT 4.645 2.215 4.775 2.345 ;
 LAYER M1 ;
 RECT 1.055 1.29 1.195 1.82 ;
 RECT 2.885 1.29 3.025 1.83 ;
 RECT 2.365 0.69 2.505 1.15 ;
 RECT 3.305 0.7 3.445 1.15 ;
 RECT 3.745 1.105 3.885 1.15 ;
 RECT 3.745 1.29 3.885 1.335 ;
 RECT 1.055 1.15 3.915 1.29 ;
 RECT 2.835 0.36 2.975 0.95 ;
 RECT 1.525 0.22 2.975 0.36 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.495 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 END
END OA222X1

MACRO OA222X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.305 2.27 2.695 2.555 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END IN5

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.65 1.085 0.93 1.415 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END IN2

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.305 2.275 1.625 2.635 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END IN4

 PIN IN6
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.725 1.455 3.035 1.725 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END IN6

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 5.03 1.645 5.17 2.8 ;
 RECT 0.115 2 0.255 2.8 ;
 RECT 1.995 2.015 2.135 2.8 ;
 RECT 3.675 2.095 3.815 2.8 ;
 RECT 4.615 2.095 4.755 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.145 1.42 4.285 2.585 ;
 RECT 4.145 1.16 4.46 1.42 ;
 RECT 4.145 0.7 4.285 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END Q

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.17 1.45 0.47 1.72 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END IN1

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 5.03 0.08 5.17 0.835 ;
 RECT 3.675 0.08 3.815 0.765 ;
 RECT 0.585 0.08 0.725 0.64 ;
 RECT 4.615 0.08 4.755 0.755 ;
 END
 END VSS

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.62 1.455 2.015 1.735 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END IN3

 OBS
 LAYER PO ;
 RECT 0.68 1.085 0.94 1.295 ;
 RECT 0.84 1.295 0.94 2.425 ;
 RECT 0.84 0.24 0.94 1.085 ;
 RECT 1.31 0.24 1.41 2.34 ;
 RECT 1.31 2.34 1.55 2.55 ;
 RECT 1.78 0.24 1.88 1.485 ;
 RECT 1.78 1.695 1.88 2.425 ;
 RECT 1.78 1.485 2.015 1.695 ;
 RECT 2.62 0.365 2.72 1.01 ;
 RECT 2.25 1.11 2.35 2.325 ;
 RECT 2.25 1.01 2.72 1.11 ;
 RECT 2.25 2.325 2.49 2.535 ;
 RECT 3.09 0.36 3.19 1.42 ;
 RECT 2.67 1.675 2.77 2.425 ;
 RECT 2.67 1.52 2.955 1.675 ;
 RECT 2.67 1.42 3.19 1.52 ;
 RECT 3.7 1.23 4.03 1.325 ;
 RECT 3.93 0.345 4.03 1.115 ;
 RECT 4.4 0.345 4.5 1.13 ;
 RECT 4.4 1.23 4.5 2.755 ;
 RECT 3.7 1.115 4.03 1.13 ;
 RECT 3.7 1.13 4.5 1.23 ;
 RECT 3.93 1.325 4.03 2.755 ;
 RECT 0.37 1.715 0.47 2.425 ;
 RECT 0.37 0.24 0.47 1.505 ;
 RECT 0.205 1.505 0.47 1.715 ;
 LAYER CO ;
 RECT 4.62 2.405 4.75 2.535 ;
 RECT 4.62 2.145 4.75 2.275 ;
 RECT 4.62 0.575 4.75 0.705 ;
 RECT 4.15 0.755 4.28 0.885 ;
 RECT 2.89 2.07 3.02 2.2 ;
 RECT 2.37 0.59 2.5 0.72 ;
 RECT 0.12 2.06 0.25 2.19 ;
 RECT 4.15 1.885 4.28 2.015 ;
 RECT 4.15 2.405 4.28 2.535 ;
 RECT 5.035 1.695 5.165 1.825 ;
 RECT 5.035 1.955 5.165 2.085 ;
 RECT 2.775 1.505 2.905 1.635 ;
 RECT 2 2.075 2.13 2.205 ;
 RECT 3.75 1.155 3.88 1.285 ;
 RECT 0.255 1.545 0.385 1.675 ;
 RECT 2.84 0.59 2.97 0.72 ;
 RECT 4.15 1.625 4.28 1.755 ;
 RECT 1.06 1.905 1.19 2.035 ;
 RECT 3.68 0.575 3.81 0.705 ;
 RECT 5.035 0.655 5.165 0.785 ;
 RECT 4.15 2.145 4.28 2.275 ;
 RECT 5.035 2.215 5.165 2.345 ;
 RECT 1.53 0.46 1.66 0.59 ;
 RECT 3.68 2.405 3.81 2.535 ;
 RECT 5.035 0.395 5.165 0.525 ;
 RECT 1.06 0.46 1.19 0.59 ;
 RECT 3.31 0.59 3.44 0.72 ;
 RECT 0.59 0.46 0.72 0.59 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 3.68 2.145 3.81 2.275 ;
 RECT 0.12 0.46 0.25 0.59 ;
 RECT 0.73 1.125 0.86 1.255 ;
 RECT 1.37 2.38 1.5 2.51 ;
 RECT 1.835 1.525 1.965 1.655 ;
 RECT 2.31 2.365 2.44 2.495 ;
 LAYER M1 ;
 RECT 2.835 0.36 2.975 0.775 ;
 RECT 1.525 0.22 2.975 0.36 ;
 RECT 1.525 0.36 1.665 0.64 ;
 RECT 0.115 0.405 0.255 0.78 ;
 RECT 1.055 0.405 1.195 0.78 ;
 RECT 1.995 0.5 2.135 0.78 ;
 RECT 0.115 0.78 2.135 0.92 ;
 RECT 2.365 0.53 2.505 1.06 ;
 RECT 1.07 1.06 3.445 1.15 ;
 RECT 3.305 1.29 3.445 2.065 ;
 RECT 3.305 0.535 3.445 1.06 ;
 RECT 2.84 2.065 3.445 2.205 ;
 RECT 1.07 1.2 1.21 1.61 ;
 RECT 1.055 1.61 1.21 1.79 ;
 RECT 1.055 1.79 1.195 2.135 ;
 RECT 1.07 1.15 3.915 1.2 ;
 RECT 3.305 1.2 3.915 1.29 ;
 RECT 3.745 1.105 3.885 1.15 ;
 RECT 3.745 1.29 3.885 1.335 ;
 END
END OA222X2

MACRO OA22X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.64 2.22 0.92 2.52 ;
 END
 ANTENNAGATEAREA 0.091 ;
 END IN2

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.28 2.12 1.56 2.445 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN4

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 RECT 1.945 1.815 2.695 1.955 ;
 RECT 3.44 1.645 3.58 2.8 ;
 RECT 0.115 1.645 0.255 2.8 ;
 RECT 2.555 1.955 2.695 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.175 1.155 0.46 1.415 ;
 END
 ANTENNAGATEAREA 0.091 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.775 2.12 2.075 2.445 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN3

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.025 1.4 3.165 2.585 ;
 RECT 3.025 1.16 3.355 1.4 ;
 RECT 3.025 0.705 3.165 1.16 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 0.585 0.08 0.725 0.73 ;
 RECT 3.44 0.08 3.58 0.835 ;
 RECT 2.555 0.08 2.695 0.76 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.84 0.33 0.94 2.22 ;
 RECT 0.69 2.22 0.94 2.32 ;
 RECT 0.69 2.32 0.92 2.43 ;
 RECT 1.31 0.33 1.41 2.22 ;
 RECT 1.31 2.22 1.54 2.43 ;
 RECT 2.81 0.35 2.91 1.115 ;
 RECT 2.81 1.325 2.91 2.755 ;
 RECT 2.68 1.115 2.91 1.325 ;
 RECT 1.78 0.33 1.88 2.22 ;
 RECT 1.775 2.22 2.005 2.43 ;
 RECT 0.37 0.33 0.47 1.13 ;
 RECT 0.37 1.34 0.47 2.32 ;
 RECT 0.23 1.13 0.47 1.34 ;
 LAYER CO ;
 RECT 0.12 1.7 0.25 1.83 ;
 RECT 0.74 2.26 0.87 2.39 ;
 RECT 1.36 2.26 1.49 2.39 ;
 RECT 3.445 0.395 3.575 0.525 ;
 RECT 1.825 2.26 1.955 2.39 ;
 RECT 3.445 2.215 3.575 2.345 ;
 RECT 0.28 1.17 0.41 1.3 ;
 RECT 3.03 0.76 3.16 0.89 ;
 RECT 2.56 2.145 2.69 2.275 ;
 RECT 0.12 1.96 0.25 2.09 ;
 RECT 3.03 1.625 3.16 1.755 ;
 RECT 3.03 2.405 3.16 2.535 ;
 RECT 3.03 2.145 3.16 2.275 ;
 RECT 3.03 1.885 3.16 2.015 ;
 RECT 1.06 1.5 1.19 1.63 ;
 RECT 3.445 1.955 3.575 2.085 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 2.73 1.155 2.86 1.285 ;
 RECT 3.445 1.695 3.575 1.825 ;
 RECT 1.06 0.55 1.19 0.68 ;
 RECT 2.56 0.58 2.69 0.71 ;
 RECT 2.56 2.405 2.69 2.535 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 2 1.82 2.13 1.95 ;
 RECT 0.12 0.55 0.25 0.68 ;
 RECT 3.445 0.655 3.575 0.785 ;
 LAYER M1 ;
 RECT 2.275 0.36 2.415 1.15 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 1.525 0.22 2.415 0.36 ;
 RECT 1.055 1.29 1.195 1.69 ;
 RECT 2.725 1.105 2.865 1.15 ;
 RECT 2.725 1.29 2.865 1.335 ;
 RECT 1.055 1.15 2.88 1.29 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.495 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 END
END OA22X1

MACRO OA22X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 3.91 1.645 4.05 2.8 ;
 RECT 1.995 2.06 2.135 2.8 ;
 RECT 0.115 2.07 0.255 2.8 ;
 RECT 2.555 2.095 2.695 2.8 ;
 RECT 3.495 2.095 3.635 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.175 1.48 0.44 1.755 ;
 END
 ANTENNAGATEAREA 0.091 ;
 END IN1

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.025 1.4 3.165 2.585 ;
 RECT 3.025 1.16 3.48 1.4 ;
 RECT 3.025 0.685 3.165 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END Q

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.95 1.475 2.29 1.72 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 3.91 0.08 4.05 0.835 ;
 RECT 0.585 0.08 0.725 0.73 ;
 RECT 2.555 0.08 2.695 0.765 ;
 RECT 3.495 0.08 3.635 0.77 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.655 1.32 0.92 1.59 ;
 END
 ANTENNAGATEAREA 0.091 ;
 END IN2

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.345 1.625 1.735 1.905 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN4

 OBS
 LAYER PO ;
 RECT 3.28 0.335 3.38 1.125 ;
 RECT 3.28 1.225 3.38 2.755 ;
 RECT 2.68 1.115 2.91 1.125 ;
 RECT 2.68 1.225 2.91 1.325 ;
 RECT 2.68 1.125 3.38 1.225 ;
 RECT 2.81 1.325 2.91 2.755 ;
 RECT 2.81 0.335 2.91 1.115 ;
 RECT 1.31 1.905 1.41 2.745 ;
 RECT 1.31 0.33 1.41 1.695 ;
 RECT 1.31 1.695 1.575 1.905 ;
 RECT 1.78 0.33 1.88 1.485 ;
 RECT 1.78 1.695 1.88 2.745 ;
 RECT 1.78 1.485 2.195 1.695 ;
 RECT 0.37 0.33 0.47 1.535 ;
 RECT 0.37 1.745 0.47 2.745 ;
 RECT 0.205 1.535 0.47 1.745 ;
 RECT 0.84 0.33 0.94 1.37 ;
 RECT 0.84 1.58 0.94 2.745 ;
 RECT 0.7 1.37 0.94 1.58 ;
 LAYER CO ;
 RECT 2 2.115 2.13 2.245 ;
 RECT 1.06 2.085 1.19 2.215 ;
 RECT 0.12 2.125 0.25 2.255 ;
 RECT 3.5 2.405 3.63 2.535 ;
 RECT 3.5 2.145 3.63 2.275 ;
 RECT 3.5 0.575 3.63 0.705 ;
 RECT 3.915 2.215 4.045 2.345 ;
 RECT 3.915 0.655 4.045 0.785 ;
 RECT 3.915 1.955 4.045 2.085 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 2.56 2.405 2.69 2.535 ;
 RECT 2.73 1.155 2.86 1.285 ;
 RECT 1.395 1.735 1.525 1.865 ;
 RECT 0.75 1.41 0.88 1.54 ;
 RECT 2 2.375 2.13 2.505 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 0.12 0.55 0.25 0.68 ;
 RECT 2.015 1.525 2.145 1.655 ;
 RECT 0.255 1.575 0.385 1.705 ;
 RECT 3.03 1.595 3.16 1.725 ;
 RECT 1.06 0.55 1.19 0.68 ;
 RECT 3.03 2.115 3.16 2.245 ;
 RECT 3.03 1.855 3.16 1.985 ;
 RECT 2.56 0.575 2.69 0.705 ;
 RECT 3.03 2.375 3.16 2.505 ;
 RECT 3.03 0.745 3.16 0.875 ;
 RECT 3.915 0.395 4.045 0.525 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 2.56 2.145 2.69 2.275 ;
 RECT 3.915 1.695 4.045 1.825 ;
 RECT 1.06 2.345 1.19 2.475 ;
 RECT 0.12 2.385 0.25 2.515 ;
 LAYER M1 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.495 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 RECT 2.275 0.36 2.415 1.15 ;
 RECT 1.525 0.22 2.415 0.36 ;
 RECT 1.06 1.29 1.2 1.645 ;
 RECT 1.055 1.645 1.2 1.785 ;
 RECT 1.055 1.785 1.195 2.535 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 1.06 1.15 2.865 1.29 ;
 RECT 2.725 1.105 2.865 1.15 ;
 RECT 2.725 1.29 2.865 1.335 ;
 END
END OA22X2

MACRO OAI21X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.17 1.35 0.46 1.755 ;
 END
 ANTENNAGATEAREA 0.062 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 RECT 0.115 1.915 0.255 2.8 ;
 RECT 3.25 1.645 3.39 2.8 ;
 RECT 1.525 1.88 1.665 2.8 ;
 RECT 2.365 2.095 2.505 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 2.365 0.08 2.505 0.905 ;
 RECT 0.585 0.08 0.725 0.74 ;
 RECT 3.25 0.08 3.39 0.835 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.835 1.4 2.975 2.585 ;
 RECT 2.835 1.16 3.195 1.4 ;
 RECT 2.835 0.705 2.975 1.16 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END QN

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.335 1.48 1.745 1.72 ;
 END
 ANTENNAGATEAREA 0.053 ;
 END IN3

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.66 2.265 0.92 2.63 ;
 END
 ANTENNAGATEAREA 0.062 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 0.84 0.33 0.94 2.4 ;
 RECT 0.71 2.4 0.94 2.61 ;
 RECT 1.31 0.33 1.41 1.495 ;
 RECT 1.31 1.705 1.41 2.28 ;
 RECT 1.31 1.495 1.55 1.705 ;
 RECT 2.47 1.085 2.72 1.295 ;
 RECT 2.62 1.295 2.72 2.755 ;
 RECT 2.62 0.325 2.72 1.085 ;
 RECT 0.37 0.33 0.47 1.535 ;
 RECT 0.37 1.745 0.47 2.5 ;
 RECT 0.205 1.535 0.47 1.745 ;
 RECT 2.15 0.505 2.25 2.185 ;
 RECT 2.02 0.295 2.25 0.505 ;
 LAYER CO ;
 RECT 0.12 1.97 0.25 2.1 ;
 RECT 2.37 2.145 2.5 2.275 ;
 RECT 1.53 1.93 1.66 2.06 ;
 RECT 0.76 2.44 0.89 2.57 ;
 RECT 1.06 0.56 1.19 0.69 ;
 RECT 3.255 0.395 3.385 0.525 ;
 RECT 2.37 2.405 2.5 2.535 ;
 RECT 2.84 2.405 2.97 2.535 ;
 RECT 2.07 0.335 2.2 0.465 ;
 RECT 2.52 1.125 2.65 1.255 ;
 RECT 1.9 0.765 2.03 0.895 ;
 RECT 0.255 1.575 0.385 1.705 ;
 RECT 2.37 0.725 2.5 0.855 ;
 RECT 1.37 1.535 1.5 1.665 ;
 RECT 2.84 1.625 2.97 1.755 ;
 RECT 2.84 1.885 2.97 2.015 ;
 RECT 3.255 1.695 3.385 1.825 ;
 RECT 0.12 0.56 0.25 0.69 ;
 RECT 3.255 0.655 3.385 0.785 ;
 RECT 0.59 0.56 0.72 0.69 ;
 RECT 1.9 1.52 2.03 1.65 ;
 RECT 2.84 2.145 2.97 2.275 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 1.06 1.925 1.19 2.055 ;
 RECT 3.255 1.955 3.385 2.085 ;
 RECT 2.84 0.755 2.97 0.885 ;
 RECT 3.255 2.215 3.385 2.345 ;
 LAYER M1 ;
 RECT 0.115 0.51 0.255 0.9 ;
 RECT 1.055 0.5 1.195 0.9 ;
 RECT 0.115 0.9 1.195 1.04 ;
 RECT 1.055 1.33 1.195 2.105 ;
 RECT 2.065 0.285 2.205 0.33 ;
 RECT 2.065 0.47 2.205 0.515 ;
 RECT 1.525 0.47 1.665 1.19 ;
 RECT 1.055 1.19 1.665 1.33 ;
 RECT 1.525 0.33 2.21 0.47 ;
 RECT 1.895 0.705 2.035 1.12 ;
 RECT 1.895 1.26 2.035 1.705 ;
 RECT 2.515 1.075 2.655 1.12 ;
 RECT 2.515 1.26 2.655 1.305 ;
 RECT 1.895 1.12 2.655 1.26 ;
 END
END OAI21X1

MACRO OAI21X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.17 1.43 0.465 1.755 ;
 END
 ANTENNAGATEAREA 0.062 ;
 END IN1

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.835 1.4 2.975 2.585 ;
 RECT 2.835 1.16 3.19 1.4 ;
 RECT 2.835 0.705 2.975 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END QN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 3.72 0.08 3.86 0.835 ;
 RECT 2.365 0.08 2.505 0.905 ;
 RECT 3.305 0.08 3.445 0.905 ;
 RECT 0.585 0.08 0.725 0.705 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 3.305 2.095 3.445 2.8 ;
 RECT 3.72 1.645 3.86 2.8 ;
 RECT 2.365 2.095 2.505 2.8 ;
 RECT 0.115 2.055 0.255 2.8 ;
 RECT 1.525 1.86 1.665 2.8 ;
 END
 END VDD

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.365 1.455 1.735 1.72 ;
 END
 ANTENNAGATEAREA 0.053 ;
 END IN3

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.645 2.26 0.96 2.62 ;
 END
 ANTENNAGATEAREA 0.062 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 2.62 0.325 2.72 1.085 ;
 RECT 2.62 1.295 2.72 2.755 ;
 RECT 3.09 1.25 3.19 2.755 ;
 RECT 2.47 1.085 2.72 1.15 ;
 RECT 2.47 1.15 3.19 1.25 ;
 RECT 2.47 1.25 2.72 1.295 ;
 RECT 3.09 0.325 3.19 1.15 ;
 RECT 1.31 0.33 1.41 1.495 ;
 RECT 1.31 1.705 1.41 2.26 ;
 RECT 1.31 1.495 1.55 1.705 ;
 RECT 2.15 0.555 2.25 2.185 ;
 RECT 2.02 0.345 2.25 0.555 ;
 RECT 0.37 0.385 0.47 1.535 ;
 RECT 0.37 1.745 0.47 2.51 ;
 RECT 0.205 1.535 0.47 1.745 ;
 RECT 0.84 0.385 0.94 2.41 ;
 RECT 0.7 2.41 0.94 2.62 ;
 LAYER CO ;
 RECT 3.725 0.655 3.855 0.785 ;
 RECT 3.725 2.215 3.855 2.345 ;
 RECT 3.725 0.395 3.855 0.525 ;
 RECT 3.31 2.405 3.44 2.535 ;
 RECT 2.84 1.625 2.97 1.755 ;
 RECT 2.52 1.125 2.65 1.255 ;
 RECT 2.07 0.385 2.2 0.515 ;
 RECT 3.725 1.695 3.855 1.825 ;
 RECT 1.37 1.535 1.5 1.665 ;
 RECT 2.37 2.145 2.5 2.275 ;
 RECT 3.725 1.955 3.855 2.085 ;
 RECT 2.84 2.405 2.97 2.535 ;
 RECT 1.53 1.91 1.66 2.04 ;
 RECT 2.37 0.725 2.5 0.855 ;
 RECT 2.84 0.755 2.97 0.885 ;
 RECT 1.9 1.52 2.03 1.65 ;
 RECT 2.84 2.145 2.97 2.275 ;
 RECT 1.06 0.64 1.19 0.77 ;
 RECT 1.9 0.765 2.03 0.895 ;
 RECT 0.59 0.525 0.72 0.655 ;
 RECT 0.255 1.575 0.385 1.705 ;
 RECT 3.31 0.725 3.44 0.855 ;
 RECT 0.75 2.45 0.88 2.58 ;
 RECT 0.12 0.525 0.25 0.655 ;
 RECT 1.06 1.9 1.19 2.03 ;
 RECT 0.12 2.11 0.25 2.24 ;
 RECT 2.37 2.405 2.5 2.535 ;
 RECT 2.84 1.885 2.97 2.015 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 3.31 2.145 3.44 2.275 ;
 LAYER M1 ;
 RECT 1.895 0.705 2.035 1.12 ;
 RECT 1.895 1.26 2.035 1.705 ;
 RECT 2.515 1.075 2.655 1.12 ;
 RECT 2.515 1.26 2.655 1.305 ;
 RECT 1.895 1.12 2.655 1.26 ;
 RECT 0.115 0.475 0.255 0.87 ;
 RECT 1.055 0.59 1.195 0.87 ;
 RECT 0.115 0.87 1.195 1.01 ;
 RECT 1.055 1.29 1.195 2.12 ;
 RECT 2.065 0.335 2.205 0.38 ;
 RECT 2.065 0.52 2.205 0.565 ;
 RECT 1.525 0.52 1.665 1.15 ;
 RECT 1.525 0.38 2.21 0.52 ;
 RECT 1.055 1.15 1.665 1.29 ;
 END
END OAI21X2

MACRO OAI221X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.655 2.095 0.95 2.48 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN2

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 3.675 2.095 3.815 2.8 ;
 RECT 1.995 1.82 2.135 2.8 ;
 RECT 4.56 1.645 4.7 2.8 ;
 RECT 0.115 1.82 0.255 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 4.56 0.08 4.7 0.835 ;
 RECT 3.675 0.08 3.815 0.905 ;
 RECT 0.585 0.08 0.725 0.705 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.145 1.4 4.285 2.585 ;
 RECT 4.145 1.16 4.475 1.4 ;
 RECT 4.145 0.705 4.285 1.16 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END QN

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.275 1.055 2.555 1.4 ;
 END
 ANTENNAGATEAREA 0.046 ;
 END IN5

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.235 1.155 1.58 1.4 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN4

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.45 2.095 1.835 2.385 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN3

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.17 1.15 0.475 1.475 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 0.84 0.33 0.94 2.16 ;
 RECT 0.71 2.16 0.94 2.37 ;
 RECT 1.78 0.33 1.88 2.14 ;
 RECT 1.645 2.14 1.88 2.35 ;
 RECT 3.46 0.615 3.56 1.905 ;
 RECT 3.31 1.905 3.56 2.065 ;
 RECT 3.31 2.065 3.54 2.115 ;
 RECT 3.93 1.295 4.03 2.755 ;
 RECT 3.93 0.325 4.03 1.085 ;
 RECT 3.78 1.085 4.03 1.295 ;
 RECT 1.31 0.33 1.41 1.175 ;
 RECT 1.31 1.385 1.41 2.235 ;
 RECT 1.31 1.175 1.55 1.385 ;
 RECT 0.37 1.39 0.47 2.235 ;
 RECT 0.37 0.33 0.47 1.18 ;
 RECT 0.235 1.18 0.47 1.39 ;
 RECT 2.25 1.275 2.35 2.235 ;
 RECT 2.62 0.49 2.72 1.055 ;
 RECT 2.25 1.155 2.49 1.275 ;
 RECT 2.25 1.055 2.72 1.155 ;
 LAYER CO ;
 RECT 1.06 0.55 1.19 0.68 ;
 RECT 4.565 2.215 4.695 2.345 ;
 RECT 4.15 2.145 4.28 2.275 ;
 RECT 4.15 1.885 4.28 2.015 ;
 RECT 4.15 1.625 4.28 1.755 ;
 RECT 3.68 0.725 3.81 0.855 ;
 RECT 0.12 0.525 0.25 0.655 ;
 RECT 1.695 2.18 1.825 2.31 ;
 RECT 2.37 0.72 2.5 0.85 ;
 RECT 2.31 1.105 2.44 1.235 ;
 RECT 2 1.875 2.13 2.005 ;
 RECT 4.15 0.755 4.28 0.885 ;
 RECT 0.12 1.88 0.25 2.01 ;
 RECT 4.15 2.405 4.28 2.535 ;
 RECT 3.21 1.52 3.34 1.65 ;
 RECT 1.06 1.725 1.19 1.855 ;
 RECT 2.84 0.72 2.97 0.85 ;
 RECT 3.21 0.755 3.34 0.885 ;
 RECT 1.37 1.215 1.5 1.345 ;
 RECT 4.565 1.955 4.695 2.085 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 0.59 0.525 0.72 0.655 ;
 RECT 0.285 1.22 0.415 1.35 ;
 RECT 3.68 2.145 3.81 2.275 ;
 RECT 3.36 1.945 3.49 2.075 ;
 RECT 3.83 1.125 3.96 1.255 ;
 RECT 4.565 1.695 4.695 1.825 ;
 RECT 2.475 1.885 2.605 2.015 ;
 RECT 0.76 2.2 0.89 2.33 ;
 RECT 4.565 0.655 4.695 0.785 ;
 RECT 3.68 2.405 3.81 2.535 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 4.565 0.395 4.695 0.525 ;
 LAYER M1 ;
 RECT 3.205 0.705 3.345 1.12 ;
 RECT 3.205 1.26 3.345 1.705 ;
 RECT 3.825 1.075 3.965 1.12 ;
 RECT 3.825 1.26 3.965 1.305 ;
 RECT 3.205 1.12 3.965 1.26 ;
 RECT 0.115 0.475 0.255 0.87 ;
 RECT 1.055 0.485 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 RECT 2.365 0.36 2.505 0.905 ;
 RECT 1.525 0.22 2.505 0.36 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 1.055 1.68 1.195 1.915 ;
 RECT 2.47 1.68 2.61 1.94 ;
 RECT 2.47 1.94 3.52 2.08 ;
 RECT 3.355 1.895 3.495 1.94 ;
 RECT 3.355 2.08 3.495 2.125 ;
 RECT 2.835 0.66 2.975 1.54 ;
 RECT 1.055 1.54 2.975 1.68 ;
 END
END OAI221X1

MACRO OAI221X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 3.675 0.08 3.815 0.735 ;
 RECT 5.03 0.08 5.17 0.835 ;
 RECT 0.585 0.08 0.725 0.73 ;
 RECT 4.615 0.08 4.755 0.905 ;
 END
 END VSS

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.25 1.46 2.605 1.72 ;
 END
 ANTENNAGATEAREA 0.046 ;
 END IN5

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.59 1.465 1.915 1.72 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN3

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.285 2.25 1.59 2.55 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN4

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.165 1.455 0.465 1.73 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN1

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.145 1.4 4.285 2.585 ;
 RECT 4.145 1.16 4.48 1.4 ;
 RECT 4.145 0.705 4.285 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 3.675 2.095 3.815 2.8 ;
 RECT 1.995 1.92 2.135 2.8 ;
 RECT 0.115 1.915 0.255 2.8 ;
 RECT 5.03 1.645 5.17 2.8 ;
 RECT 4.615 2.095 4.755 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.575 2.265 0.945 2.55 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 1.78 0.33 1.88 1.485 ;
 RECT 1.78 1.695 1.88 2.375 ;
 RECT 1.62 1.485 1.88 1.695 ;
 RECT 1.31 0.33 1.41 2.275 ;
 RECT 1.31 2.275 1.55 2.485 ;
 RECT 3.46 0.615 3.56 1.91 ;
 RECT 3.31 1.91 3.56 2.065 ;
 RECT 3.31 2.065 3.54 2.12 ;
 RECT 0.37 0.33 0.47 1.48 ;
 RECT 0.37 1.69 0.47 2.375 ;
 RECT 0.205 1.48 0.47 1.69 ;
 RECT 2.62 0.495 2.72 1.055 ;
 RECT 2.25 1.68 2.35 2.375 ;
 RECT 2.25 1.155 2.35 1.47 ;
 RECT 2.25 1.47 2.49 1.68 ;
 RECT 2.25 1.055 2.72 1.155 ;
 RECT 0.84 0.33 0.94 2.275 ;
 RECT 0.7 2.275 0.94 2.485 ;
 RECT 3.93 0.325 4.03 1.085 ;
 RECT 3.93 1.295 4.03 2.755 ;
 RECT 4.4 1.25 4.5 2.755 ;
 RECT 3.78 1.085 4.03 1.15 ;
 RECT 3.78 1.15 4.5 1.25 ;
 RECT 3.78 1.25 4.03 1.295 ;
 RECT 4.4 0.325 4.5 1.15 ;
 LAYER CO ;
 RECT 4.62 0.725 4.75 0.855 ;
 RECT 4.62 2.405 4.75 2.535 ;
 RECT 4.62 2.145 4.75 2.275 ;
 RECT 0.75 2.315 0.88 2.445 ;
 RECT 5.035 1.695 5.165 1.825 ;
 RECT 5.035 0.655 5.165 0.785 ;
 RECT 5.035 0.395 5.165 0.525 ;
 RECT 5.035 2.215 5.165 2.345 ;
 RECT 5.035 1.955 5.165 2.085 ;
 RECT 4.15 1.625 4.28 1.755 ;
 RECT 3.21 0.755 3.34 0.885 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 2.31 1.51 2.44 1.64 ;
 RECT 4.15 2.145 4.28 2.275 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 1.67 1.525 1.8 1.655 ;
 RECT 3.68 0.555 3.81 0.685 ;
 RECT 2.84 0.73 2.97 0.86 ;
 RECT 1.06 1.875 1.19 2.005 ;
 RECT 2.37 0.73 2.5 0.86 ;
 RECT 4.15 0.755 4.28 0.885 ;
 RECT 2 1.975 2.13 2.105 ;
 RECT 0.12 1.975 0.25 2.105 ;
 RECT 3.36 1.95 3.49 2.08 ;
 RECT 0.255 1.52 0.385 1.65 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 4.15 2.405 4.28 2.535 ;
 RECT 3.21 1.52 3.34 1.65 ;
 RECT 1.06 0.56 1.19 0.69 ;
 RECT 3.68 2.145 3.81 2.275 ;
 RECT 3.83 1.125 3.96 1.255 ;
 RECT 4.15 1.885 4.28 2.015 ;
 RECT 2.475 2.025 2.605 2.155 ;
 RECT 0.12 0.56 0.25 0.69 ;
 RECT 3.68 2.405 3.81 2.535 ;
 RECT 1.37 2.315 1.5 2.445 ;
 LAYER M1 ;
 RECT 2.365 0.36 2.505 0.91 ;
 RECT 1.525 0.22 2.505 0.36 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.51 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 RECT 3.205 0.705 3.345 1.12 ;
 RECT 3.205 1.26 3.345 1.705 ;
 RECT 3.825 1.075 3.965 1.12 ;
 RECT 3.825 1.26 3.965 1.305 ;
 RECT 3.205 1.12 3.965 1.26 ;
 RECT 1.055 1.29 1.195 2.065 ;
 RECT 3.355 2.09 3.495 2.13 ;
 RECT 2.84 1.95 3.52 2.02 ;
 RECT 2.84 1.29 2.98 1.95 ;
 RECT 3.355 1.9 3.495 1.95 ;
 RECT 1.055 1.15 2.98 1.29 ;
 RECT 2.425 2.02 3.52 2.09 ;
 RECT 2.425 2.09 2.98 2.16 ;
 RECT 2.835 0.665 2.975 1.15 ;
 END
END OAI221X2

MACRO OAI222X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.49 2.095 0.88 2.515 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END IN2

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.235 1.43 2.555 1.72 ;
 END
 ANTENNAGATEAREA 0.035 ;
 END IN5

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 1.995 1.86 2.135 2.8 ;
 RECT 0.115 1.84 0.255 2.8 ;
 RECT 4.145 2.095 4.285 2.8 ;
 RECT 5.03 1.645 5.17 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 5.03 0.08 5.17 0.835 ;
 RECT 4.145 0.08 4.285 0.75 ;
 RECT 0.585 0.08 0.725 0.73 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.615 1.41 4.755 2.585 ;
 RECT 4.615 1.11 5.105 1.41 ;
 RECT 4.615 0.705 4.755 1.11 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END QN

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.35 1.44 1.75 1.735 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END IN4

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.46 2.11 1.855 2.41 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END IN3

 PIN IN6
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.57 2.2 2.935 2.55 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END IN6

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.12 1.16 0.465 1.435 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 4.4 0.325 4.5 1.085 ;
 RECT 4.4 1.295 4.5 2.755 ;
 RECT 4.25 1.085 4.5 1.295 ;
 RECT 1.31 1.44 1.58 1.65 ;
 RECT 1.31 1.65 1.41 2.265 ;
 RECT 1.31 0.41 1.41 1.44 ;
 RECT 0.37 0.41 0.47 1.215 ;
 RECT 0.37 1.425 0.47 2.265 ;
 RECT 0.205 1.215 0.47 1.425 ;
 RECT 3.93 0.615 4.03 1.905 ;
 RECT 3.78 1.905 4.03 2.07 ;
 RECT 3.78 2.07 4.01 2.115 ;
 RECT 2.67 1.52 2.77 2.2 ;
 RECT 3.09 0.64 3.19 1.42 ;
 RECT 2.67 1.42 3.19 1.52 ;
 RECT 2.67 2.2 2.9 2.41 ;
 RECT 1.78 0.41 1.88 2.17 ;
 RECT 1.65 2.17 1.88 2.38 ;
 RECT 2.25 1.24 2.35 1.44 ;
 RECT 2.25 1.44 2.49 1.65 ;
 RECT 2.25 1.65 2.35 2.175 ;
 RECT 2.62 0.64 2.72 1.14 ;
 RECT 2.25 1.14 2.72 1.24 ;
 RECT 0.84 0.41 0.94 2.195 ;
 RECT 0.65 2.195 0.94 2.405 ;
 LAYER CO ;
 RECT 1.4 1.48 1.53 1.61 ;
 RECT 5.035 0.655 5.165 0.785 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 4.3 1.125 4.43 1.255 ;
 RECT 4.62 2.405 4.75 2.535 ;
 RECT 4.62 2.145 4.75 2.275 ;
 RECT 4.62 0.755 4.75 0.885 ;
 RECT 4.62 1.885 4.75 2.015 ;
 RECT 4.62 1.625 4.75 1.755 ;
 RECT 0.255 1.255 0.385 1.385 ;
 RECT 5.035 0.395 5.165 0.525 ;
 RECT 0.12 0.55 0.25 0.68 ;
 RECT 4.15 0.565 4.28 0.695 ;
 RECT 1.06 1.825 1.19 1.955 ;
 RECT 2.72 2.24 2.85 2.37 ;
 RECT 2.84 0.78 2.97 0.91 ;
 RECT 4.15 2.405 4.28 2.535 ;
 RECT 1.7 2.21 1.83 2.34 ;
 RECT 5.035 2.215 5.165 2.345 ;
 RECT 2.31 1.48 2.44 1.61 ;
 RECT 0.12 1.9 0.25 2.03 ;
 RECT 3.83 1.945 3.96 2.075 ;
 RECT 3.68 0.755 3.81 0.885 ;
 RECT 0.7 2.235 0.83 2.365 ;
 RECT 2 1.91 2.13 2.04 ;
 RECT 4.15 2.145 4.28 2.275 ;
 RECT 5.035 1.695 5.165 1.825 ;
 RECT 3.31 0.78 3.44 0.91 ;
 RECT 3.68 1.52 3.81 1.65 ;
 RECT 2.37 0.78 2.5 0.91 ;
 RECT 5.035 1.955 5.165 2.085 ;
 RECT 2.89 1.865 3.02 1.995 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 1.06 0.55 1.19 0.68 ;
 LAYER M1 ;
 RECT 2.835 0.36 2.975 0.96 ;
 RECT 1.525 0.22 2.975 0.36 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 3.675 0.705 3.815 1.12 ;
 RECT 3.675 1.26 3.815 1.705 ;
 RECT 4.295 1.075 4.435 1.12 ;
 RECT 4.295 1.26 4.435 1.305 ;
 RECT 3.675 1.12 4.435 1.26 ;
 RECT 1.055 1.29 1.195 2.005 ;
 RECT 3.825 1.895 3.965 1.94 ;
 RECT 3.825 2.08 3.965 2.125 ;
 RECT 2.365 0.73 2.505 1.15 ;
 RECT 3.305 1.29 3.445 1.86 ;
 RECT 2.84 1.94 3.98 2 ;
 RECT 2.84 1.86 3.445 1.94 ;
 RECT 3.305 2 3.98 2.08 ;
 RECT 3.305 0.725 3.445 1.15 ;
 RECT 1.055 1.15 3.445 1.29 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.495 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 END
END OAI222X1

MACRO OAI222X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.08 BY 2.88 ;
 PIN IN6
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.58 1.45 2.88 1.76 ;
 END
 ANTENNAGATEAREA 0.039 ;
 END IN6

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.56 1.16 4.955 1.425 ;
 RECT 4.615 1.425 4.755 2.585 ;
 RECT 4.615 0.705 4.755 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END QN

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.275 2.105 2.555 2.445 ;
 END
 ANTENNAGATEAREA 0.039 ;
 END IN5

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.365 1.455 1.75 1.745 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END IN4

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.45 2.12 1.855 2.405 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.08 0.08 ;
 RECT 5.5 0.08 5.64 0.835 ;
 RECT 0.585 0.08 0.725 0.73 ;
 RECT 4.145 0.08 4.285 0.83 ;
 RECT 5.085 0.08 5.225 0.83 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.16 0.475 1.435 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.495 2.185 0.94 2.425 ;
 END
 ANTENNAGATEAREA 0.044 ;
 END IN2

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.08 2.96 ;
 RECT 4.145 2.095 4.285 2.8 ;
 RECT 5.5 1.645 5.64 2.8 ;
 RECT 0.115 1.835 0.255 2.8 ;
 RECT 1.995 1.87 2.135 2.8 ;
 RECT 5.085 2.095 5.225 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 2.62 0.555 2.72 1.055 ;
 RECT 2.62 1.155 2.72 1.165 ;
 RECT 2.25 1.155 2.35 2.195 ;
 RECT 2.25 1.055 2.72 1.155 ;
 RECT 2.25 2.195 2.49 2.405 ;
 RECT 2.67 1.67 2.77 2.295 ;
 RECT 3.09 0.555 3.19 1.42 ;
 RECT 2.67 1.52 2.9 1.67 ;
 RECT 2.67 1.42 3.19 1.52 ;
 RECT 3.93 0.615 4.03 1.905 ;
 RECT 3.78 1.905 4.03 2.065 ;
 RECT 3.78 2.065 4.01 2.115 ;
 RECT 4.4 0.325 4.5 1.085 ;
 RECT 4.4 1.295 4.5 2.755 ;
 RECT 4.87 1.25 4.97 2.755 ;
 RECT 4.225 1.085 4.5 1.15 ;
 RECT 4.225 1.15 4.97 1.25 ;
 RECT 4.225 1.25 4.5 1.295 ;
 RECT 4.87 0.325 4.97 1.15 ;
 RECT 1.31 1.495 1.55 1.705 ;
 RECT 1.31 1.705 1.41 2.295 ;
 RECT 1.31 0.41 1.41 1.495 ;
 RECT 0.37 1.425 0.47 2.295 ;
 RECT 0.37 0.41 0.47 1.215 ;
 RECT 0.205 1.215 0.47 1.425 ;
 RECT 0.84 0.41 0.94 2.195 ;
 RECT 0.7 2.195 0.94 2.405 ;
 RECT 1.78 0.41 1.88 2.195 ;
 RECT 1.59 2.195 1.88 2.405 ;
 LAYER CO ;
 RECT 4.62 1.885 4.75 2.015 ;
 RECT 4.62 1.625 4.75 1.755 ;
 RECT 0.12 1.895 0.25 2.025 ;
 RECT 5.09 0.64 5.22 0.77 ;
 RECT 5.09 2.405 5.22 2.535 ;
 RECT 5.09 2.145 5.22 2.275 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 3.68 0.755 3.81 0.885 ;
 RECT 2.89 1.945 3.02 2.075 ;
 RECT 5.505 1.695 5.635 1.825 ;
 RECT 0.75 2.235 0.88 2.365 ;
 RECT 4.62 2.405 4.75 2.535 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 5.505 0.655 5.635 0.785 ;
 RECT 5.505 0.395 5.635 0.525 ;
 RECT 4.15 2.145 4.28 2.275 ;
 RECT 3.83 1.945 3.96 2.075 ;
 RECT 4.275 1.125 4.405 1.255 ;
 RECT 4.15 0.64 4.28 0.77 ;
 RECT 3.31 0.695 3.44 0.825 ;
 RECT 0.12 0.55 0.25 0.68 ;
 RECT 4.15 2.405 4.28 2.535 ;
 RECT 2.31 2.235 2.44 2.365 ;
 RECT 1.64 2.235 1.77 2.365 ;
 RECT 2.37 0.695 2.5 0.825 ;
 RECT 2 1.93 2.13 2.06 ;
 RECT 4.62 0.755 4.75 0.885 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 2.72 1.5 2.85 1.63 ;
 RECT 3.68 1.52 3.81 1.65 ;
 RECT 1.06 1.855 1.19 1.985 ;
 RECT 0.255 1.255 0.385 1.385 ;
 RECT 1.06 0.55 1.19 0.68 ;
 RECT 1.37 1.535 1.5 1.665 ;
 RECT 5.505 2.215 5.635 2.345 ;
 RECT 4.62 2.145 4.75 2.275 ;
 RECT 5.505 1.955 5.635 2.085 ;
 RECT 2.84 0.695 2.97 0.825 ;
 LAYER M1 ;
 RECT 2.835 0.36 2.975 0.875 ;
 RECT 1.525 0.22 2.975 0.36 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 3.675 0.705 3.815 1.12 ;
 RECT 3.675 1.26 3.815 1.705 ;
 RECT 4.27 1.075 4.41 1.12 ;
 RECT 4.27 1.26 4.41 1.305 ;
 RECT 3.675 1.12 4.42 1.26 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.5 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 RECT 1.055 1.29 1.195 2.035 ;
 RECT 2.365 0.645 2.505 1.15 ;
 RECT 3.305 1.29 3.445 1.94 ;
 RECT 2.84 1.94 3.98 2.08 ;
 RECT 3.825 1.895 3.965 1.94 ;
 RECT 3.825 2.08 3.965 2.125 ;
 RECT 3.305 0.645 3.445 1.15 ;
 RECT 1.055 1.15 3.445 1.29 ;
 END
END OAI222X2

MACRO OAI22X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.45 2.085 1.85 2.405 ;
 END
 ANTENNAGATEAREA 0.073 ;
 END IN3

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.495 1.4 3.635 2.585 ;
 RECT 3.495 1.15 3.835 1.4 ;
 RECT 3.495 0.705 3.635 1.15 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END QN

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.095 1.16 0.475 1.485 ;
 END
 ANTENNAGATEAREA 0.064 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 0.115 1.845 0.255 2.8 ;
 RECT 3.91 1.645 4.05 2.8 ;
 RECT 1.995 1.835 2.135 2.8 ;
 RECT 3.025 2.095 3.165 2.8 ;
 END
 END VDD

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.265 1.15 1.595 1.405 ;
 END
 ANTENNAGATEAREA 0.073 ;
 END IN4

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.66 2.095 0.95 2.425 ;
 END
 ANTENNAGATEAREA 0.064 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 3.91 0.08 4.05 0.835 ;
 RECT 3.025 0.08 3.165 0.905 ;
 RECT 0.585 0.08 0.725 0.73 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.37 0.41 0.47 1.215 ;
 RECT 0.37 1.425 0.47 2.26 ;
 RECT 0.205 1.215 0.47 1.425 ;
 RECT 1.31 0.32 1.41 1.175 ;
 RECT 1.31 1.385 1.41 2.26 ;
 RECT 1.31 1.175 1.55 1.385 ;
 RECT 3.13 1.085 3.38 1.295 ;
 RECT 3.28 1.295 3.38 2.755 ;
 RECT 3.28 0.295 3.38 1.085 ;
 RECT 2.81 0.555 2.91 2.035 ;
 RECT 2.675 0.455 2.91 0.555 ;
 RECT 2.675 0.345 2.905 0.455 ;
 RECT 1.78 0.32 1.88 2.18 ;
 RECT 1.62 2.18 1.88 2.26 ;
 RECT 1.62 2.26 1.85 2.39 ;
 RECT 0.84 0.41 0.94 2.16 ;
 RECT 0.7 2.16 0.94 2.37 ;
 LAYER CO ;
 RECT 3.5 2.405 3.63 2.535 ;
 RECT 3.03 0.725 3.16 0.855 ;
 RECT 3.915 0.655 4.045 0.785 ;
 RECT 1.06 1.725 1.19 1.855 ;
 RECT 2 1.89 2.13 2.02 ;
 RECT 1.37 1.215 1.5 1.345 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 0.12 1.905 0.25 2.035 ;
 RECT 3.18 1.125 3.31 1.255 ;
 RECT 3.5 0.755 3.63 0.885 ;
 RECT 2.56 1.52 2.69 1.65 ;
 RECT 0.255 1.255 0.385 1.385 ;
 RECT 3.5 2.145 3.63 2.275 ;
 RECT 3.5 1.885 3.63 2.015 ;
 RECT 0.75 2.2 0.88 2.33 ;
 RECT 3.5 1.625 3.63 1.755 ;
 RECT 3.915 0.395 4.045 0.525 ;
 RECT 3.915 1.695 4.045 1.825 ;
 RECT 3.03 2.145 3.16 2.275 ;
 RECT 1.67 2.22 1.8 2.35 ;
 RECT 3.03 2.405 3.16 2.535 ;
 RECT 2.56 0.755 2.69 0.885 ;
 RECT 2 0.555 2.13 0.685 ;
 RECT 3.915 2.215 4.045 2.345 ;
 RECT 1.53 0.54 1.66 0.67 ;
 RECT 1.06 0.55 1.19 0.68 ;
 RECT 2.725 0.385 2.855 0.515 ;
 RECT 3.915 1.955 4.045 2.085 ;
 RECT 0.12 0.55 0.25 0.68 ;
 LAYER M1 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.5 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 RECT 1.055 1.685 1.195 1.915 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 2.275 0.36 2.415 0.38 ;
 RECT 2.275 0.52 2.415 1.545 ;
 RECT 2.72 0.335 2.86 0.38 ;
 RECT 2.72 0.52 2.86 0.565 ;
 RECT 1.055 1.545 2.415 1.685 ;
 RECT 2.275 0.38 2.865 0.52 ;
 RECT 1.525 0.22 2.415 0.36 ;
 RECT 2.555 0.705 2.695 1.12 ;
 RECT 2.555 1.26 2.695 1.705 ;
 RECT 3.175 1.075 3.315 1.12 ;
 RECT 3.175 1.26 3.315 1.305 ;
 RECT 2.555 1.12 3.315 1.26 ;
 END
END OAI22X1

MACRO OAI22X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 2.88 ;
 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.715 1.46 2.07 1.72 ;
 END
 ANTENNAGATEAREA 0.073 ;
 END IN3

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 0.115 1.935 0.255 2.8 ;
 RECT 4.38 1.645 4.52 2.8 ;
 RECT 1.995 1.9 2.135 2.8 ;
 RECT 3.025 2.095 3.165 2.8 ;
 RECT 3.965 2.095 4.105 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 3.025 0.08 3.165 0.905 ;
 RECT 0.585 0.08 0.725 0.73 ;
 RECT 4.38 0.08 4.52 0.835 ;
 RECT 3.965 0.08 4.105 0.755 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.495 1.425 3.635 2.585 ;
 RECT 3.495 1.14 3.835 1.425 ;
 RECT 3.495 0.705 3.635 1.14 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END QN

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.29 2.34 1.645 2.58 ;
 END
 ANTENNAGATEAREA 0.073 ;
 END IN4

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.495 2.26 0.94 2.575 ;
 END
 ANTENNAGATEAREA 0.064 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.165 1.225 0.47 1.585 ;
 END
 ANTENNAGATEAREA 0.064 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 0.84 0.41 0.94 2.355 ;
 RECT 0.7 2.355 0.94 2.575 ;
 RECT 1.31 0.33 1.41 2.355 ;
 RECT 1.31 2.355 1.55 2.565 ;
 RECT 1.78 0.33 1.88 1.485 ;
 RECT 1.78 1.695 1.88 2.565 ;
 RECT 1.78 1.485 2.015 1.695 ;
 RECT 3.13 1.25 3.38 1.295 ;
 RECT 3.75 0.32 3.85 1.15 ;
 RECT 3.75 1.25 3.85 2.755 ;
 RECT 3.28 0.32 3.38 1.085 ;
 RECT 3.13 1.085 3.38 1.15 ;
 RECT 3.28 1.295 3.38 2.755 ;
 RECT 3.13 1.15 3.85 1.25 ;
 RECT 0.37 1.49 0.47 2.565 ;
 RECT 0.37 0.41 0.47 1.28 ;
 RECT 0.205 1.28 0.47 1.49 ;
 RECT 2.81 0.555 2.91 2.045 ;
 RECT 2.68 0.345 2.91 0.555 ;
 LAYER CO ;
 RECT 3.97 0.575 4.1 0.705 ;
 RECT 3.97 2.145 4.1 2.275 ;
 RECT 3.97 2.405 4.1 2.535 ;
 RECT 0.12 2.025 0.25 2.155 ;
 RECT 3.03 2.145 3.16 2.275 ;
 RECT 2 2.01 2.13 2.14 ;
 RECT 1.835 1.525 1.965 1.655 ;
 RECT 0.75 2.395 0.88 2.525 ;
 RECT 1.06 0.56 1.19 0.69 ;
 RECT 4.385 0.395 4.515 0.525 ;
 RECT 3.03 2.405 3.16 2.535 ;
 RECT 3.5 2.405 3.63 2.535 ;
 RECT 2.73 0.385 2.86 0.515 ;
 RECT 3.18 1.125 3.31 1.255 ;
 RECT 2.56 0.755 2.69 0.885 ;
 RECT 0.255 1.32 0.385 1.45 ;
 RECT 3.03 0.725 3.16 0.855 ;
 RECT 1.37 2.395 1.5 2.525 ;
 RECT 3.5 1.625 3.63 1.755 ;
 RECT 3.5 1.885 3.63 2.015 ;
 RECT 2 0.55 2.13 0.68 ;
 RECT 4.385 1.695 4.515 1.825 ;
 RECT 0.12 0.55 0.25 0.68 ;
 RECT 4.385 0.655 4.515 0.785 ;
 RECT 0.59 0.55 0.72 0.68 ;
 RECT 2.56 1.52 2.69 1.65 ;
 RECT 3.5 2.145 3.63 2.275 ;
 RECT 1.53 0.55 1.66 0.68 ;
 RECT 1.06 1.91 1.19 2.04 ;
 RECT 4.385 1.955 4.515 2.085 ;
 RECT 3.5 0.755 3.63 0.885 ;
 RECT 4.385 2.215 4.515 2.345 ;
 LAYER M1 ;
 RECT 0.115 0.5 0.255 0.87 ;
 RECT 1.055 0.505 1.195 0.87 ;
 RECT 1.995 0.5 2.135 0.87 ;
 RECT 0.115 0.87 2.135 1.01 ;
 RECT 1.055 1.29 1.195 2.115 ;
 RECT 1.525 0.36 1.665 0.73 ;
 RECT 2.725 0.335 2.865 0.38 ;
 RECT 2.725 0.52 2.865 0.565 ;
 RECT 2.275 0.52 2.415 1.15 ;
 RECT 2.275 0.36 2.415 0.38 ;
 RECT 1.055 1.15 2.415 1.29 ;
 RECT 2.275 0.38 2.865 0.52 ;
 RECT 1.525 0.22 2.415 0.36 ;
 RECT 2.555 0.705 2.695 1.12 ;
 RECT 2.555 1.26 2.695 1.705 ;
 RECT 3.175 1.075 3.315 1.12 ;
 RECT 3.175 1.26 3.315 1.305 ;
 RECT 2.555 1.12 3.315 1.26 ;
 END
END OAI22X2

MACRO SDFFARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 13.12 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 13.12 2.96 ;
 RECT 1.27 2.005 1.41 2.8 ;
 RECT 7.265 2.635 7.525 2.8 ;
 RECT 3.855 2.34 4.105 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 3.18 1.98 3.32 2.8 ;
 RECT 9.915 1.955 10.055 2.8 ;
 RECT 11.095 2.06 11.235 2.8 ;
 RECT 12.62 1.73 12.76 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 13.12 0.08 ;
 RECT 6.525 0.08 6.76 0.595 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 10.01 0.08 10.15 0.6 ;
 RECT 3.925 0.08 4.065 0.39 ;
 RECT 12.705 0.08 12.845 0.88 ;
 RECT 11.115 0.08 11.255 0.67 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.57 0.785 10.545 0.925 ;
 RECT 10.405 0.225 10.545 0.785 ;
 RECT 5.965 0.735 7.04 0.875 ;
 RECT 9.26 0.36 9.71 0.64 ;
 RECT 9.57 0.64 9.71 0.785 ;
 RECT 6.9 0.36 7.04 0.735 ;
 RECT 5.965 0.445 6.105 0.735 ;
 RECT 6.935 0.22 9.71 0.225 ;
 RECT 6.9 0.225 9.71 0.36 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 2.105 2.015 2.365 ;
 RECT 2.575 1.615 2.715 1.72 ;
 RECT 1.875 1.72 2.715 1.89 ;
 RECT 1.875 1.89 2.015 2.105 ;
 RECT 1.875 1.11 2.015 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.24 1.155 2.6 1.415 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.76 2.405 11.9 2.57 ;
 RECT 11.475 2.07 11.9 2.405 ;
 RECT 11.76 0.55 11.9 2.07 ;
 END
 ANTENNADIFFAREA 0.505 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.145 2.075 12.48 2.415 ;
 RECT 12.145 2.415 12.285 2.61 ;
 RECT 12.145 0.7 12.285 2.075 ;
 END
 ANTENNADIFFAREA 0.483 ;
 END Q

 OBS
 LAYER PO ;
 RECT 5.595 1.475 5.825 1.71 ;
 RECT 7.635 0.575 8.54 0.675 ;
 RECT 8.44 0.675 8.54 1.35 ;
 RECT 9.775 0.265 9.875 1.32 ;
 RECT 7.635 0.46 7.865 0.575 ;
 RECT 7.635 0.675 7.865 0.69 ;
 RECT 8.44 0.265 8.54 0.575 ;
 RECT 8.885 1.545 8.985 2.405 ;
 RECT 8.44 0.165 9.875 0.265 ;
 RECT 8.44 1.35 8.73 1.445 ;
 RECT 8.44 1.445 8.985 1.45 ;
 RECT 8.63 1.45 8.985 1.545 ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 2.665 1.865 2.765 2.48 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 4.28 1.265 4.38 1.52 ;
 RECT 3.78 1.52 4.38 1.62 ;
 RECT 4.215 1.62 4.315 2.68 ;
 RECT 6.895 1.79 6.995 2.68 ;
 RECT 3.78 1.44 4.025 1.52 ;
 RECT 3.78 1.62 4.025 1.69 ;
 RECT 5.145 0.705 5.245 1.165 ;
 RECT 4.28 0.585 4.38 1.165 ;
 RECT 5.145 0.47 5.43 0.705 ;
 RECT 4.215 2.68 6.995 2.78 ;
 RECT 4.28 1.165 5.245 1.265 ;
 RECT 2.245 1.41 2.345 1.645 ;
 RECT 2.665 0.655 2.765 1.18 ;
 RECT 2.195 1.745 2.295 2.47 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.245 1.18 2.765 1.41 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 4.6 0.285 4.7 0.51 ;
 RECT 4.6 0.185 6.435 0.285 ;
 RECT 6.335 0.285 6.435 1.24 ;
 RECT 4.56 0.51 4.805 0.755 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.245 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 5.1 1.595 5.2 2.48 ;
 RECT 4.56 1.445 4.805 1.495 ;
 RECT 4.56 1.495 5.2 1.595 ;
 RECT 4.56 1.595 4.805 1.69 ;
 RECT 9.7 1.575 9.8 2.585 ;
 RECT 8.48 2.47 8.7 2.585 ;
 RECT 8.48 2.685 8.7 2.71 ;
 RECT 8.48 2.585 9.8 2.685 ;
 RECT 8.91 0.685 9.01 1.255 ;
 RECT 8.835 0.455 9.065 0.685 ;
 RECT 7.95 1.64 8.39 1.865 ;
 RECT 8.155 1.865 8.39 1.87 ;
 RECT 7.95 1.105 8.175 1.64 ;
 RECT 7.86 0.875 8.175 1.105 ;
 RECT 11.18 1.05 11.645 1.28 ;
 RECT 11.545 0.135 11.645 1.05 ;
 RECT 11.545 1.28 11.645 2.79 ;
 RECT 12.405 0.32 12.505 1.19 ;
 RECT 12.405 1.425 12.505 2.79 ;
 RECT 12.39 1.19 12.6 1.425 ;
 RECT 10.79 1.32 10.89 2.7 ;
 RECT 10.49 0.47 10.59 1.22 ;
 RECT 10.49 1.22 10.89 1.32 ;
 RECT 10.36 0.23 10.59 0.47 ;
 RECT 6.035 0.695 6.135 1.61 ;
 RECT 6.07 1.71 6.17 2.48 ;
 RECT 6.035 1.61 6.17 1.71 ;
 RECT 5.915 0.465 6.155 0.695 ;
 RECT 9.38 0.645 9.48 1.18 ;
 RECT 9.38 1.39 9.48 2.295 ;
 RECT 9.36 1.18 9.595 1.39 ;
 RECT 10.19 0.65 10.29 1.71 ;
 RECT 10.19 1.71 10.435 1.95 ;
 RECT 10.19 1.95 10.29 2.7 ;
 RECT 7.2 1.61 7.465 1.82 ;
 RECT 7.365 1.82 7.465 2.49 ;
 RECT 6.995 0.635 7.095 1.51 ;
 RECT 6.995 1.51 7.465 1.61 ;
 RECT 5.595 1.33 5.735 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.635 0.65 5.735 1.33 ;
 LAYER CO ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 3.925 2.345 4.055 2.475 ;
 RECT 4.615 1.49 4.745 1.62 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 3.295 1.535 3.425 1.665 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 8.635 1.815 8.765 1.945 ;
 RECT 12.43 1.24 12.56 1.37 ;
 RECT 12.71 0.68 12.84 0.81 ;
 RECT 11.765 2.35 11.895 2.48 ;
 RECT 4.615 0.555 4.745 0.685 ;
 RECT 7.675 0.51 7.805 0.64 ;
 RECT 10.26 1.765 10.39 1.895 ;
 RECT 12.625 2.06 12.755 2.19 ;
 RECT 11.765 0.615 11.895 0.745 ;
 RECT 11.765 1.535 11.895 1.665 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 2.4 1.23 2.53 1.36 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 8.21 1.69 8.34 1.82 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 6.575 0.455 6.705 0.585 ;
 RECT 8.53 2.525 8.66 2.655 ;
 RECT 9.41 1.22 9.54 1.35 ;
 RECT 10.71 0.87 10.84 1 ;
 RECT 9.92 2.01 10.05 2.14 ;
 RECT 11.1 2.19 11.23 2.32 ;
 RECT 12.625 2.32 12.755 2.45 ;
 RECT 12.15 0.75 12.28 0.88 ;
 RECT 11.23 1.1 11.36 1.23 ;
 RECT 12.625 1.8 12.755 1.93 ;
 RECT 7.59 0.88 7.72 1.01 ;
 RECT 7.585 2.015 7.715 2.145 ;
 RECT 3.93 0.21 4.06 0.34 ;
 RECT 7.315 2.64 7.445 2.77 ;
 RECT 11.765 1.795 11.895 1.925 ;
 RECT 11.12 0.485 11.25 0.615 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 7.93 0.915 8.06 1.045 ;
 RECT 10.41 0.285 10.54 0.415 ;
 RECT 10.015 0.4 10.145 0.53 ;
 RECT 5.97 0.515 6.1 0.645 ;
 RECT 6.295 1.825 6.425 1.955 ;
 RECT 5.815 2.125 5.945 2.255 ;
 RECT 9.13 1.875 9.26 2.005 ;
 RECT 9.13 0.87 9.26 1 ;
 RECT 8.66 0.87 8.79 1 ;
 RECT 8.885 0.505 9.015 0.635 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 10.54 2.17 10.67 2.3 ;
 RECT 7.255 1.63 7.385 1.76 ;
 RECT 5.645 1.525 5.775 1.655 ;
 RECT 3.66 1.995 3.79 2.125 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 6.645 2.125 6.775 2.255 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 12.15 1.565 12.28 1.695 ;
 RECT 12.15 1.83 12.28 1.96 ;
 RECT 12.15 2.09 12.28 2.22 ;
 RECT 12.15 2.39 12.28 2.52 ;
 RECT 11.765 2.085 11.895 2.215 ;
 RECT 4.435 1.825 4.565 1.955 ;
 RECT 5.25 0.525 5.38 0.655 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 LAYER M1 ;
 RECT 10.705 0.815 11.535 0.955 ;
 RECT 11.395 0.36 11.535 0.815 ;
 RECT 9.405 1.17 9.545 1.395 ;
 RECT 9.405 1.395 10.845 1.535 ;
 RECT 10.705 0.955 10.845 1.395 ;
 RECT 10.535 1.535 10.675 2.36 ;
 RECT 11.395 0.22 12.565 0.36 ;
 RECT 12.425 0.36 12.565 1.45 ;
 RECT 5.745 2.12 6.845 2.26 ;
 RECT 5.18 0.52 5.825 0.66 ;
 RECT 5.685 0.66 5.825 1.015 ;
 RECT 7.18 0.505 7.855 0.645 ;
 RECT 5.685 1.015 7.32 1.155 ;
 RECT 7.18 0.645 7.32 1.015 ;
 RECT 7.58 1.015 8.13 1.05 ;
 RECT 7.58 1.05 7.72 1.3 ;
 RECT 7.58 1.44 7.72 2.215 ;
 RECT 6.305 1.3 7.72 1.44 ;
 RECT 7.52 0.91 8.13 1.015 ;
 RECT 7.52 0.875 7.79 0.91 ;
 RECT 5.575 1.52 6.445 1.66 ;
 RECT 6.305 1.44 6.445 1.52 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 9.125 1.815 9.335 1.87 ;
 RECT 9.125 0.805 9.265 1.675 ;
 RECT 9.055 1.87 9.335 2.01 ;
 RECT 10.815 1.92 10.955 2.505 ;
 RECT 9.125 1.675 10.395 1.815 ;
 RECT 10.255 2.505 10.955 2.645 ;
 RECT 10.255 1.815 10.395 2.505 ;
 RECT 11.05 1.235 11.19 1.78 ;
 RECT 11.05 1.095 11.43 1.235 ;
 RECT 10.815 1.78 11.19 1.92 ;
 RECT 8.14 1.685 8.795 1.81 ;
 RECT 8.655 1.005 8.795 1.685 ;
 RECT 8.14 1.81 8.835 1.825 ;
 RECT 8.565 1.825 8.835 1.95 ;
 RECT 8.585 0.865 8.865 1.005 ;
 RECT 3.7 1.63 3.84 1.99 ;
 RECT 3.7 1.475 4.045 1.63 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.59 1.99 3.84 2.13 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 5.36 0.805 5.5 1.22 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 5.185 1.36 5.325 1.82 ;
 RECT 5.185 1.82 7.39 1.96 ;
 RECT 7.25 1.58 7.39 1.82 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.365 2.11 2.995 2.195 ;
 RECT 2.365 2.195 2.99 2.25 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 4.89 0.36 5.03 2.035 ;
 RECT 3.46 0.53 4.345 0.67 ;
 RECT 4.205 0.22 5.03 0.36 ;
 RECT 4.205 0.36 4.345 0.53 ;
 RECT 4.845 2.035 5.03 2.17 ;
 RECT 4.845 2.17 4.985 2.305 ;
 RECT 4.495 0.5 4.75 0.965 ;
 RECT 4.495 1.96 4.635 2.51 ;
 RECT 4.495 1.67 4.635 1.82 ;
 RECT 4.495 0.965 4.635 1.44 ;
 RECT 4.495 1.44 4.75 1.67 ;
 RECT 4.365 1.82 4.635 1.96 ;
 RECT 4.495 2.51 7.125 2.65 ;
 RECT 6.985 2.495 7.125 2.51 ;
 RECT 6.985 2.355 8 2.495 ;
 RECT 8.46 2.24 8.6 2.52 ;
 RECT 7.86 2.24 8 2.355 ;
 RECT 7.86 1.35 8 2.1 ;
 RECT 7.86 2.1 8.6 2.24 ;
 RECT 7.86 1.21 8.44 1.35 ;
 RECT 8.46 2.52 8.73 2.66 ;
 RECT 8.58 0.5 9.09 0.58 ;
 RECT 8.3 0.58 9.09 0.64 ;
 RECT 8.3 0.64 8.76 0.72 ;
 RECT 8.3 0.72 8.44 1.21 ;
 END
END SDFFARX1

MACRO SDFFARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 13.76 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 13.76 2.96 ;
 RECT 7.265 2.635 7.525 2.8 ;
 RECT 3.855 2.34 4.105 2.8 ;
 RECT 1.27 2.005 1.41 2.8 ;
 RECT 3.18 1.98 3.32 2.8 ;
 RECT 9.915 1.955 10.055 2.8 ;
 RECT 11.095 2.06 11.235 2.8 ;
 RECT 13.235 1.73 13.375 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 12.23 1.465 12.37 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 13.76 0.08 ;
 RECT 6.525 0.08 6.76 0.595 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 13.515 0.08 13.655 0.88 ;
 RECT 11.115 0.08 11.255 0.67 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 12.365 0.08 12.505 0.3 ;
 RECT 3.925 0.08 4.065 0.39 ;
 RECT 10.015 0.08 10.155 0.58 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.57 0.785 10.545 0.925 ;
 RECT 10.405 0.225 10.545 0.785 ;
 RECT 5.965 0.735 7.04 0.875 ;
 RECT 9.275 0.36 9.71 0.645 ;
 RECT 9.57 0.645 9.71 0.785 ;
 RECT 6.9 0.36 7.04 0.735 ;
 RECT 5.965 0.445 6.105 0.735 ;
 RECT 6.935 0.22 9.71 0.225 ;
 RECT 6.9 0.225 9.71 0.36 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.6 2.07 2.015 2.41 ;
 RECT 2.575 1.615 2.715 1.72 ;
 RECT 1.875 1.72 2.715 1.89 ;
 RECT 1.875 1.89 2.015 2.07 ;
 RECT 1.875 1.11 2.015 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.255 1.155 2.6 1.415 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.68 2.24 11.995 2.57 ;
 RECT 11.76 0.72 11.9 2.24 ;
 END
 ANTENNADIFFAREA 0.616 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.635 2.09 12.96 2.4 ;
 RECT 12.7 2.4 12.84 2.61 ;
 RECT 12.7 0.98 13.085 1.12 ;
 RECT 12.7 1.12 12.84 2.09 ;
 RECT 12.945 0.72 13.085 0.98 ;
 END
 ANTENNADIFFAREA 0.666 ;
 END Q

 OBS
 LAYER PO ;
 RECT 6.895 1.79 6.995 2.68 ;
 RECT 5.145 0.47 5.43 0.705 ;
 RECT 5.145 0.705 5.245 1.165 ;
 RECT 3.78 1.44 4.025 1.52 ;
 RECT 3.78 1.62 4.025 1.69 ;
 RECT 4.28 0.585 4.38 1.165 ;
 RECT 4.215 2.68 6.995 2.78 ;
 RECT 4.28 1.165 5.245 1.265 ;
 RECT 5.1 1.595 5.2 2.48 ;
 RECT 4.56 1.445 4.805 1.495 ;
 RECT 4.56 1.495 5.2 1.595 ;
 RECT 4.56 1.595 4.805 1.69 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 2.245 1.41 2.345 1.645 ;
 RECT 2.665 0.655 2.765 1.18 ;
 RECT 2.195 1.745 2.295 2.47 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.245 1.18 2.765 1.41 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 11.18 1.05 11.645 1.135 ;
 RECT 11.18 1.135 12.115 1.235 ;
 RECT 11.545 0.2 11.645 1.05 ;
 RECT 11.545 1.28 11.645 2.79 ;
 RECT 11.18 1.235 11.645 1.28 ;
 RECT 12.015 0.2 12.115 1.135 ;
 RECT 12.015 1.235 12.115 2.79 ;
 RECT 13.19 1.19 13.4 1.265 ;
 RECT 13.3 0.38 13.4 1.19 ;
 RECT 13.02 1.365 13.4 1.425 ;
 RECT 13.02 1.425 13.12 2.79 ;
 RECT 12.73 0.38 12.83 1.265 ;
 RECT 12.485 1.265 13.4 1.365 ;
 RECT 12.485 1.365 12.585 2.79 ;
 RECT 9.38 0.645 9.48 1.18 ;
 RECT 9.38 1.39 9.48 2.295 ;
 RECT 9.36 1.18 9.595 1.39 ;
 RECT 8.91 0.685 9.01 1.255 ;
 RECT 8.835 0.455 9.065 0.685 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.245 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 6.335 0.285 6.435 1.24 ;
 RECT 4.6 0.185 6.435 0.285 ;
 RECT 4.6 0.285 4.7 0.51 ;
 RECT 4.56 0.51 4.805 0.755 ;
 RECT 10.19 0.65 10.29 1.71 ;
 RECT 10.19 1.71 10.435 1.95 ;
 RECT 10.19 1.95 10.29 2.7 ;
 RECT 9.7 1.575 9.8 2.585 ;
 RECT 8.48 2.47 8.7 2.585 ;
 RECT 8.48 2.685 8.7 2.71 ;
 RECT 8.48 2.585 9.8 2.685 ;
 RECT 7.635 0.575 8.54 0.675 ;
 RECT 8.44 0.675 8.54 1.35 ;
 RECT 9.775 0.265 9.875 1.32 ;
 RECT 7.635 0.46 7.865 0.575 ;
 RECT 7.635 0.675 7.865 0.69 ;
 RECT 8.44 0.265 8.54 0.575 ;
 RECT 8.885 1.545 8.985 2.405 ;
 RECT 8.44 0.165 9.875 0.265 ;
 RECT 8.44 1.35 8.73 1.445 ;
 RECT 8.44 1.445 8.985 1.45 ;
 RECT 8.63 1.45 8.985 1.545 ;
 RECT 7.2 1.61 7.465 1.82 ;
 RECT 7.365 1.82 7.465 2.49 ;
 RECT 6.995 0.635 7.095 1.51 ;
 RECT 6.995 1.51 7.465 1.61 ;
 RECT 5.595 1.33 5.735 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.635 0.65 5.735 1.33 ;
 RECT 5.595 1.475 5.825 1.71 ;
 RECT 7.955 1.64 8.39 1.87 ;
 RECT 7.955 1.105 8.175 1.64 ;
 RECT 7.86 0.875 8.175 1.105 ;
 RECT 10.79 1.32 10.89 2.7 ;
 RECT 10.49 0.47 10.59 1.22 ;
 RECT 10.49 1.22 10.89 1.32 ;
 RECT 10.36 0.23 10.59 0.47 ;
 RECT 6.035 0.695 6.135 1.61 ;
 RECT 6.07 1.71 6.17 2.48 ;
 RECT 6.035 1.61 6.17 1.71 ;
 RECT 5.915 0.465 6.155 0.695 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 2.665 1.865 2.765 2.48 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 4.28 1.265 4.38 1.52 ;
 RECT 3.78 1.52 4.38 1.62 ;
 RECT 4.215 1.62 4.315 2.68 ;
 LAYER CO ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 3.295 1.535 3.425 1.665 ;
 RECT 3.66 1.995 3.79 2.125 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 5.25 0.525 5.38 0.655 ;
 RECT 13.24 2.32 13.37 2.45 ;
 RECT 12.95 0.77 13.08 0.9 ;
 RECT 11.23 1.1 11.36 1.23 ;
 RECT 13.24 1.8 13.37 1.93 ;
 RECT 13.24 2.06 13.37 2.19 ;
 RECT 11.765 0.77 11.895 0.9 ;
 RECT 11.765 1.535 11.895 1.665 ;
 RECT 11.765 1.795 11.895 1.925 ;
 RECT 11.12 0.485 11.25 0.615 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 12.705 2.39 12.835 2.52 ;
 RECT 11.765 2.085 11.895 2.215 ;
 RECT 4.615 0.555 4.745 0.685 ;
 RECT 7.675 0.51 7.805 0.64 ;
 RECT 10.26 1.765 10.39 1.895 ;
 RECT 8.635 1.815 8.765 1.945 ;
 RECT 13.23 1.24 13.36 1.37 ;
 RECT 9.13 1.875 9.26 2.005 ;
 RECT 9.13 0.87 9.26 1 ;
 RECT 6.295 1.825 6.425 1.955 ;
 RECT 5.815 2.125 5.945 2.255 ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 3.925 2.345 4.055 2.475 ;
 RECT 10.54 2.17 10.67 2.3 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 8.53 2.525 8.66 2.655 ;
 RECT 5.97 0.515 6.1 0.645 ;
 RECT 6.575 0.455 6.705 0.585 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 7.255 1.63 7.385 1.76 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 8.21 1.69 8.34 1.82 ;
 RECT 7.93 0.915 8.06 1.045 ;
 RECT 10.41 0.285 10.54 0.415 ;
 RECT 12.37 0.12 12.5 0.25 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 10.02 0.4 10.15 0.53 ;
 RECT 12.235 1.535 12.365 1.665 ;
 RECT 12.235 2.085 12.365 2.215 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 5.645 1.525 5.775 1.655 ;
 RECT 7.59 0.88 7.72 1.01 ;
 RECT 7.585 2.015 7.715 2.145 ;
 RECT 3.93 0.21 4.06 0.34 ;
 RECT 7.315 2.64 7.445 2.77 ;
 RECT 6.645 2.125 6.775 2.255 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 2.4 1.23 2.53 1.36 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 12.705 1.565 12.835 1.695 ;
 RECT 12.705 1.83 12.835 1.96 ;
 RECT 12.705 2.09 12.835 2.22 ;
 RECT 4.435 1.825 4.565 1.955 ;
 RECT 13.52 0.68 13.65 0.81 ;
 RECT 11.765 2.35 11.895 2.48 ;
 RECT 8.66 0.87 8.79 1 ;
 RECT 8.885 0.505 9.015 0.635 ;
 RECT 9.41 1.22 9.54 1.35 ;
 RECT 10.71 0.87 10.84 1 ;
 RECT 9.92 2.01 10.05 2.14 ;
 RECT 11.1 2.19 11.23 2.32 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 12.235 1.795 12.365 1.925 ;
 RECT 12.235 2.35 12.365 2.48 ;
 RECT 4.615 1.49 4.745 1.62 ;
 LAYER M1 ;
 RECT 7.58 1.05 7.72 1.3 ;
 RECT 6.305 1.3 7.72 1.44 ;
 RECT 7.58 1.44 7.72 2.215 ;
 RECT 7.52 0.91 8.13 1.015 ;
 RECT 7.52 0.875 7.79 0.91 ;
 RECT 7.58 1.015 8.13 1.05 ;
 RECT 5.575 1.52 6.445 1.66 ;
 RECT 6.305 1.44 6.445 1.52 ;
 RECT 5.745 2.12 6.845 2.26 ;
 RECT 5.18 0.52 5.825 0.66 ;
 RECT 5.685 0.66 5.825 1.015 ;
 RECT 7.18 0.505 7.855 0.645 ;
 RECT 5.685 1.015 7.32 1.155 ;
 RECT 7.18 0.645 7.32 1.015 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.365 2.11 2.995 2.195 ;
 RECT 2.365 2.195 2.99 2.25 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 4.89 0.36 5.03 2.035 ;
 RECT 3.46 0.53 4.345 0.67 ;
 RECT 4.205 0.22 5.03 0.36 ;
 RECT 4.205 0.36 4.345 0.53 ;
 RECT 4.845 2.035 5.03 2.17 ;
 RECT 4.845 2.17 4.985 2.305 ;
 RECT 4.495 0.5 4.75 0.965 ;
 RECT 4.495 1.96 4.635 2.51 ;
 RECT 4.495 0.965 4.635 1.44 ;
 RECT 4.495 1.67 4.635 1.82 ;
 RECT 4.495 1.44 4.75 1.67 ;
 RECT 4.365 1.82 4.635 1.96 ;
 RECT 4.495 2.51 7.125 2.65 ;
 RECT 6.985 2.495 7.125 2.51 ;
 RECT 7.86 1.21 8.44 1.35 ;
 RECT 7.86 1.35 8 2.1 ;
 RECT 7.86 2.1 8.6 2.24 ;
 RECT 7.86 2.24 8 2.355 ;
 RECT 8.46 2.24 8.6 2.52 ;
 RECT 6.985 2.355 8 2.495 ;
 RECT 8.58 0.5 9.09 0.58 ;
 RECT 8.3 0.58 9.09 0.64 ;
 RECT 8.3 0.64 8.76 0.72 ;
 RECT 8.46 2.52 8.73 2.66 ;
 RECT 8.3 0.72 8.44 1.21 ;
 RECT 3.7 1.63 3.84 1.99 ;
 RECT 3.7 1.475 4.045 1.63 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.59 1.99 3.84 2.13 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 9.125 1.815 9.335 1.87 ;
 RECT 9.125 0.805 9.265 1.675 ;
 RECT 9.055 1.87 9.335 2.01 ;
 RECT 10.815 1.92 10.955 2.505 ;
 RECT 9.125 1.675 10.395 1.815 ;
 RECT 10.255 2.505 10.955 2.645 ;
 RECT 10.255 1.815 10.395 2.505 ;
 RECT 11.05 1.235 11.19 1.78 ;
 RECT 11.05 1.095 11.43 1.235 ;
 RECT 10.815 1.78 11.19 1.92 ;
 RECT 8.14 1.685 8.795 1.81 ;
 RECT 8.655 1.005 8.795 1.685 ;
 RECT 8.14 1.81 8.835 1.825 ;
 RECT 8.565 1.825 8.835 1.95 ;
 RECT 8.585 0.865 8.865 1.005 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 5.36 0.805 5.5 1.22 ;
 RECT 5.185 1.36 5.325 1.82 ;
 RECT 5.185 1.82 7.39 1.96 ;
 RECT 7.25 1.58 7.39 1.82 ;
 RECT 9.405 1.17 9.545 1.395 ;
 RECT 9.405 1.395 10.845 1.535 ;
 RECT 10.705 0.955 10.845 1.395 ;
 RECT 10.535 1.535 10.675 2.36 ;
 RECT 11.395 0.58 11.535 0.815 ;
 RECT 10.705 0.815 11.535 0.955 ;
 RECT 13.225 0.58 13.365 1.45 ;
 RECT 11.395 0.44 13.365 0.58 ;
 END
END SDFFARX2

MACRO SDFFASRSX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 14.72 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 14.72 2.96 ;
 RECT 7.265 2.635 7.525 2.8 ;
 RECT 11.075 2.21 11.215 2.8 ;
 RECT 12.195 2.06 12.335 2.8 ;
 RECT 13.72 1.485 13.86 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 3.18 1.93 3.32 2.8 ;
 RECT 4.025 1.93 4.165 2.8 ;
 RECT 8.285 2.38 8.425 2.8 ;
 RECT 1.27 2.005 1.41 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 14.72 0.08 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 3.88 0.08 4.11 0.39 ;
 RECT 10.545 0.08 10.8 1.005 ;
 RECT 13.645 0.08 13.93 0.275 ;
 RECT 6.525 0.08 6.76 0.37 ;
 RECT 12.215 0.08 12.355 0.565 ;
 RECT 0.3 0.08 0.44 0.81 ;
 RECT 1.27 0.08 1.41 1.055 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.195 0.97 10.335 1.16 ;
 RECT 5.92 0.51 7.075 0.65 ;
 RECT 10.195 1.16 11.485 1.3 ;
 RECT 6.935 0.36 7.075 0.51 ;
 RECT 9.41 0.36 9.76 0.65 ;
 RECT 9.62 0.97 9.76 0.975 ;
 RECT 9.62 0.83 10.335 0.97 ;
 RECT 9.62 0.65 9.76 0.83 ;
 RECT 6.935 0.22 9.715 0.225 ;
 RECT 6.935 0.225 9.76 0.36 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.575 2.04 2.015 2.415 ;
 RECT 2.575 1.86 2.715 1.89 ;
 RECT 1.875 1.72 2.715 1.86 ;
 RECT 2.575 1.615 2.715 1.72 ;
 RECT 1.875 1.86 2.015 2.04 ;
 RECT 1.875 1.11 2.015 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.2 1.155 2.715 1.43 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.92 0.32 10.255 0.67 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END SETB

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.09 1.11 14.415 1.475 ;
 RECT 14.19 1.475 14.33 2.585 ;
 RECT 14.19 0.705 14.33 1.11 ;
 END
 ANTENNADIFFAREA 0.462 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.78 1.44 12.92 2.575 ;
 RECT 12.78 1.12 13.105 1.44 ;
 RECT 12.78 0.5 12.92 1.12 ;
 END
 ANTENNADIFFAREA 0.64 ;
 END QN

 PIN S0
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.12 2.07 13.475 2.405 ;
 RECT 13.245 2.405 13.385 2.58 ;
 RECT 13.245 0.7 13.385 2.07 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END S0

 OBS
 LAYER PO ;
 RECT 8.62 0.265 8.72 0.535 ;
 RECT 7.635 0.46 7.865 0.535 ;
 RECT 7.635 0.535 8.72 0.635 ;
 RECT 7.635 0.635 7.865 0.69 ;
 RECT 9.065 1.545 9.165 2.175 ;
 RECT 8.62 0.165 10.475 0.265 ;
 RECT 8.62 1.35 8.91 1.445 ;
 RECT 8.62 1.445 9.165 1.45 ;
 RECT 8.81 1.45 9.165 1.545 ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 2.665 1.865 2.765 2.48 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 5.1 1.655 5.2 2.495 ;
 RECT 4.575 1.555 5.2 1.655 ;
 RECT 4.575 1.655 4.82 1.8 ;
 RECT 9.56 0.645 9.66 1.24 ;
 RECT 9.56 1.24 9.805 1.45 ;
 RECT 9.56 1.45 9.66 2.37 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 7.645 1.33 7.745 1.565 ;
 RECT 7.835 1.665 7.935 2.69 ;
 RECT 10.035 0.67 10.135 2.69 ;
 RECT 7.15 0.635 7.25 1.23 ;
 RECT 7.15 1.23 7.745 1.33 ;
 RECT 7.645 1.565 7.935 1.665 ;
 RECT 7.835 2.69 10.135 2.79 ;
 RECT 9.955 0.46 10.185 0.67 ;
 RECT 6.335 0.285 6.435 1.24 ;
 RECT 4.6 0.185 6.435 0.285 ;
 RECT 4.6 0.285 4.7 0.525 ;
 RECT 4.56 0.525 4.79 0.76 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.255 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 7.2 1.61 7.465 1.82 ;
 RECT 7.365 1.82 7.465 2.49 ;
 RECT 6.795 0.625 6.895 1.51 ;
 RECT 6.795 1.51 7.465 1.61 ;
 RECT 10.645 2.47 10.96 2.71 ;
 RECT 10.86 1.96 10.96 2.47 ;
 RECT 8.045 0.865 8.44 1.095 ;
 RECT 8.115 1.095 8.44 1.64 ;
 RECT 8.115 1.64 8.575 1.87 ;
 RECT 11.325 0.65 11.425 1.11 ;
 RECT 11.89 1.35 11.99 2.63 ;
 RECT 11.255 1.11 11.485 1.25 ;
 RECT 11.255 1.25 11.99 1.35 ;
 RECT 6.035 0.695 6.135 1.61 ;
 RECT 6.07 1.71 6.17 2.48 ;
 RECT 6.035 1.61 6.17 1.71 ;
 RECT 5.915 0.465 6.155 0.695 ;
 RECT 9.09 0.685 9.19 1.255 ;
 RECT 9.015 0.455 9.245 0.685 ;
 RECT 10.87 1.57 11.43 1.67 ;
 RECT 11.205 1.67 11.43 1.94 ;
 RECT 11.33 1.94 11.43 2.63 ;
 RECT 10.87 0.65 10.97 1.57 ;
 RECT 5.595 1.33 5.735 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.635 0.65 5.735 1.33 ;
 RECT 5.595 1.475 5.825 1.71 ;
 RECT 12.28 1.06 12.63 1.29 ;
 RECT 12.53 0.145 12.63 1.06 ;
 RECT 12.53 1.29 12.63 2.775 ;
 RECT 13.505 1.01 14.075 1.245 ;
 RECT 13.975 0.31 14.075 1.01 ;
 RECT 13.975 1.245 14.075 2.775 ;
 RECT 13.505 0.31 13.605 1.01 ;
 RECT 13.505 1.245 13.605 2.775 ;
 RECT 2.54 1.2 2.765 1.245 ;
 RECT 2.665 0.655 2.765 1.2 ;
 RECT 2.54 1.345 2.765 1.43 ;
 RECT 2.245 1.345 2.345 1.645 ;
 RECT 2.195 1.745 2.295 2.465 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.245 1.245 2.765 1.345 ;
 RECT 4.28 1.31 4.38 1.52 ;
 RECT 3.78 1.52 4.38 1.62 ;
 RECT 4.28 1.62 4.38 2.685 ;
 RECT 6.895 1.79 6.995 2.685 ;
 RECT 5.145 0.47 5.43 0.705 ;
 RECT 5.145 0.705 5.245 1.21 ;
 RECT 4.28 0.585 4.38 1.21 ;
 RECT 3.78 1.44 4.025 1.52 ;
 RECT 3.78 1.62 4.025 1.69 ;
 RECT 4.28 2.685 6.995 2.785 ;
 RECT 4.28 1.21 5.245 1.31 ;
 RECT 8.62 0.635 8.72 1.35 ;
 RECT 10.375 0.265 10.475 1.22 ;
 LAYER CO ;
 RECT 5.25 0.525 5.38 0.655 ;
 RECT 14.195 2.35 14.325 2.48 ;
 RECT 14.195 2.085 14.325 2.215 ;
 RECT 13.725 1.555 13.855 1.685 ;
 RECT 13.725 1.825 13.855 1.955 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 13.25 1.555 13.38 1.685 ;
 RECT 0.305 0.61 0.435 0.74 ;
 RECT 13.25 1.825 13.38 1.955 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 12.785 1.555 12.915 1.685 ;
 RECT 11.64 2.13 11.77 2.26 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 10.71 2.525 10.84 2.655 ;
 RECT 8.815 1.815 8.945 1.945 ;
 RECT 8.29 2.44 8.42 2.57 ;
 RECT 14.195 0.765 14.325 0.895 ;
 RECT 13.72 1.06 13.85 1.19 ;
 RECT 13.725 0.14 13.855 0.27 ;
 RECT 13.25 0.75 13.38 0.88 ;
 RECT 12.33 1.11 12.46 1.24 ;
 RECT 12.785 0.55 12.915 0.68 ;
 RECT 12.785 1.825 12.915 1.955 ;
 RECT 12.785 2.085 12.915 2.215 ;
 RECT 12.22 0.365 12.35 0.495 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 8.395 1.69 8.525 1.82 ;
 RECT 8.115 0.915 8.245 1.045 ;
 RECT 11.305 1.165 11.435 1.295 ;
 RECT 10.62 0.87 10.75 1 ;
 RECT 5.97 0.515 6.1 0.645 ;
 RECT 6.575 0.23 6.705 0.36 ;
 RECT 7.685 0.51 7.815 0.64 ;
 RECT 9.31 1.765 9.44 1.895 ;
 RECT 9.31 0.87 9.44 1 ;
 RECT 14.195 1.825 14.325 1.955 ;
 RECT 9.78 2.02 9.91 2.15 ;
 RECT 14.195 1.555 14.325 1.685 ;
 RECT 9.065 0.505 9.195 0.635 ;
 RECT 13.725 2.35 13.855 2.48 ;
 RECT 13.725 2.085 13.855 2.215 ;
 RECT 11.64 0.87 11.77 1 ;
 RECT 13.25 2.35 13.38 2.48 ;
 RECT 10.61 2.19 10.74 2.32 ;
 RECT 13.25 2.085 13.38 2.215 ;
 RECT 11.255 1.76 11.385 1.89 ;
 RECT 7.255 1.63 7.385 1.76 ;
 RECT 12.785 2.35 12.915 2.48 ;
 RECT 5.645 1.525 5.775 1.655 ;
 RECT 7.59 0.88 7.72 1.01 ;
 RECT 7.585 2.015 7.715 2.145 ;
 RECT 3.93 0.255 4.06 0.385 ;
 RECT 7.315 2.64 7.445 2.77 ;
 RECT 6.645 2.105 6.775 2.235 ;
 RECT 10.26 1.92 10.39 2.05 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 8.84 0.87 8.97 1 ;
 RECT 2.58 1.25 2.71 1.38 ;
 RECT 9.62 1.28 9.75 1.41 ;
 RECT 11.08 2.28 11.21 2.41 ;
 RECT 0.305 0.35 0.435 0.48 ;
 RECT 12.2 2.13 12.33 2.26 ;
 RECT 10.005 0.5 10.135 0.63 ;
 RECT 6.295 1.825 6.425 1.955 ;
 RECT 5.815 2.105 5.945 2.235 ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 4.03 2.005 4.16 2.135 ;
 RECT 4.61 0.58 4.74 0.71 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 4.63 1.6 4.76 1.73 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 3.305 1.535 3.435 1.665 ;
 RECT 3.66 1.995 3.79 2.125 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 1.995 3.315 2.125 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 4.5 2.015 4.63 2.145 ;
 LAYER M1 ;
 RECT 5.745 2.1 6.845 2.24 ;
 RECT 5.18 0.52 5.78 0.66 ;
 RECT 5.64 0.66 5.78 0.79 ;
 RECT 7.215 0.505 7.885 0.645 ;
 RECT 5.64 0.79 7.355 0.93 ;
 RECT 7.215 0.645 7.355 0.79 ;
 RECT 9.425 2.32 9.565 2.52 ;
 RECT 7.925 2.18 9.495 2.185 ;
 RECT 7.925 2.185 9.565 2.24 ;
 RECT 8.78 2.24 9.565 2.32 ;
 RECT 7.925 1.35 8.065 2.1 ;
 RECT 7.925 2.24 8.065 2.295 ;
 RECT 4.495 2.43 8.065 2.435 ;
 RECT 6.985 2.295 8.065 2.43 ;
 RECT 4.495 2.435 7.125 2.57 ;
 RECT 8.48 0.5 9.27 0.64 ;
 RECT 7.925 2.1 8.92 2.18 ;
 RECT 8.48 0.64 8.62 1.21 ;
 RECT 7.925 1.21 8.62 1.35 ;
 RECT 4.495 1.78 4.635 2.43 ;
 RECT 4.495 0.84 4.745 1.035 ;
 RECT 4.605 0.51 4.745 0.84 ;
 RECT 4.495 1.035 4.635 1.55 ;
 RECT 4.495 1.55 4.765 1.78 ;
 RECT 9.425 2.52 10.92 2.66 ;
 RECT 9.615 1.21 9.755 1.44 ;
 RECT 11.635 0.82 12.635 0.965 ;
 RECT 12.495 0.36 12.635 0.82 ;
 RECT 11.635 0.965 11.775 1.44 ;
 RECT 11.635 1.58 11.775 2.33 ;
 RECT 9.615 1.44 11.775 1.58 ;
 RECT 12.495 0.22 13.49 0.36 ;
 RECT 13.35 0.36 13.49 0.42 ;
 RECT 13.685 0.56 13.825 1.055 ;
 RECT 13.62 1.055 13.915 1.195 ;
 RECT 13.35 0.42 13.825 0.56 ;
 RECT 9.775 2.155 9.96 2.22 ;
 RECT 9.775 2.22 10.795 2.36 ;
 RECT 10.555 2.185 10.795 2.22 ;
 RECT 9.73 2.015 9.96 2.155 ;
 RECT 7.52 0.875 8.315 1.05 ;
 RECT 7.58 1.325 7.72 2.01 ;
 RECT 6.97 1.185 7.72 1.325 ;
 RECT 7.52 1.05 7.72 1.185 ;
 RECT 5.575 1.52 7.11 1.66 ;
 RECT 6.97 1.325 7.11 1.52 ;
 RECT 7.53 2.01 7.785 2.15 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 9.305 0.805 9.445 1.72 ;
 RECT 9.305 1.9 9.515 1.905 ;
 RECT 9.235 1.86 9.515 1.9 ;
 RECT 10.21 1.86 10.44 2.055 ;
 RECT 9.305 1.72 11.495 1.76 ;
 RECT 9.235 1.76 11.495 1.86 ;
 RECT 11.915 1.92 12.055 2.505 ;
 RECT 11.355 1.935 11.495 2.505 ;
 RECT 11.195 1.86 11.495 1.935 ;
 RECT 11.355 2.505 12.055 2.645 ;
 RECT 12.15 1.245 12.29 1.78 ;
 RECT 12.15 1.105 12.53 1.245 ;
 RECT 11.915 1.78 12.29 1.92 ;
 RECT 8.835 1.005 8.975 1.685 ;
 RECT 8.325 1.685 8.975 1.81 ;
 RECT 8.325 1.81 9.015 1.825 ;
 RECT 8.745 1.825 9.015 1.95 ;
 RECT 8.765 0.865 9.045 1.005 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.365 2.11 2.995 2.25 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 3.46 0.53 4.41 0.67 ;
 RECT 4.89 0.36 5.03 1.175 ;
 RECT 4.905 1.27 5.045 2.1 ;
 RECT 4.27 0.36 4.41 0.53 ;
 RECT 4.27 0.22 5.03 0.36 ;
 RECT 4.78 2.1 5.05 2.24 ;
 RECT 4.89 1.175 5.045 1.27 ;
 RECT 3.7 1.63 3.84 1.925 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.655 1.925 3.84 2.175 ;
 RECT 3.7 1.475 4.045 1.63 ;
 RECT 5.185 1.82 7.39 1.96 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 5.36 0.805 5.5 1.22 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 7.25 1.58 7.39 1.82 ;
 RECT 5.185 1.36 5.325 1.82 ;
 END
END SDFFASRSX1

MACRO SDFFASRSX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 15.68 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 15.68 2.96 ;
 RECT 7.265 2.635 7.525 2.8 ;
 RECT 12.195 2.06 12.335 2.8 ;
 RECT 14.195 1.485 14.335 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 3.18 1.93 3.32 2.8 ;
 RECT 4.025 1.93 4.165 2.8 ;
 RECT 13.25 1.505 13.39 2.8 ;
 RECT 15.135 1.485 15.275 2.8 ;
 RECT 8.285 2.38 8.425 2.8 ;
 RECT 1.27 2.005 1.41 2.8 ;
 RECT 11.075 2.145 11.215 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 15.68 0.08 ;
 RECT 13.175 0.08 13.46 0.255 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 6.525 0.08 6.76 0.37 ;
 RECT 14.12 0.08 14.405 0.275 ;
 RECT 3.88 0.08 4.11 0.39 ;
 RECT 10.545 0.08 10.8 1.005 ;
 RECT 12.03 0.08 12.17 0.625 ;
 RECT 0.3 0.08 0.44 0.81 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 15.135 0.08 15.275 0.945 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.935 0.22 9.9 0.36 ;
 RECT 8.025 0.36 8.33 0.46 ;
 RECT 5.92 0.51 7.075 0.65 ;
 RECT 9.76 0.83 10.335 0.97 ;
 RECT 10.195 0.97 10.335 1.16 ;
 RECT 10.195 1.16 11.485 1.3 ;
 RECT 6.935 0.36 7.075 0.51 ;
 RECT 9.76 0.36 9.9 0.83 ;
 END
 ANTENNAGATEAREA 0.11 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.615 2.04 2.015 2.415 ;
 RECT 2.575 1.86 2.715 1.89 ;
 RECT 1.875 1.72 2.715 1.86 ;
 RECT 2.575 1.615 2.715 1.72 ;
 RECT 1.875 1.86 2.015 2.04 ;
 RECT 1.875 1.11 2.015 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.2 1.165 2.715 1.43 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.625 2.42 9.285 2.66 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END SETB

 PIN S0
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.665 1.11 14.98 1.475 ;
 RECT 14.665 1.475 14.805 2.585 ;
 RECT 14.665 0.705 14.805 1.11 ;
 END
 ANTENNADIFFAREA 0.58 ;
 END S0

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.78 1.425 12.92 2.575 ;
 RECT 12.78 1.105 13.11 1.425 ;
 RECT 12.78 0.965 12.92 1.105 ;
 RECT 12.59 0.825 12.915 0.9 ;
 RECT 12.59 0.9 12.92 0.965 ;
 RECT 12.59 0.5 12.73 0.825 ;
 END
 ANTENNADIFFAREA 0.766 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.72 2.38 13.86 2.58 ;
 RECT 13.72 2.015 14.055 2.38 ;
 RECT 13.72 0.7 13.86 2.015 ;
 END
 ANTENNADIFFAREA 0.588 ;
 END Q

 OBS
 LAYER PO ;
 RECT 6.895 1.79 6.995 2.685 ;
 RECT 4.28 0.585 4.38 1.21 ;
 RECT 3.78 1.44 4.025 1.52 ;
 RECT 3.78 1.62 4.025 1.69 ;
 RECT 4.28 2.685 6.995 2.785 ;
 RECT 4.28 1.21 5.245 1.31 ;
 RECT 6.335 0.285 6.435 1.24 ;
 RECT 4.6 0.185 6.435 0.285 ;
 RECT 4.6 0.285 4.7 0.525 ;
 RECT 4.56 0.525 4.79 0.76 ;
 RECT 5.1 1.655 5.2 2.495 ;
 RECT 4.575 1.655 4.82 1.8 ;
 RECT 4.575 1.555 5.2 1.655 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.255 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 12.53 1.36 12.63 2.775 ;
 RECT 12.285 1.23 12.63 1.36 ;
 RECT 12.955 0.2 13.055 1.13 ;
 RECT 13.035 1.23 13.135 2.775 ;
 RECT 12.285 0.2 12.385 1.13 ;
 RECT 12.285 1.13 13.135 1.23 ;
 RECT 2.665 0.655 2.765 1.2 ;
 RECT 2.54 1.2 2.765 1.245 ;
 RECT 2.54 1.345 2.765 1.43 ;
 RECT 2.245 1.345 2.345 1.645 ;
 RECT 2.245 1.245 2.765 1.345 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.195 1.745 2.295 2.465 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 6.035 0.695 6.135 1.61 ;
 RECT 6.07 1.71 6.17 2.48 ;
 RECT 6.035 1.61 6.17 1.71 ;
 RECT 5.915 0.465 6.155 0.695 ;
 RECT 9.56 0.645 9.66 1.24 ;
 RECT 9.56 1.24 9.805 1.45 ;
 RECT 9.56 1.45 9.66 2.37 ;
 RECT 9.09 0.685 9.19 1.255 ;
 RECT 9.015 0.455 9.245 0.685 ;
 RECT 8.62 0.635 8.72 1.35 ;
 RECT 10.375 0.265 10.475 1.22 ;
 RECT 8.62 0.265 8.72 0.535 ;
 RECT 7.635 0.46 7.865 0.535 ;
 RECT 7.635 0.535 8.72 0.635 ;
 RECT 7.635 0.635 7.865 0.69 ;
 RECT 9.065 1.545 9.165 2.205 ;
 RECT 8.62 0.165 10.475 0.265 ;
 RECT 8.62 1.35 8.91 1.445 ;
 RECT 8.62 1.445 9.165 1.45 ;
 RECT 8.81 1.45 9.165 1.545 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 11.255 1.25 11.99 1.35 ;
 RECT 11.89 1.35 11.99 2.63 ;
 RECT 11.255 1.11 11.485 1.25 ;
 RECT 11.325 0.65 11.425 1.11 ;
 RECT 5.595 1.33 5.735 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.635 0.65 5.735 1.33 ;
 RECT 5.595 1.475 5.825 1.71 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 7.67 1.33 7.77 1.565 ;
 RECT 7.875 1.665 7.975 2.69 ;
 RECT 10.035 0.635 10.135 2.69 ;
 RECT 8.625 2.435 8.855 2.69 ;
 RECT 7.15 0.635 7.25 1.23 ;
 RECT 7.15 1.23 7.77 1.33 ;
 RECT 7.67 1.565 7.975 1.665 ;
 RECT 7.875 2.69 10.135 2.79 ;
 RECT 7.2 1.61 7.465 1.82 ;
 RECT 7.365 1.82 7.465 2.49 ;
 RECT 6.795 0.625 6.895 1.51 ;
 RECT 6.795 1.51 7.465 1.61 ;
 RECT 10.645 2.47 10.96 2.71 ;
 RECT 10.86 1.96 10.96 2.47 ;
 RECT 14.45 0.31 14.55 1.01 ;
 RECT 13.98 1.01 14.55 1.13 ;
 RECT 14.45 1.245 14.55 2.775 ;
 RECT 13.98 1.23 14.55 1.245 ;
 RECT 13.98 0.31 14.08 1.01 ;
 RECT 13.98 1.245 14.08 2.775 ;
 RECT 13.505 1.13 15.02 1.23 ;
 RECT 14.92 0.31 15.02 1.13 ;
 RECT 14.92 1.23 15.02 2.775 ;
 RECT 13.505 0.31 13.605 1.13 ;
 RECT 13.505 1.23 13.605 2.775 ;
 RECT 8.155 1.64 8.575 1.87 ;
 RECT 8.155 1.095 8.36 1.64 ;
 RECT 8.045 0.865 8.36 1.095 ;
 RECT 10.87 1.57 11.43 1.67 ;
 RECT 11.205 1.67 11.43 1.94 ;
 RECT 10.87 0.65 10.97 1.57 ;
 RECT 11.33 1.94 11.43 2.63 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 2.665 1.865 2.765 2.48 ;
 RECT 4.28 1.31 4.38 1.52 ;
 RECT 3.78 1.52 4.38 1.62 ;
 RECT 4.28 1.62 4.38 2.685 ;
 RECT 5.145 0.47 5.43 0.705 ;
 RECT 5.145 0.705 5.245 1.21 ;
 LAYER CO ;
 RECT 11.255 1.76 11.385 1.89 ;
 RECT 10.71 2.525 10.84 2.655 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 14.195 1.06 14.325 1.19 ;
 RECT 14.2 0.14 14.33 0.27 ;
 RECT 13.725 0.75 13.855 0.88 ;
 RECT 13.255 2.35 13.385 2.48 ;
 RECT 13.255 1.825 13.385 1.955 ;
 RECT 12.595 0.55 12.725 0.68 ;
 RECT 12.785 1.825 12.915 1.955 ;
 RECT 12.785 2.085 12.915 2.215 ;
 RECT 12.035 0.445 12.165 0.575 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 5.25 0.525 5.38 0.655 ;
 RECT 14.67 2.35 14.8 2.48 ;
 RECT 14.67 1.825 14.8 1.955 ;
 RECT 14.67 2.085 14.8 2.215 ;
 RECT 14.67 1.555 14.8 1.685 ;
 RECT 14.2 1.555 14.33 1.685 ;
 RECT 14.2 2.35 14.33 2.48 ;
 RECT 9.31 1.765 9.44 1.895 ;
 RECT 9.31 0.87 9.44 1 ;
 RECT 10.26 1.92 10.39 2.05 ;
 RECT 9.78 2.02 9.91 2.15 ;
 RECT 8.84 0.87 8.97 1 ;
 RECT 9.065 0.505 9.195 0.635 ;
 RECT 13.725 2.085 13.855 2.215 ;
 RECT 5.815 2.105 5.945 2.235 ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 4.03 2.005 4.16 2.135 ;
 RECT 4.61 0.58 4.74 0.71 ;
 RECT 8.29 2.44 8.42 2.57 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 7.315 2.64 7.445 2.77 ;
 RECT 6.645 2.105 6.775 2.235 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 4.63 1.6 4.76 1.73 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 3.305 1.535 3.435 1.665 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 8.815 1.815 8.945 1.945 ;
 RECT 13.255 0.12 13.385 0.25 ;
 RECT 15.14 0.74 15.27 0.87 ;
 RECT 15.14 1.555 15.27 1.685 ;
 RECT 15.14 2.35 15.27 2.48 ;
 RECT 15.14 1.825 15.27 1.955 ;
 RECT 15.14 2.085 15.27 2.215 ;
 RECT 13.255 1.555 13.385 1.685 ;
 RECT 12.335 1.18 12.465 1.31 ;
 RECT 13.255 2.085 13.385 2.215 ;
 RECT 8.115 0.915 8.245 1.045 ;
 RECT 11.305 1.165 11.435 1.295 ;
 RECT 10.62 0.87 10.75 1 ;
 RECT 5.97 0.515 6.1 0.645 ;
 RECT 6.575 0.23 6.705 0.36 ;
 RECT 7.685 0.51 7.815 0.64 ;
 RECT 0.305 0.61 0.435 0.74 ;
 RECT 0.305 0.35 0.435 0.48 ;
 RECT 9.62 1.28 9.75 1.41 ;
 RECT 11.64 0.87 11.77 1 ;
 RECT 11.08 2.215 11.21 2.345 ;
 RECT 10.61 2.19 10.74 2.32 ;
 RECT 12.2 2.13 12.33 2.26 ;
 RECT 6.295 1.825 6.425 1.955 ;
 RECT 7.255 1.63 7.385 1.76 ;
 RECT 5.645 1.525 5.775 1.655 ;
 RECT 7.59 0.88 7.72 1.01 ;
 RECT 7.585 2.015 7.715 2.145 ;
 RECT 3.93 0.255 4.06 0.385 ;
 RECT 14.2 1.825 14.33 1.955 ;
 RECT 14.67 0.765 14.8 0.895 ;
 RECT 3.185 1.995 3.315 2.125 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 8.395 1.69 8.525 1.82 ;
 RECT 4.5 2.015 4.63 2.145 ;
 RECT 12.785 2.35 12.915 2.48 ;
 RECT 12.785 1.555 12.915 1.685 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 2.58 1.25 2.71 1.38 ;
 RECT 14.2 2.085 14.33 2.215 ;
 RECT 13.725 1.555 13.855 1.685 ;
 RECT 13.725 2.35 13.855 2.48 ;
 RECT 13.725 1.825 13.855 1.955 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 8.685 2.485 8.815 2.615 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.66 1.995 3.79 2.125 ;
 RECT 11.64 2.13 11.77 2.26 ;
 LAYER M1 ;
 RECT 5.745 2.1 6.845 2.24 ;
 RECT 5.18 0.52 5.78 0.66 ;
 RECT 5.64 0.66 5.78 0.79 ;
 RECT 7.215 0.505 7.865 0.645 ;
 RECT 5.64 0.79 7.355 0.93 ;
 RECT 7.215 0.645 7.355 0.79 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.365 2.11 2.995 2.25 ;
 RECT 3.46 0.53 4.41 0.67 ;
 RECT 4.89 0.36 5.03 1.175 ;
 RECT 4.905 1.27 5.045 2.1 ;
 RECT 4.27 0.36 4.41 0.53 ;
 RECT 4.27 0.22 5.03 0.36 ;
 RECT 4.78 2.1 5.05 2.24 ;
 RECT 4.89 1.175 5.045 1.27 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 12.875 0.555 13.57 0.65 ;
 RECT 12.31 0.36 12.45 0.82 ;
 RECT 11.635 0.82 12.45 0.965 ;
 RECT 12.875 0.36 13.015 0.51 ;
 RECT 12.31 0.22 13.015 0.36 ;
 RECT 11.635 0.965 11.775 1.44 ;
 RECT 11.635 1.58 11.775 2.33 ;
 RECT 9.615 1.44 11.775 1.58 ;
 RECT 9.615 1.21 9.755 1.44 ;
 RECT 14.17 0.555 14.31 1.055 ;
 RECT 14.095 1.055 14.39 1.195 ;
 RECT 13.43 0.415 14.31 0.51 ;
 RECT 12.875 0.51 14.31 0.555 ;
 RECT 9.775 2.155 9.96 2.22 ;
 RECT 9.775 2 9.915 2.015 ;
 RECT 9.775 2.22 10.795 2.36 ;
 RECT 10.555 2.185 10.795 2.22 ;
 RECT 9.73 2.015 9.96 2.155 ;
 RECT 8.835 1.005 8.975 1.685 ;
 RECT 8.325 1.685 8.975 1.81 ;
 RECT 8.325 1.81 9.015 1.825 ;
 RECT 8.745 1.825 9.015 1.95 ;
 RECT 8.765 0.865 9.045 1.005 ;
 RECT 5.185 1.82 7.39 1.96 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 5.36 0.805 5.5 1.22 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 7.25 1.575 7.39 1.82 ;
 RECT 5.185 1.36 5.325 1.82 ;
 RECT 7.52 0.875 8.315 1.05 ;
 RECT 7.58 1.325 7.72 2.01 ;
 RECT 6.97 1.185 7.72 1.325 ;
 RECT 7.52 1.05 7.72 1.185 ;
 RECT 5.575 1.52 7.11 1.66 ;
 RECT 6.97 1.325 7.11 1.52 ;
 RECT 7.53 2.01 7.785 2.15 ;
 RECT 9.305 1.72 11.495 1.76 ;
 RECT 9.235 1.76 11.495 1.86 ;
 RECT 11.915 1.92 12.055 2.505 ;
 RECT 11.355 1.935 11.495 2.505 ;
 RECT 11.195 1.86 11.495 1.935 ;
 RECT 11.355 2.505 12.055 2.645 ;
 RECT 9.305 1.9 9.515 1.905 ;
 RECT 9.305 0.805 9.445 1.72 ;
 RECT 9.235 1.86 9.515 1.9 ;
 RECT 10.21 1.86 10.44 2.055 ;
 RECT 12.15 1.315 12.29 1.78 ;
 RECT 12.15 1.175 12.54 1.315 ;
 RECT 11.915 1.78 12.29 1.92 ;
 RECT 7.925 1.35 8.065 2.1 ;
 RECT 7.925 2.24 8.065 2.295 ;
 RECT 4.495 2.43 8.065 2.435 ;
 RECT 6.985 2.295 8.065 2.43 ;
 RECT 4.495 2.435 7.125 2.57 ;
 RECT 4.495 1.78 4.635 2.43 ;
 RECT 4.495 0.84 4.745 1.035 ;
 RECT 4.605 0.51 4.745 0.84 ;
 RECT 4.495 1.035 4.635 1.55 ;
 RECT 4.495 1.55 4.765 1.78 ;
 RECT 8.48 0.64 8.62 1.21 ;
 RECT 7.925 1.21 8.62 1.35 ;
 RECT 9.425 2.24 9.565 2.52 ;
 RECT 8.48 0.5 9.27 0.64 ;
 RECT 7.925 2.1 9.565 2.24 ;
 RECT 9.425 2.52 10.92 2.66 ;
 RECT 3.7 1.63 3.84 1.925 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.655 1.925 3.84 2.175 ;
 RECT 3.7 1.475 4.045 1.63 ;
 END
END SDFFASRSX2

MACRO SDFFASRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 14.08 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 14.08 2.96 ;
 RECT 7.265 2.635 7.525 2.8 ;
 RECT 11.075 2.21 11.215 2.8 ;
 RECT 12.195 2.06 12.335 2.8 ;
 RECT 13.72 1.485 13.86 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 3.18 1.93 3.32 2.8 ;
 RECT 4.025 1.93 4.165 2.8 ;
 RECT 1.27 1.985 1.41 2.8 ;
 RECT 8.285 2.38 8.425 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 14.08 0.08 ;
 RECT 6.525 0.08 6.76 0.37 ;
 RECT 3.88 0.08 4.11 0.39 ;
 RECT 10.545 0.08 10.8 1.005 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 12.215 0.08 12.355 0.565 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 13.835 0.08 13.975 0.86 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.92 0.51 7.075 0.65 ;
 RECT 10.195 1.16 11.485 1.3 ;
 RECT 6.935 0.22 9.815 0.36 ;
 RECT 9.44 0.36 9.815 0.65 ;
 RECT 10.195 1.06 10.335 1.16 ;
 RECT 9.675 0.65 9.815 0.92 ;
 RECT 9.675 0.92 10.335 1.06 ;
 RECT 6.935 0.36 7.075 0.51 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.615 2.04 2.015 2.415 ;
 RECT 2.575 1.86 2.715 1.89 ;
 RECT 1.875 1.72 2.715 1.86 ;
 RECT 2.575 1.615 2.715 1.72 ;
 RECT 1.875 1.86 2.015 2.04 ;
 RECT 1.875 1.11 2.015 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.2 1.155 2.715 1.43 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.955 0.445 10.23 0.76 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.78 1.445 12.92 2.575 ;
 RECT 12.78 1.105 13.09 1.445 ;
 RECT 12.78 0.5 12.92 1.105 ;
 END
 ANTENNADIFFAREA 0.64 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.12 2.075 13.455 2.4 ;
 RECT 13.245 2.4 13.385 2.58 ;
 RECT 13.145 0.7 13.285 0.745 ;
 RECT 13.245 0.93 13.385 2.075 ;
 RECT 13.145 0.745 13.385 0.93 ;
 END
 ANTENNADIFFAREA 0.469 ;
 END Q

 OBS
 LAYER PO ;
 RECT 2.54 1.2 2.765 1.245 ;
 RECT 2.54 1.345 2.765 1.43 ;
 RECT 2.245 1.345 2.345 1.645 ;
 RECT 2.195 1.745 2.295 2.465 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.245 1.245 2.765 1.345 ;
 RECT 11.255 1.25 11.99 1.35 ;
 RECT 11.89 1.35 11.99 2.63 ;
 RECT 11.255 1.11 11.485 1.25 ;
 RECT 11.325 0.65 11.425 1.11 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 4.28 1.62 4.38 2.685 ;
 RECT 4.28 1.31 4.38 1.52 ;
 RECT 3.78 1.52 4.38 1.62 ;
 RECT 6.895 1.79 6.995 2.685 ;
 RECT 4.28 2.685 6.995 2.775 ;
 RECT 4.28 2.775 6.945 2.785 ;
 RECT 3.78 1.44 4.025 1.52 ;
 RECT 3.78 1.62 4.025 1.69 ;
 RECT 5.145 0.705 5.245 1.21 ;
 RECT 4.28 0.585 4.38 1.21 ;
 RECT 5.145 0.47 5.43 0.705 ;
 RECT 4.28 1.21 5.245 1.31 ;
 RECT 7.67 1.33 7.77 1.565 ;
 RECT 7.86 1.665 7.96 2.69 ;
 RECT 10.035 0.73 10.135 2.69 ;
 RECT 7.15 0.635 7.25 1.23 ;
 RECT 7.15 1.23 7.77 1.33 ;
 RECT 7.67 1.565 7.96 1.665 ;
 RECT 7.86 2.69 10.135 2.79 ;
 RECT 9.965 0.52 10.195 0.73 ;
 RECT 6.335 0.285 6.435 1.24 ;
 RECT 4.6 0.185 6.435 0.285 ;
 RECT 4.6 0.285 4.7 0.525 ;
 RECT 4.56 0.525 4.79 0.76 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 10.645 2.47 10.96 2.71 ;
 RECT 10.86 1.96 10.96 2.47 ;
 RECT 12.53 0.145 12.63 1.06 ;
 RECT 12.53 1.29 12.63 2.775 ;
 RECT 12.28 1.06 12.63 1.29 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 2.665 1.865 2.765 2.48 ;
 RECT 6.035 0.695 6.135 1.61 ;
 RECT 6.07 1.71 6.17 2.48 ;
 RECT 6.035 1.61 6.17 1.71 ;
 RECT 5.915 0.465 6.155 0.695 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 8.045 0.865 8.36 1.095 ;
 RECT 8.14 1.095 8.36 1.64 ;
 RECT 8.14 1.64 8.575 1.87 ;
 RECT 9.56 0.645 9.66 1.24 ;
 RECT 9.56 1.24 9.805 1.45 ;
 RECT 9.56 1.45 9.66 2.37 ;
 RECT 9.09 0.685 9.19 1.255 ;
 RECT 9.015 0.455 9.245 0.685 ;
 RECT 7.2 1.61 7.465 1.82 ;
 RECT 7.365 1.82 7.465 2.49 ;
 RECT 6.795 0.625 6.895 1.51 ;
 RECT 6.795 1.51 7.465 1.61 ;
 RECT 5.595 1.33 5.735 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.635 0.65 5.735 1.33 ;
 RECT 5.595 1.475 5.825 1.71 ;
 RECT 11.205 1.67 11.43 1.94 ;
 RECT 11.33 1.94 11.43 2.63 ;
 RECT 10.87 0.65 10.97 1.57 ;
 RECT 10.87 1.57 11.43 1.67 ;
 RECT 13.4 0.35 13.5 1.01 ;
 RECT 13.505 1.245 13.605 2.775 ;
 RECT 13.4 1.01 13.815 1.245 ;
 RECT 5.1 1.655 5.2 2.495 ;
 RECT 4.575 1.655 4.82 1.8 ;
 RECT 4.575 1.555 5.2 1.655 ;
 RECT 8.62 0.635 8.72 1.35 ;
 RECT 9.065 1.545 9.165 2.175 ;
 RECT 10.375 0.265 10.475 1.22 ;
 RECT 8.62 0.265 8.72 0.535 ;
 RECT 7.635 0.46 7.865 0.535 ;
 RECT 7.635 0.535 8.72 0.635 ;
 RECT 7.635 0.635 7.865 0.69 ;
 RECT 8.62 0.165 10.475 0.265 ;
 RECT 8.81 1.45 9.165 1.545 ;
 RECT 8.62 1.35 8.91 1.445 ;
 RECT 8.62 1.445 9.165 1.45 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.255 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 2.665 0.655 2.765 1.2 ;
 LAYER CO ;
 RECT 13.635 1.06 13.765 1.19 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 12.785 2.085 12.915 2.215 ;
 RECT 12.22 0.365 12.35 0.495 ;
 RECT 8.115 0.915 8.245 1.045 ;
 RECT 11.305 1.165 11.435 1.295 ;
 RECT 10.62 0.87 10.75 1 ;
 RECT 5.97 0.515 6.1 0.645 ;
 RECT 8.395 1.69 8.525 1.82 ;
 RECT 9.31 1.765 9.44 1.895 ;
 RECT 9.31 0.87 9.44 1 ;
 RECT 10.26 1.92 10.39 2.05 ;
 RECT 9.78 2.02 9.91 2.15 ;
 RECT 8.84 0.87 8.97 1 ;
 RECT 9.065 0.505 9.195 0.635 ;
 RECT 6.575 0.23 6.705 0.36 ;
 RECT 7.685 0.51 7.815 0.64 ;
 RECT 13.725 1.555 13.855 1.685 ;
 RECT 13.725 2.35 13.855 2.48 ;
 RECT 13.725 1.825 13.855 1.955 ;
 RECT 13.725 2.085 13.855 2.215 ;
 RECT 13.25 1.555 13.38 1.685 ;
 RECT 13.25 2.35 13.38 2.48 ;
 RECT 9.62 1.28 9.75 1.41 ;
 RECT 11.64 0.87 11.77 1 ;
 RECT 11.08 2.28 11.21 2.41 ;
 RECT 10.61 2.19 10.74 2.32 ;
 RECT 12.2 2.13 12.33 2.26 ;
 RECT 11.64 2.13 11.77 2.26 ;
 RECT 11.255 1.76 11.385 1.89 ;
 RECT 13.25 1.825 13.38 1.955 ;
 RECT 13.25 2.085 13.38 2.215 ;
 RECT 12.785 1.555 12.915 1.685 ;
 RECT 12.785 2.35 12.915 2.48 ;
 RECT 7.255 1.63 7.385 1.76 ;
 RECT 5.645 1.525 5.775 1.655 ;
 RECT 7.59 0.88 7.72 1.01 ;
 RECT 7.585 2.015 7.715 2.145 ;
 RECT 3.93 0.255 4.06 0.385 ;
 RECT 7.315 2.64 7.445 2.77 ;
 RECT 6.295 1.825 6.425 1.955 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 4.63 1.6 4.76 1.73 ;
 RECT 3.305 1.535 3.435 1.665 ;
 RECT 3.66 1.995 3.79 2.125 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 1.995 3.315 2.125 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 4.5 2.015 4.63 2.145 ;
 RECT 5.25 0.525 5.38 0.655 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 10.71 2.525 10.84 2.655 ;
 RECT 10.015 0.56 10.145 0.69 ;
 RECT 5.815 2.105 5.945 2.235 ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 4.03 2.005 4.16 2.135 ;
 RECT 4.61 0.58 4.74 0.71 ;
 RECT 6.645 2.105 6.775 2.235 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 2.58 1.25 2.71 1.38 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 13.15 0.75 13.28 0.88 ;
 RECT 12.33 1.11 12.46 1.24 ;
 RECT 12.785 0.55 12.915 0.68 ;
 RECT 12.785 1.825 12.915 1.955 ;
 RECT 8.815 1.77 8.945 1.9 ;
 RECT 8.29 2.44 8.42 2.57 ;
 RECT 13.84 0.68 13.97 0.81 ;
 LAYER M1 ;
 RECT 5.745 2.1 6.845 2.24 ;
 RECT 5.18 0.52 5.78 0.66 ;
 RECT 5.64 0.66 5.78 0.79 ;
 RECT 7.215 0.505 7.88 0.645 ;
 RECT 5.64 0.79 7.355 0.93 ;
 RECT 7.215 0.645 7.355 0.79 ;
 RECT 7.925 2.185 9.565 2.24 ;
 RECT 7.925 2.1 9.56 2.185 ;
 RECT 9.425 2.24 9.565 2.52 ;
 RECT 7.925 1.35 8.065 2.1 ;
 RECT 7.925 2.24 8.065 2.295 ;
 RECT 4.495 2.43 8.065 2.435 ;
 RECT 6.985 2.295 8.065 2.43 ;
 RECT 4.495 2.435 7.125 2.57 ;
 RECT 8.48 0.5 9.27 0.64 ;
 RECT 8.48 0.64 8.62 1.21 ;
 RECT 7.925 1.21 8.62 1.35 ;
 RECT 4.495 1.78 4.635 2.43 ;
 RECT 4.495 0.84 4.745 1.035 ;
 RECT 4.605 0.51 4.745 0.84 ;
 RECT 4.495 1.035 4.635 1.55 ;
 RECT 4.495 1.55 4.765 1.78 ;
 RECT 9.425 2.52 10.92 2.66 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.365 2.11 2.995 2.25 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 3.46 0.53 4.41 0.67 ;
 RECT 4.89 0.36 5.03 1.175 ;
 RECT 4.905 1.27 5.045 2.1 ;
 RECT 4.27 0.36 4.41 0.53 ;
 RECT 4.27 0.22 5.03 0.36 ;
 RECT 4.78 2.1 5.05 2.24 ;
 RECT 4.89 1.175 5.045 1.27 ;
 RECT 9.775 2.155 9.96 2.22 ;
 RECT 9.775 2 9.915 2.015 ;
 RECT 9.775 2.22 10.795 2.36 ;
 RECT 10.555 2.185 10.795 2.22 ;
 RECT 9.73 2.015 9.96 2.155 ;
 RECT 8.325 1.685 8.975 1.765 ;
 RECT 8.835 1.005 8.975 1.685 ;
 RECT 8.325 1.765 9.015 1.825 ;
 RECT 8.745 1.825 9.015 1.905 ;
 RECT 8.765 0.865 9.045 1.005 ;
 RECT 3.7 1.63 3.84 1.925 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.655 1.925 3.84 2.175 ;
 RECT 3.7 1.475 4.045 1.63 ;
 RECT 7.52 0.875 8.315 1.05 ;
 RECT 6.97 1.185 7.72 1.325 ;
 RECT 7.58 1.325 7.72 2.01 ;
 RECT 7.52 1.05 7.72 1.185 ;
 RECT 5.575 1.52 7.11 1.66 ;
 RECT 6.97 1.325 7.11 1.52 ;
 RECT 7.53 2.01 7.785 2.15 ;
 RECT 9.615 1.21 9.755 1.44 ;
 RECT 11.635 0.82 12.635 0.965 ;
 RECT 12.495 0.36 12.635 0.82 ;
 RECT 11.635 0.965 11.775 1.44 ;
 RECT 11.635 1.58 11.775 2.33 ;
 RECT 9.615 1.44 11.775 1.58 ;
 RECT 13.53 0.56 13.67 1.055 ;
 RECT 12.495 0.22 13.335 0.36 ;
 RECT 13.195 0.42 13.67 0.56 ;
 RECT 13.195 0.36 13.335 0.42 ;
 RECT 13.53 1.055 13.83 1.195 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 5.36 0.805 5.5 1.22 ;
 RECT 5.185 1.82 7.39 1.96 ;
 RECT 7.25 1.58 7.39 1.82 ;
 RECT 5.185 1.36 5.325 1.82 ;
 RECT 9.305 0.805 9.445 1.72 ;
 RECT 9.305 1.9 9.515 1.905 ;
 RECT 9.235 1.86 9.515 1.9 ;
 RECT 9.305 1.72 11.495 1.76 ;
 RECT 9.235 1.76 11.495 1.86 ;
 RECT 11.915 1.92 12.055 2.505 ;
 RECT 11.195 1.86 11.495 1.935 ;
 RECT 11.355 1.935 11.495 2.505 ;
 RECT 11.355 2.505 12.055 2.645 ;
 RECT 10.21 1.86 10.44 2.055 ;
 RECT 12.15 1.245 12.29 1.78 ;
 RECT 12.15 1.105 12.53 1.245 ;
 RECT 11.915 1.78 12.29 1.92 ;
 END
END SDFFASRX1

MACRO SDFFASRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 14.72 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 14.72 2.96 ;
 RECT 7.265 2.635 7.525 2.8 ;
 RECT 8.285 2.38 8.425 2.8 ;
 RECT 11.075 2.21 11.215 2.8 ;
 RECT 12.195 2.06 12.335 2.8 ;
 RECT 14.195 1.485 14.335 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 3.18 1.93 3.32 2.8 ;
 RECT 4.025 1.93 4.165 2.8 ;
 RECT 13.25 1.485 13.39 2.8 ;
 RECT 1.27 1.985 1.41 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 14.72 0.08 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 3.88 0.08 4.11 0.39 ;
 RECT 10.545 0.08 10.8 1.005 ;
 RECT 6.525 0.08 6.76 0.37 ;
 RECT 13.38 0.08 13.615 0.37 ;
 RECT 12.215 0.08 12.355 0.565 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 14.475 0.08 14.615 0.86 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.195 0.97 10.335 1.16 ;
 RECT 5.92 0.51 7.075 0.65 ;
 RECT 10.195 1.16 11.485 1.3 ;
 RECT 6.935 0.36 7.075 0.51 ;
 RECT 9.415 0.36 9.8 0.63 ;
 RECT 6.935 0.22 9.8 0.36 ;
 RECT 9.66 0.63 9.8 0.83 ;
 RECT 9.66 0.83 10.335 0.97 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.615 2.04 2.015 2.415 ;
 RECT 2.575 1.86 2.715 1.89 ;
 RECT 1.875 1.72 2.715 1.86 ;
 RECT 2.575 1.615 2.715 1.72 ;
 RECT 1.875 1.86 2.015 2.04 ;
 RECT 1.875 1.11 2.015 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.2 1.16 2.715 1.43 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.945 0.33 10.26 0.685 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.78 1.425 12.92 2.575 ;
 RECT 12.78 1.105 13.09 1.425 ;
 RECT 12.78 0.5 12.92 1.105 ;
 END
 ANTENNADIFFAREA 0.672 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.72 2.015 14.045 2.38 ;
 RECT 13.72 0.6 14.21 0.74 ;
 RECT 13.72 2.38 13.86 2.58 ;
 RECT 13.72 0.74 13.86 2.015 ;
 END
 ANTENNADIFFAREA 0.568 ;
 END Q

 OBS
 LAYER PO ;
 RECT 3.78 1.44 4.025 1.52 ;
 RECT 3.78 1.62 4.025 1.69 ;
 RECT 4.28 1.21 5.245 1.31 ;
 RECT 8.62 0.635 8.72 1.35 ;
 RECT 10.375 0.265 10.475 1.22 ;
 RECT 8.62 0.265 8.72 0.535 ;
 RECT 7.635 0.46 7.865 0.535 ;
 RECT 7.635 0.535 8.72 0.635 ;
 RECT 7.635 0.635 7.865 0.69 ;
 RECT 9.065 1.545 9.165 2.195 ;
 RECT 8.62 0.165 10.475 0.265 ;
 RECT 8.62 1.35 8.91 1.445 ;
 RECT 8.62 1.445 9.165 1.45 ;
 RECT 8.81 1.45 9.165 1.545 ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 2.665 1.865 2.765 2.48 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 7.67 1.33 7.77 1.565 ;
 RECT 7.84 1.665 7.94 2.69 ;
 RECT 10.035 0.685 10.135 2.69 ;
 RECT 7.15 0.635 7.25 1.23 ;
 RECT 7.15 1.23 7.77 1.33 ;
 RECT 7.67 1.565 7.94 1.665 ;
 RECT 7.84 2.69 10.135 2.79 ;
 RECT 9.965 0.475 10.195 0.685 ;
 RECT 6.335 0.285 6.435 1.24 ;
 RECT 4.6 0.185 6.435 0.285 ;
 RECT 4.6 0.285 4.7 0.525 ;
 RECT 4.56 0.525 4.79 0.76 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.255 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 11.255 1.25 11.99 1.35 ;
 RECT 11.89 1.35 11.99 2.63 ;
 RECT 11.255 1.11 11.485 1.25 ;
 RECT 11.325 0.65 11.425 1.11 ;
 RECT 5.1 1.655 5.2 2.495 ;
 RECT 4.575 1.555 5.2 1.655 ;
 RECT 4.575 1.655 4.82 1.8 ;
 RECT 10.645 2.47 10.96 2.71 ;
 RECT 10.86 1.96 10.96 2.47 ;
 RECT 8.12 1.64 8.575 1.87 ;
 RECT 8.12 1.095 8.36 1.64 ;
 RECT 8.045 0.865 8.36 1.095 ;
 RECT 6.035 0.695 6.135 1.61 ;
 RECT 6.07 1.71 6.17 2.48 ;
 RECT 6.035 1.61 6.17 1.71 ;
 RECT 5.915 0.465 6.155 0.695 ;
 RECT 9.56 0.645 9.66 1.24 ;
 RECT 9.56 1.24 9.805 1.45 ;
 RECT 9.56 1.45 9.66 2.37 ;
 RECT 9.09 0.685 9.19 1.255 ;
 RECT 9.015 0.455 9.245 0.685 ;
 RECT 10.87 1.57 11.43 1.67 ;
 RECT 11.205 1.67 11.43 1.94 ;
 RECT 11.33 1.94 11.43 2.63 ;
 RECT 10.87 0.65 10.97 1.57 ;
 RECT 7.2 1.61 7.465 1.82 ;
 RECT 7.365 1.82 7.465 2.49 ;
 RECT 6.795 0.625 6.895 1.51 ;
 RECT 6.795 1.51 7.465 1.61 ;
 RECT 5.595 1.33 5.735 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.635 0.65 5.735 1.33 ;
 RECT 5.595 1.475 5.825 1.71 ;
 RECT 12.28 1.06 12.63 1.1 ;
 RECT 12.28 1.1 13.135 1.2 ;
 RECT 12.28 1.2 12.63 1.29 ;
 RECT 13.035 0.12 13.135 1.1 ;
 RECT 13.035 1.2 13.135 2.775 ;
 RECT 12.53 0.125 12.63 1.06 ;
 RECT 12.53 1.29 12.63 2.775 ;
 RECT 13.505 1.3 13.605 2.775 ;
 RECT 13.345 1.2 13.605 1.3 ;
 RECT 14.26 0.35 14.36 1.1 ;
 RECT 13.345 1.1 14.36 1.2 ;
 RECT 13.79 0.35 13.89 1.1 ;
 RECT 13.345 1.065 13.6 1.1 ;
 RECT 13.98 1.2 14.08 2.775 ;
 RECT 2.54 1.2 2.765 1.245 ;
 RECT 2.665 0.655 2.765 1.2 ;
 RECT 2.54 1.345 2.765 1.43 ;
 RECT 2.245 1.345 2.345 1.645 ;
 RECT 2.195 1.745 2.295 2.465 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.245 1.245 2.765 1.345 ;
 RECT 4.28 1.62 4.38 2.685 ;
 RECT 4.28 1.31 4.38 1.52 ;
 RECT 3.78 1.52 4.38 1.62 ;
 RECT 5.145 0.47 5.43 0.705 ;
 RECT 5.145 0.705 5.245 1.21 ;
 RECT 4.28 2.685 6.995 2.785 ;
 RECT 6.895 1.79 6.995 2.685 ;
 RECT 4.28 0.585 4.38 1.21 ;
 LAYER CO ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 4.63 1.6 4.76 1.73 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 3.305 1.535 3.435 1.665 ;
 RECT 3.66 1.995 3.79 2.125 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 1.995 3.315 2.125 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 13.43 0.23 13.56 0.36 ;
 RECT 13.255 1.555 13.385 1.685 ;
 RECT 13.255 2.35 13.385 2.48 ;
 RECT 13.255 1.825 13.385 1.955 ;
 RECT 13.255 2.085 13.385 2.215 ;
 RECT 4.5 2.015 4.63 2.145 ;
 RECT 5.25 0.525 5.38 0.655 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 2.58 1.25 2.71 1.38 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 10.71 2.525 10.84 2.655 ;
 RECT 8.815 1.815 8.945 1.945 ;
 RECT 8.29 2.44 8.42 2.57 ;
 RECT 14.01 0.605 14.14 0.735 ;
 RECT 12.785 0.55 12.915 0.68 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 8.395 1.69 8.525 1.82 ;
 RECT 10.62 0.87 10.75 1 ;
 RECT 7.685 0.51 7.815 0.64 ;
 RECT 9.78 2.02 9.91 2.15 ;
 RECT 8.84 0.87 8.97 1 ;
 RECT 9.065 0.505 9.195 0.635 ;
 RECT 9.62 1.28 9.75 1.41 ;
 RECT 11.64 0.87 11.77 1 ;
 RECT 11.08 2.28 11.21 2.41 ;
 RECT 10.61 2.19 10.74 2.32 ;
 RECT 12.2 2.13 12.33 2.26 ;
 RECT 11.64 2.13 11.77 2.26 ;
 RECT 11.255 1.76 11.385 1.89 ;
 RECT 7.255 1.63 7.385 1.76 ;
 RECT 5.645 1.525 5.775 1.655 ;
 RECT 7.59 0.88 7.72 1.01 ;
 RECT 7.585 2.015 7.715 2.145 ;
 RECT 3.93 0.255 4.06 0.385 ;
 RECT 7.315 2.64 7.445 2.77 ;
 RECT 6.645 2.105 6.775 2.235 ;
 RECT 10.015 0.515 10.145 0.645 ;
 RECT 14.48 0.68 14.61 0.81 ;
 RECT 13.385 1.115 13.515 1.245 ;
 RECT 12.33 1.11 12.46 1.24 ;
 RECT 12.785 1.825 12.915 1.955 ;
 RECT 12.785 2.085 12.915 2.215 ;
 RECT 12.22 0.365 12.35 0.495 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 8.115 0.915 8.245 1.045 ;
 RECT 11.305 1.165 11.435 1.295 ;
 RECT 5.97 0.515 6.1 0.645 ;
 RECT 6.575 0.23 6.705 0.36 ;
 RECT 9.31 1.765 9.44 1.895 ;
 RECT 9.31 0.87 9.44 1 ;
 RECT 10.26 1.92 10.39 2.05 ;
 RECT 14.2 1.555 14.33 1.685 ;
 RECT 14.2 2.35 14.33 2.48 ;
 RECT 14.2 1.825 14.33 1.955 ;
 RECT 14.2 2.085 14.33 2.215 ;
 RECT 13.725 1.555 13.855 1.685 ;
 RECT 13.725 2.35 13.855 2.48 ;
 RECT 13.725 1.825 13.855 1.955 ;
 RECT 13.725 2.085 13.855 2.215 ;
 RECT 12.785 1.555 12.915 1.685 ;
 RECT 12.785 2.35 12.915 2.48 ;
 RECT 6.295 1.825 6.425 1.955 ;
 RECT 5.815 2.105 5.945 2.235 ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 4.03 2.005 4.16 2.135 ;
 RECT 4.61 0.58 4.74 0.71 ;
 RECT 5.345 2.07 5.475 2.2 ;
 LAYER M1 ;
 RECT 5.18 0.52 5.78 0.66 ;
 RECT 5.64 0.66 5.78 0.79 ;
 RECT 5.64 0.79 7.355 0.93 ;
 RECT 7.215 0.505 7.89 0.645 ;
 RECT 7.215 0.645 7.355 0.79 ;
 RECT 5.745 2.1 6.845 2.24 ;
 RECT 9.425 2.32 9.565 2.52 ;
 RECT 7.925 2.18 9.495 2.185 ;
 RECT 7.925 2.185 9.565 2.24 ;
 RECT 8.78 2.24 9.565 2.32 ;
 RECT 4.495 2.43 8.065 2.435 ;
 RECT 7.925 1.35 8.065 2.1 ;
 RECT 7.925 2.24 8.065 2.295 ;
 RECT 6.985 2.295 8.065 2.43 ;
 RECT 4.495 2.435 7.125 2.57 ;
 RECT 8.48 0.5 9.27 0.64 ;
 RECT 7.925 2.1 8.92 2.18 ;
 RECT 8.48 0.64 8.62 1.21 ;
 RECT 7.925 1.21 8.62 1.35 ;
 RECT 4.495 1.78 4.635 2.43 ;
 RECT 4.495 0.84 4.745 1.035 ;
 RECT 4.605 0.51 4.745 0.84 ;
 RECT 4.495 1.035 4.635 1.55 ;
 RECT 4.495 1.55 4.765 1.78 ;
 RECT 9.425 2.52 10.92 2.66 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.365 2.11 2.995 2.25 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 3.46 0.53 4.41 0.67 ;
 RECT 4.89 0.36 5.03 1.175 ;
 RECT 4.905 1.27 5.045 2.1 ;
 RECT 4.27 0.36 4.41 0.53 ;
 RECT 4.27 0.22 5.03 0.36 ;
 RECT 4.78 2.1 5.05 2.24 ;
 RECT 4.89 1.175 5.045 1.27 ;
 RECT 3.7 1.63 3.84 1.925 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.655 1.925 3.84 2.175 ;
 RECT 3.7 1.475 4.045 1.63 ;
 RECT 7.52 0.875 8.315 1.05 ;
 RECT 7.58 1.325 7.72 2.01 ;
 RECT 6.97 1.185 7.72 1.325 ;
 RECT 7.52 1.05 7.72 1.185 ;
 RECT 5.575 1.52 7.11 1.66 ;
 RECT 6.97 1.325 7.11 1.52 ;
 RECT 7.53 2.01 7.785 2.15 ;
 RECT 9.615 1.21 9.755 1.44 ;
 RECT 11.635 0.82 12.635 0.965 ;
 RECT 12.495 0.36 12.635 0.82 ;
 RECT 13.09 0.36 13.23 0.67 ;
 RECT 12.495 0.22 13.23 0.36 ;
 RECT 11.635 0.965 11.775 1.44 ;
 RECT 11.635 1.58 11.775 2.33 ;
 RECT 9.615 1.44 11.775 1.58 ;
 RECT 13.25 0.81 13.39 1.11 ;
 RECT 13.25 1.11 13.58 1.25 ;
 RECT 13.09 0.67 13.39 0.81 ;
 RECT 9.775 2.155 9.96 2.22 ;
 RECT 9.775 2 9.915 2.015 ;
 RECT 10.555 2.185 10.795 2.22 ;
 RECT 9.775 2.22 10.795 2.36 ;
 RECT 9.73 2.015 9.96 2.155 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 5.36 0.805 5.5 1.22 ;
 RECT 5.185 1.82 7.39 1.96 ;
 RECT 7.25 1.58 7.39 1.82 ;
 RECT 5.185 1.36 5.325 1.82 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 9.305 0.805 9.445 1.72 ;
 RECT 9.305 1.9 9.515 1.905 ;
 RECT 9.235 1.86 9.515 1.9 ;
 RECT 9.305 1.72 11.495 1.76 ;
 RECT 9.235 1.76 11.495 1.86 ;
 RECT 11.915 1.92 12.055 2.505 ;
 RECT 11.355 1.935 11.495 2.505 ;
 RECT 11.195 1.86 11.495 1.935 ;
 RECT 11.355 2.505 12.055 2.645 ;
 RECT 10.21 1.86 10.44 2.055 ;
 RECT 12.15 1.245 12.29 1.78 ;
 RECT 12.15 1.105 12.53 1.245 ;
 RECT 11.915 1.78 12.29 1.92 ;
 RECT 8.835 1.005 8.975 1.685 ;
 RECT 8.325 1.685 8.975 1.81 ;
 RECT 8.325 1.81 9.015 1.825 ;
 RECT 8.745 1.825 9.015 1.95 ;
 RECT 8.765 0.865 9.045 1.005 ;
 END
END SDFFASRX2

MACRO SDFFASX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 12.8 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 12.8 2.96 ;
 RECT 1.51 2.025 1.65 2.8 ;
 RECT 4.075 2.36 4.325 2.8 ;
 RECT 6.415 2.635 6.675 2.8 ;
 RECT 11.855 1.48 11.995 2.8 ;
 RECT 7.405 2.38 7.545 2.8 ;
 RECT 3.42 2 3.56 2.8 ;
 RECT 0.54 1.76 0.68 2.8 ;
 RECT 10.18 2.055 10.32 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 12.8 0.08 ;
 RECT 3.995 0.08 4.225 0.385 ;
 RECT 11.95 0.08 12.09 0.76 ;
 RECT 3.42 0.08 3.56 0.53 ;
 RECT 6.385 0.08 6.525 0.38 ;
 RECT 0.54 0.08 0.68 0.83 ;
 RECT 9.695 0.08 9.835 1.07 ;
 RECT 1.51 0.08 1.65 1.075 ;
 END
 END VSS

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.96 0.325 9.285 0.735 ;
 END
 ANTENNAGATEAREA 0.088 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.19 0.52 11.525 0.77 ;
 RECT 11.3 0.77 11.44 2.51 ;
 END
 ANTENNADIFFAREA 0.611 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.2 2.065 12.475 2.385 ;
 RECT 12.335 0.77 12.56 0.91 ;
 RECT 12.42 0.555 12.56 0.77 ;
 RECT 12.335 2.385 12.475 2.52 ;
 RECT 12.335 0.91 12.475 2.065 ;
 END
 ANTENNADIFFAREA 0.466 ;
 END Q

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.515 1.5 1.925 1.88 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.9 2.115 2.255 2.385 ;
 RECT 2.815 1.655 2.955 1.74 ;
 RECT 2.115 1.74 2.955 1.91 ;
 RECT 2.115 1.91 2.255 2.115 ;
 RECT 2.115 1.13 2.255 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.4 1.415 2.86 1.505 ;
 RECT 2.4 1.505 2.67 1.6 ;
 RECT 2.405 1.17 2.86 1.415 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.52 1.47 3.885 1.805 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 OBS
 LAYER PO ;
 RECT 5.34 1.77 5.44 2.495 ;
 RECT 8.665 0.645 8.765 1.24 ;
 RECT 8.665 1.24 8.91 1.45 ;
 RECT 8.665 1.45 8.765 2.37 ;
 RECT 8.195 0.685 8.295 1.23 ;
 RECT 8.12 0.455 8.35 0.685 ;
 RECT 7.725 0.265 7.825 0.575 ;
 RECT 7.075 0.575 7.825 0.675 ;
 RECT 7.725 0.675 7.825 1.35 ;
 RECT 8.17 1.545 8.27 2.415 ;
 RECT 9.48 0.265 9.58 1.32 ;
 RECT 7.075 0.455 7.305 0.575 ;
 RECT 7.075 0.675 7.305 0.685 ;
 RECT 7.915 1.45 8.27 1.545 ;
 RECT 7.725 0.165 9.58 0.265 ;
 RECT 7.725 1.35 8.015 1.445 ;
 RECT 7.725 1.445 8.27 1.45 ;
 RECT 10.31 1.63 10.535 1.94 ;
 RECT 10.435 1.94 10.535 2.66 ;
 RECT 9.95 0.65 10.05 1.53 ;
 RECT 9.95 1.53 10.535 1.63 ;
 RECT 12.205 0.215 12.305 1.035 ;
 RECT 12.115 1.27 12.215 2.79 ;
 RECT 11.955 1.035 12.305 1.27 ;
 RECT 11.565 0.145 11.665 1.18 ;
 RECT 11.565 1.28 11.665 2.79 ;
 RECT 10.985 1.18 11.665 1.28 ;
 RECT 10.985 1.28 11.195 1.415 ;
 RECT 2.1 0.66 2.2 1.165 ;
 RECT 2.06 1.165 2.305 1.405 ;
 RECT 3 0.195 3.305 0.425 ;
 RECT 3.205 0.425 3.305 2.485 ;
 RECT 3.68 0.675 3.78 1.5 ;
 RECT 3.485 1.5 3.78 1.74 ;
 RECT 3.68 1.74 3.78 2.39 ;
 RECT 7.1 1.375 7.2 2.69 ;
 RECT 6.795 1.275 7.2 1.375 ;
 RECT 7.1 2.69 9.24 2.79 ;
 RECT 9.14 0.73 9.24 2.69 ;
 RECT 6.795 0.635 6.895 1.275 ;
 RECT 9.01 0.52 9.24 0.73 ;
 RECT 7.38 1.64 7.76 1.87 ;
 RECT 7.38 1.095 7.545 1.64 ;
 RECT 7.275 0.865 7.545 1.095 ;
 RECT 4.455 1.69 4.555 2.685 ;
 RECT 4.455 1.355 4.555 1.44 ;
 RECT 5.385 0.705 5.485 1.255 ;
 RECT 6.14 1.795 6.24 2.685 ;
 RECT 5.385 0.47 5.67 0.705 ;
 RECT 4.455 2.685 6.24 2.785 ;
 RECT 4.455 1.255 5.485 1.355 ;
 RECT 4.205 1.44 4.555 1.69 ;
 RECT 4.52 0.515 4.62 1.255 ;
 RECT 6.495 0.625 6.595 1.58 ;
 RECT 6.625 1.82 6.725 2.39 ;
 RECT 6.495 1.58 6.735 1.82 ;
 RECT 5.835 1.43 5.935 1.475 ;
 RECT 5.835 1.71 5.935 2.505 ;
 RECT 5.855 0.65 5.955 1.33 ;
 RECT 5.835 1.33 5.955 1.43 ;
 RECT 5.705 1.475 5.935 1.71 ;
 RECT 2.485 1.43 2.585 1.665 ;
 RECT 2.905 0.675 3.005 1.2 ;
 RECT 2.435 1.765 2.535 2.49 ;
 RECT 2.435 1.665 2.585 1.765 ;
 RECT 2.485 1.2 3.005 1.43 ;
 RECT 6.17 0.285 6.27 1.24 ;
 RECT 4.84 0.185 6.27 0.285 ;
 RECT 4.84 0.285 4.94 0.5 ;
 RECT 4.8 0.5 5.03 0.735 ;
 RECT 2.905 1.885 3.005 2.5 ;
 RECT 2.765 1.655 3.005 1.885 ;
 RECT 9.75 2.47 10.065 2.71 ;
 RECT 9.965 1.88 10.065 2.47 ;
 RECT 1.295 1.495 1.865 1.77 ;
 RECT 1.295 0.655 1.395 1.495 ;
 RECT 1.295 1.77 1.395 2.485 ;
 RECT 1.765 0.675 1.865 1.495 ;
 RECT 1.765 1.77 1.865 2.485 ;
 RECT 4.735 1.67 5.44 1.77 ;
 RECT 4.735 1.77 4.98 1.92 ;
 LAYER CO ;
 RECT 7.015 0.88 7.145 1.01 ;
 RECT 11.305 1.53 11.435 1.66 ;
 RECT 6.39 0.2 6.52 0.33 ;
 RECT 4.675 2.23 4.805 2.36 ;
 RECT 5.49 0.525 5.62 0.655 ;
 RECT 8.4 1.815 8.53 1.945 ;
 RECT 8.415 0.87 8.545 1 ;
 RECT 9.365 1.965 9.495 2.095 ;
 RECT 8.885 1.965 9.015 2.095 ;
 RECT 12.34 1.53 12.47 1.66 ;
 RECT 12.34 1.79 12.47 1.92 ;
 RECT 12.34 2.05 12.47 2.18 ;
 RECT 12.34 2.31 12.47 2.44 ;
 RECT 11.86 1.53 11.99 1.66 ;
 RECT 11.86 1.79 11.99 1.92 ;
 RECT 11.86 2.05 11.99 2.18 ;
 RECT 11.86 2.31 11.99 2.44 ;
 RECT 11.305 2.05 11.435 2.18 ;
 RECT 11.305 2.31 11.435 2.44 ;
 RECT 10.745 2.13 10.875 2.26 ;
 RECT 11.995 1.085 12.125 1.215 ;
 RECT 12.425 0.625 12.555 0.755 ;
 RECT 11.955 0.56 12.085 0.69 ;
 RECT 7.58 1.69 7.71 1.82 ;
 RECT 2.12 1.215 2.25 1.345 ;
 RECT 0.545 0.37 0.675 0.5 ;
 RECT 1.515 2.075 1.645 2.205 ;
 RECT 1.52 1.57 1.65 1.7 ;
 RECT 2.82 1.705 2.95 1.835 ;
 RECT 3.425 2.07 3.555 2.2 ;
 RECT 4.275 1.495 4.405 1.625 ;
 RECT 4.145 2.365 4.275 2.495 ;
 RECT 5.585 2.07 5.715 2.2 ;
 RECT 0.545 2.365 0.675 2.495 ;
 RECT 3.9 2.015 4.03 2.145 ;
 RECT 1.515 0.895 1.645 1.025 ;
 RECT 10.36 1.76 10.49 1.89 ;
 RECT 6.565 1.63 6.695 1.76 ;
 RECT 5.755 1.525 5.885 1.655 ;
 RECT 6.85 2.015 6.98 2.145 ;
 RECT 4.045 0.25 4.175 0.38 ;
 RECT 6.465 2.64 6.595 2.77 ;
 RECT 9.7 0.87 9.83 1 ;
 RECT 0.545 0.63 0.675 0.76 ;
 RECT 0.545 1.845 0.675 1.975 ;
 RECT 5.605 0.88 5.735 1.01 ;
 RECT 5.09 2.105 5.22 2.235 ;
 RECT 5.135 0.88 5.265 1.01 ;
 RECT 0.545 2.105 0.675 2.235 ;
 RECT 4.03 0.895 4.16 1.025 ;
 RECT 4.85 0.555 4.98 0.685 ;
 RECT 4.805 1.725 4.935 1.855 ;
 RECT 1.045 2.075 1.175 2.205 ;
 RECT 1.045 0.895 1.175 1.025 ;
 RECT 9.815 2.525 9.945 2.655 ;
 RECT 4.74 0.905 4.87 1.035 ;
 RECT 11.305 0.585 11.435 0.715 ;
 RECT 7.945 0.87 8.075 1 ;
 RECT 8.17 0.505 8.3 0.635 ;
 RECT 8.725 1.28 8.855 1.41 ;
 RECT 10.17 0.87 10.3 1 ;
 RECT 10.185 2.115 10.315 2.245 ;
 RECT 9.715 2.11 9.845 2.24 ;
 RECT 11.305 1.79 11.435 1.92 ;
 RECT 7.92 1.815 8.05 1.945 ;
 RECT 7.41 2.44 7.54 2.57 ;
 RECT 7.34 0.915 7.47 1.045 ;
 RECT 7.125 0.505 7.255 0.635 ;
 RECT 11.025 1.23 11.155 1.36 ;
 RECT 3.425 0.265 3.555 0.395 ;
 RECT 3.05 0.245 3.18 0.375 ;
 RECT 3.535 1.555 3.665 1.685 ;
 RECT 2.46 0.895 2.59 1.025 ;
 RECT 2.655 2.135 2.785 2.265 ;
 RECT 2.64 1.25 2.77 1.38 ;
 RECT 9.06 0.56 9.19 0.69 ;
 LAYER M1 ;
 RECT 5.42 0.52 7.33 0.66 ;
 RECT 7.045 0.47 7.33 0.52 ;
 RECT 5.425 1.805 6.7 1.945 ;
 RECT 5.425 1.945 5.79 1.96 ;
 RECT 5.425 1.22 5.74 1.36 ;
 RECT 5.6 0.805 5.74 1.22 ;
 RECT 5.51 1.96 5.79 2.215 ;
 RECT 5.425 1.36 5.565 1.805 ;
 RECT 6.56 1.56 6.7 1.805 ;
 RECT 10.74 1.005 10.88 1.395 ;
 RECT 8.72 1.395 10.88 1.535 ;
 RECT 10.74 1.535 10.88 2.32 ;
 RECT 10.74 0.38 10.88 0.865 ;
 RECT 10.12 0.865 10.88 1.005 ;
 RECT 8.72 1.21 8.86 1.395 ;
 RECT 11.67 0.38 11.81 1.15 ;
 RECT 10.74 0.24 11.81 0.38 ;
 RECT 11.99 1.02 12.13 1.15 ;
 RECT 11.67 1.15 12.13 1.29 ;
 RECT 1.825 0.38 1.965 1.22 ;
 RECT 1.04 1.22 1.965 1.36 ;
 RECT 1.04 0.82 1.18 1.22 ;
 RECT 1.04 1.36 1.18 2.325 ;
 RECT 1.825 0.24 3.25 0.38 ;
 RECT 8.41 0.805 8.55 1.675 ;
 RECT 9.315 1.815 9.545 2.1 ;
 RECT 8.34 1.815 8.62 1.95 ;
 RECT 8.34 1.675 10.6 1.815 ;
 RECT 11.02 1.18 11.16 2.505 ;
 RECT 10.3 1.815 10.6 1.915 ;
 RECT 10.46 1.915 10.6 2.505 ;
 RECT 10.46 2.505 11.16 2.645 ;
 RECT 8.88 2.1 9.065 2.24 ;
 RECT 9.71 2.03 9.85 2.24 ;
 RECT 8.835 1.96 9.065 2.1 ;
 RECT 8.88 2.24 9.85 2.38 ;
 RECT 7.57 1.685 8.08 1.81 ;
 RECT 7.57 1.81 8.12 1.825 ;
 RECT 7.94 0.78 8.08 1.685 ;
 RECT 7.57 1.615 7.71 1.685 ;
 RECT 7.57 1.825 7.71 1.895 ;
 RECT 7.85 1.825 8.12 1.95 ;
 RECT 6.845 1.04 7.52 1.05 ;
 RECT 6.28 0.91 7.52 1.04 ;
 RECT 6.28 0.9 7.15 0.91 ;
 RECT 6.845 1.08 6.985 2.2 ;
 RECT 6.845 1.05 7.15 1.08 ;
 RECT 5.705 1.52 6.42 1.66 ;
 RECT 7.01 0.81 7.15 0.9 ;
 RECT 6.28 1.04 6.42 1.52 ;
 RECT 4.025 0.845 4.165 1.125 ;
 RECT 4.025 1.125 4.41 1.265 ;
 RECT 4.27 1.265 4.41 2.01 ;
 RECT 3.83 2.01 4.41 2.15 ;
 RECT 7.125 1.36 7.265 2.1 ;
 RECT 7.125 2.24 7.265 2.355 ;
 RECT 6.05 2.355 7.265 2.495 ;
 RECT 4.67 2.515 6.19 2.655 ;
 RECT 4.735 0.735 4.875 1.72 ;
 RECT 4.735 1.72 4.985 1.775 ;
 RECT 4.67 1.775 4.985 1.86 ;
 RECT 4.67 1.86 4.875 2.005 ;
 RECT 4.67 2.005 4.81 2.515 ;
 RECT 4.845 0.505 4.985 0.535 ;
 RECT 6.05 2.495 6.19 2.515 ;
 RECT 4.735 0.535 4.985 0.735 ;
 RECT 7.125 2.185 8.67 2.24 ;
 RECT 7.125 2.1 8.66 2.185 ;
 RECT 8.53 2.24 8.67 2.52 ;
 RECT 7.66 0.5 8.375 0.64 ;
 RECT 7.66 0.64 7.8 1.22 ;
 RECT 7.125 1.22 7.8 1.36 ;
 RECT 8.53 2.52 10.025 2.66 ;
 RECT 3.7 0.665 3.84 0.895 ;
 RECT 2.395 0.895 3.84 1.03 ;
 RECT 3.095 1.03 3.84 1.035 ;
 RECT 3.095 1.035 3.235 2.13 ;
 RECT 2.395 0.89 3.235 0.895 ;
 RECT 2.585 2.13 3.235 2.27 ;
 RECT 3.7 0.525 4.59 0.665 ;
 RECT 4.45 0.36 4.59 0.525 ;
 RECT 5.13 0.36 5.27 0.875 ;
 RECT 5.145 1.015 5.285 2.035 ;
 RECT 4.45 0.22 5.27 0.36 ;
 RECT 5.085 0.875 5.34 1.015 ;
 RECT 5.085 2.035 5.285 2.305 ;
 END
END SDFFASX1

MACRO INVX16
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.96 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 4.345 0.08 4.485 0.77 ;
 RECT 3.405 0.08 3.545 0.77 ;
 RECT 2.465 0.08 2.605 0.77 ;
 RECT 1.525 0.08 1.665 0.77 ;
 RECT 7.165 0.08 7.305 0.77 ;
 RECT 5.285 0.08 5.425 0.77 ;
 RECT 6.225 0.08 6.365 0.77 ;
 RECT 0.585 0.08 0.725 0.77 ;
 RECT 8.375 0.08 8.515 0.77 ;
 RECT 0 -0.08 8.96 0.08 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.065 1.37 7.34 1.72 ;
 RECT 0.305 1.23 7.495 1.37 ;
 END
 ANTENNAGATEAREA 2.576 ;
 END INP

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.755 1.715 6.835 1.855 ;
 RECT 3.875 1.715 4.955 1.855 ;
 RECT 1.995 1.715 3.075 1.855 ;
 RECT 0.115 1.715 1.195 1.855 ;
 RECT 7.635 1.13 8.185 1.43 ;
 RECT 6.695 0.625 6.835 0.94 ;
 RECT 6.695 1.86 7.775 2 ;
 RECT 5.755 0.64 5.895 0.94 ;
 RECT 4.815 0.625 4.955 0.94 ;
 RECT 2.935 0.625 3.075 0.94 ;
 RECT 3.875 0.64 4.015 0.94 ;
 RECT 5.755 1.585 5.895 1.715 ;
 RECT 6.695 1.855 6.835 1.86 ;
 RECT 1.995 0.64 2.135 0.94 ;
 RECT 1.055 0.625 1.195 0.94 ;
 RECT 0.115 0.64 0.255 0.94 ;
 RECT 4.815 1.86 5.895 2 ;
 RECT 3.875 1.585 4.015 1.715 ;
 RECT 4.815 1.855 4.955 1.86 ;
 RECT 2.935 1.86 4.015 2 ;
 RECT 2.935 2 3.075 2.31 ;
 RECT 1.995 1.585 2.135 1.715 ;
 RECT 2.935 1.855 3.075 1.86 ;
 RECT 1.055 1.86 2.135 2 ;
 RECT 1.055 1.855 1.195 1.86 ;
 RECT 0.115 1.855 0.255 2.31 ;
 RECT 7.635 1.08 7.775 1.13 ;
 RECT 7.635 0.64 7.775 0.94 ;
 RECT 0.115 0.94 7.775 1.08 ;
 RECT 6.695 2 6.835 2.31 ;
 RECT 7.635 2 7.775 2.04 ;
 RECT 7.635 1.43 7.775 1.86 ;
 RECT 5.755 1.855 5.895 1.86 ;
 RECT 5.755 2 5.895 2.31 ;
 RECT 4.815 2 4.955 2.31 ;
 RECT 3.875 1.855 4.015 1.86 ;
 RECT 3.875 2 4.015 2.31 ;
 RECT 1.995 1.855 2.135 1.86 ;
 RECT 1.995 2 2.135 2.31 ;
 RECT 1.055 2 1.195 2.31 ;
 END
 ANTENNADIFFAREA 5.138 ;
 END ZN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 3.405 2.345 3.545 2.8 ;
 RECT 5.285 2.345 5.425 2.8 ;
 RECT 1.525 2.345 1.665 2.8 ;
 RECT 7.165 2.345 7.305 2.8 ;
 RECT 4.345 2.065 4.485 2.8 ;
 RECT 2.465 2.065 2.605 2.8 ;
 RECT 6.225 2.065 6.365 2.8 ;
 RECT 0.585 2.065 0.725 2.8 ;
 RECT 8.37 1.915 8.51 2.8 ;
 RECT 0 2.8 8.96 2.96 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 3.66 0.275 3.76 1.185 ;
 RECT 3.505 1.185 3.76 1.415 ;
 RECT 3.66 1.415 3.76 2.79 ;
 RECT 3.19 0.275 3.29 1.185 ;
 RECT 3.19 1.415 3.29 2.79 ;
 RECT 3.095 1.185 3.325 1.415 ;
 RECT 2.72 0.275 2.82 1.185 ;
 RECT 2.72 1.415 2.82 2.79 ;
 RECT 2.685 1.185 2.915 1.415 ;
 RECT 2.25 0.275 2.35 1.185 ;
 RECT 2.25 1.185 2.505 1.415 ;
 RECT 2.25 1.415 2.35 2.79 ;
 RECT 1.78 0.275 1.88 1.185 ;
 RECT 1.625 1.185 1.88 1.415 ;
 RECT 1.78 1.415 1.88 2.79 ;
 RECT 1.31 0.275 1.41 1.185 ;
 RECT 1.31 1.415 1.41 2.79 ;
 RECT 1.2 1.185 1.43 1.415 ;
 RECT 0.37 0.275 0.47 1.185 ;
 RECT 0.37 1.415 0.47 2.79 ;
 RECT 0.305 1.185 0.535 1.415 ;
 RECT 5.54 0.275 5.64 1.185 ;
 RECT 5.385 1.185 5.64 1.415 ;
 RECT 5.54 1.415 5.64 2.79 ;
 RECT 5.07 0.275 5.17 1.185 ;
 RECT 5.07 1.415 5.17 2.79 ;
 RECT 4.96 1.185 5.19 1.415 ;
 RECT 6.01 0.275 6.11 1.185 ;
 RECT 6.01 1.185 6.265 1.415 ;
 RECT 6.01 1.415 6.11 2.79 ;
 RECT 4.13 0.275 4.23 1.185 ;
 RECT 4.13 1.185 4.745 1.415 ;
 RECT 4.13 1.415 4.23 2.79 ;
 RECT 4.6 0.275 4.7 1.185 ;
 RECT 4.6 1.415 4.7 2.79 ;
 RECT 7.42 0.275 7.52 1.185 ;
 RECT 7.265 1.185 7.52 1.415 ;
 RECT 7.42 1.415 7.52 2.79 ;
 RECT 6.95 0.275 7.05 1.185 ;
 RECT 6.95 1.415 7.05 2.79 ;
 RECT 6.855 1.185 7.085 1.415 ;
 RECT 0.84 0.275 0.94 1.185 ;
 RECT 0.84 1.415 0.94 2.79 ;
 RECT 0.755 1.185 0.985 1.415 ;
 RECT 6.48 0.275 6.58 1.185 ;
 RECT 6.48 1.415 6.58 2.79 ;
 RECT 6.445 1.185 6.675 1.415 ;
 LAYER CO ;
 RECT 3.88 1.86 4.01 1.99 ;
 RECT 2.47 2.115 2.6 2.245 ;
 RECT 2.94 2.13 3.07 2.26 ;
 RECT 3.555 1.235 3.685 1.365 ;
 RECT 3.145 1.235 3.275 1.365 ;
 RECT 2.735 1.235 2.865 1.365 ;
 RECT 2.325 1.235 2.455 1.365 ;
 RECT 0.59 0.59 0.72 0.72 ;
 RECT 5.29 0.59 5.42 0.72 ;
 RECT 0.59 2.425 0.72 2.555 ;
 RECT 0.355 1.235 0.485 1.365 ;
 RECT 0.805 1.235 0.935 1.365 ;
 RECT 0.12 2.13 0.25 2.26 ;
 RECT 1.53 2.44 1.66 2.57 ;
 RECT 1.675 1.235 1.805 1.365 ;
 RECT 2 1.86 2.13 1.99 ;
 RECT 1.06 1.86 1.19 1.99 ;
 RECT 1.25 1.235 1.38 1.365 ;
 RECT 6.7 0.675 6.83 0.805 ;
 RECT 0.12 1.86 0.25 1.99 ;
 RECT 0.59 2.115 0.72 2.245 ;
 RECT 2 0.69 2.13 0.82 ;
 RECT 0.12 0.69 0.25 0.82 ;
 RECT 1.06 2.13 1.19 2.26 ;
 RECT 1.53 0.59 1.66 0.72 ;
 RECT 7.17 0.59 7.3 0.72 ;
 RECT 3.88 1.86 4.01 1.99 ;
 RECT 3.88 0.69 4.01 0.82 ;
 RECT 6.23 2.425 6.36 2.555 ;
 RECT 5.76 1.86 5.89 1.99 ;
 RECT 4.35 2.115 4.48 2.245 ;
 RECT 4.82 2.13 4.95 2.26 ;
 RECT 5.435 1.235 5.565 1.365 ;
 RECT 5.01 1.235 5.14 1.365 ;
 RECT 4.565 1.235 4.695 1.365 ;
 RECT 6.495 1.235 6.625 1.365 ;
 RECT 6.085 1.235 6.215 1.365 ;
 RECT 6.7 1.86 6.83 1.99 ;
 RECT 5.76 1.86 5.89 1.99 ;
 RECT 7.64 0.69 7.77 0.82 ;
 RECT 5.76 0.69 5.89 0.82 ;
 RECT 6.23 0.59 6.36 0.72 ;
 RECT 2 1.86 2.13 1.99 ;
 RECT 7.64 1.86 7.77 1.99 ;
 RECT 4.82 1.86 4.95 1.99 ;
 RECT 4.35 0.59 4.48 0.72 ;
 RECT 3.88 2.13 4.01 2.26 ;
 RECT 7.17 2.44 7.3 2.57 ;
 RECT 6.23 2.115 6.36 2.245 ;
 RECT 5.76 2.13 5.89 2.26 ;
 RECT 5.76 0.69 5.89 0.82 ;
 RECT 6.7 2.13 6.83 2.26 ;
 RECT 4.82 0.675 4.95 0.805 ;
 RECT 5.29 2.44 5.42 2.57 ;
 RECT 4.35 2.425 4.48 2.555 ;
 RECT 4.205 1.235 4.335 1.365 ;
 RECT 2.94 1.86 3.07 1.99 ;
 RECT 2.47 0.59 2.6 0.72 ;
 RECT 2 2.13 2.13 2.26 ;
 RECT 3.88 0.69 4.01 0.82 ;
 RECT 2.94 0.675 3.07 0.805 ;
 RECT 3.41 2.44 3.54 2.57 ;
 RECT 3.41 0.59 3.54 0.72 ;
 RECT 2.47 2.425 2.6 2.555 ;
 RECT 1.06 0.675 1.19 0.805 ;
 RECT 2 0.69 2.13 0.82 ;
 RECT 8.38 0.59 8.51 0.72 ;
 RECT 8.38 0.32 8.51 0.45 ;
 RECT 8.375 2.235 8.505 2.365 ;
 RECT 8.375 1.965 8.505 2.095 ;
 RECT 7.315 1.235 7.445 1.365 ;
 RECT 6.905 1.235 7.035 1.365 ;
 END
END INVX16

MACRO INVX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.24 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.24 2.96 ;
 RECT 1.75 1.92 1.89 2.8 ;
 RECT 0.74 1.91 0.88 2.8 ;
 END
 END VDD

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.545 1.085 1.08 1.4 ;
 END
 ANTENNAGATEAREA 0.322 ;
 END INP

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.24 0.08 ;
 RECT 0.74 0.08 0.88 0.86 ;
 RECT 1.745 0.08 1.885 0.795 ;
 END
 END VSS

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.23 1.1 1.625 1.485 ;
 RECT 1.23 0.64 1.37 1.1 ;
 RECT 1.23 1.485 1.37 1.545 ;
 RECT 0.25 1.685 0.39 2.14 ;
 RECT 0.25 0.64 0.39 1.545 ;
 RECT 1.23 1.685 1.37 1.87 ;
 RECT 0.25 1.545 1.37 1.685 ;
 END
 ANTENNADIFFAREA 0.966 ;
 END ZN

 OBS
 LAYER PO ;
 RECT 0.505 0.275 0.605 0.975 ;
 RECT 1.015 0.275 1.115 0.975 ;
 RECT 0.505 0.82 0.605 2.74 ;
 RECT 1.015 0.82 1.115 2.74 ;
 RECT 0.555 1.125 1.07 1.355 ;
 LAYER CO ;
 RECT 1.755 1.97 1.885 2.1 ;
 RECT 1.755 2.24 1.885 2.37 ;
 RECT 1.75 0.345 1.88 0.475 ;
 RECT 1.75 0.615 1.88 0.745 ;
 RECT 0.6 1.175 0.73 1.305 ;
 RECT 0.89 1.175 1.02 1.305 ;
 RECT 0.745 1.96 0.875 2.09 ;
 RECT 0.255 1.69 0.385 1.82 ;
 RECT 0.255 0.69 0.385 0.82 ;
 RECT 0.255 1.96 0.385 2.09 ;
 RECT 0.745 2.27 0.875 2.4 ;
 RECT 1.235 1.69 1.365 1.82 ;
 RECT 0.745 0.68 0.875 0.81 ;
 RECT 0.745 1.96 0.875 2.09 ;
 RECT 1.235 0.69 1.365 0.82 ;
 RECT 0.745 2.27 0.875 2.4 ;
 RECT 0.89 1.175 1.02 1.305 ;
 END
END INVX2

MACRO SDFFNARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 13.76 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 13.76 2.96 ;
 RECT 3.785 2.62 4.035 2.8 ;
 RECT 7.265 2.635 7.525 2.8 ;
 RECT 1.27 2.005 1.41 2.8 ;
 RECT 11.095 2.06 11.235 2.8 ;
 RECT 13.235 1.73 13.375 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 12.23 1.465 12.37 2.8 ;
 RECT 3.18 1.98 3.32 2.8 ;
 RECT 9.915 2.09 10.055 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 13.76 0.08 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 6.525 0.08 6.76 0.37 ;
 RECT 11.115 0.08 11.255 0.815 ;
 RECT 0.3 0.08 0.44 0.81 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 12.365 0.08 12.505 0.3 ;
 RECT 3.925 0.08 4.065 0.39 ;
 RECT 9.99 0.08 10.13 0.58 ;
 RECT 13.515 0.08 13.655 0.88 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.57 0.785 10.545 0.925 ;
 RECT 10.405 0.225 10.545 0.785 ;
 RECT 5.965 0.51 7.04 0.65 ;
 RECT 9.265 0.36 9.71 0.64 ;
 RECT 9.57 0.64 9.71 0.785 ;
 RECT 6.9 0.36 7.04 0.51 ;
 RECT 5.965 0.35 6.105 0.51 ;
 RECT 6.9 0.22 9.71 0.36 ;
 END
 ANTENNAGATEAREA 0.177 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.192 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.555 2.105 2.015 2.365 ;
 RECT 2.575 1.785 2.715 1.825 ;
 RECT 1.875 1.615 2.715 1.785 ;
 RECT 2.575 1.55 2.715 1.615 ;
 RECT 1.875 1.785 2.015 2.105 ;
 RECT 1.875 1.11 2.015 1.615 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.245 1.15 2.715 1.39 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.76 0.72 11.9 2.07 ;
 RECT 11.565 2.07 11.9 2.57 ;
 END
 ANTENNADIFFAREA 0.544 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.645 2.015 12.955 2.38 ;
 RECT 12.7 2.38 12.84 2.61 ;
 RECT 12.7 0.98 13.085 1.12 ;
 RECT 12.7 1.12 12.84 2.015 ;
 RECT 12.945 0.72 13.085 0.98 ;
 END
 ANTENNADIFFAREA 0.652 ;
 END Q

 OBS
 LAYER PO ;
 RECT 4.215 1.62 4.315 2.265 ;
 RECT 4.28 0.09 6.435 0.19 ;
 RECT 6.335 0.19 6.435 1.155 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.79 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.79 ;
 RECT 2.665 0.655 2.765 1.13 ;
 RECT 2.245 1.245 2.775 1.36 ;
 RECT 2.245 1.36 2.345 1.645 ;
 RECT 2.255 1.13 2.775 1.245 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.195 1.745 2.295 2.79 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 2.965 0.405 3.065 2.79 ;
 RECT 2.525 1.56 2.765 1.79 ;
 RECT 2.665 1.79 2.765 2.79 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 8.155 1.105 8.255 1.64 ;
 RECT 7.86 0.875 8.255 1.105 ;
 RECT 8.155 1.64 8.39 1.87 ;
 RECT 6.895 1.53 6.995 2.69 ;
 RECT 4.495 2.69 6.995 2.78 ;
 RECT 4.495 2.07 4.725 2.69 ;
 RECT 4.555 2.78 6.995 2.79 ;
 RECT 5.635 0.56 5.735 1.27 ;
 RECT 5.595 1.505 5.695 2.51 ;
 RECT 5.595 1.27 5.825 1.505 ;
 RECT 11.545 1.42 11.645 2.79 ;
 RECT 11.18 1.235 11.645 1.42 ;
 RECT 11.18 1.19 12.115 1.235 ;
 RECT 11.545 1.135 12.115 1.19 ;
 RECT 12.015 0.2 12.115 1.135 ;
 RECT 12.015 1.235 12.115 2.79 ;
 RECT 11.545 0.2 11.645 1.135 ;
 RECT 5.145 0.605 5.245 1.155 ;
 RECT 5.145 0.37 5.43 0.605 ;
 RECT 4.56 1.085 4.805 1.155 ;
 RECT 4.56 1.265 4.805 1.325 ;
 RECT 4.56 1.155 5.245 1.265 ;
 RECT 10.19 0.65 10.29 1.51 ;
 RECT 10.19 1.75 10.29 2.79 ;
 RECT 10.07 1.51 10.3 1.75 ;
 RECT 7.2 1.41 7.465 1.64 ;
 RECT 7.365 1.23 7.465 1.41 ;
 RECT 6.995 0.525 7.095 1.13 ;
 RECT 6.995 1.13 7.465 1.23 ;
 RECT 7.365 1.64 7.465 2.52 ;
 RECT 10.79 1.32 10.89 2.79 ;
 RECT 10.49 0.47 10.59 1.22 ;
 RECT 10.49 1.22 10.89 1.32 ;
 RECT 10.36 0.23 10.59 0.47 ;
 RECT 9.38 0.37 9.48 1.18 ;
 RECT 9.38 1.39 9.48 2.51 ;
 RECT 9.36 1.18 9.595 1.39 ;
 RECT 8.91 0.685 9.01 1.22 ;
 RECT 8.835 0.455 9.065 0.685 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.245 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 6.035 0.6 6.135 1.335 ;
 RECT 6.07 1.435 6.17 2.51 ;
 RECT 6.035 1.335 6.17 1.435 ;
 RECT 5.915 0.37 6.155 0.6 ;
 RECT 7.6 0.575 8.54 0.675 ;
 RECT 8.44 0.675 8.54 1.35 ;
 RECT 9.775 0.19 9.875 1.32 ;
 RECT 7.6 0.46 7.845 0.575 ;
 RECT 7.6 0.675 7.845 0.69 ;
 RECT 8.44 0.19 8.54 0.575 ;
 RECT 8.885 1.5 8.985 2.51 ;
 RECT 8.44 0.09 9.875 0.19 ;
 RECT 8.44 1.35 8.73 1.4 ;
 RECT 8.44 1.4 8.985 1.45 ;
 RECT 8.63 1.45 8.985 1.5 ;
 RECT 13.3 0.105 13.4 1.19 ;
 RECT 13.02 1.365 13.4 1.425 ;
 RECT 12.73 0.115 12.83 1.265 ;
 RECT 12.485 1.265 13.4 1.365 ;
 RECT 12.485 1.365 12.585 2.79 ;
 RECT 13.19 1.19 13.4 1.265 ;
 RECT 13.02 1.425 13.12 2.79 ;
 RECT 9.7 1.57 9.8 2.69 ;
 RECT 8.48 2.47 8.7 2.69 ;
 RECT 8.48 2.69 9.8 2.79 ;
 RECT 5.1 1.605 5.2 2.51 ;
 RECT 3.78 1.52 5.2 1.605 ;
 RECT 3.78 1.605 4.38 1.62 ;
 RECT 3.78 1.44 4.025 1.52 ;
 RECT 5.1 1.475 5.2 1.505 ;
 RECT 4.28 1.505 5.2 1.52 ;
 RECT 4.28 0.19 4.38 1.505 ;
 RECT 3.78 1.62 4.025 1.69 ;
 LAYER CO ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 13.24 1.8 13.37 1.93 ;
 RECT 13.24 2.06 13.37 2.19 ;
 RECT 10.54 2.17 10.67 2.3 ;
 RECT 7.255 1.45 7.385 1.58 ;
 RECT 5.645 1.32 5.775 1.45 ;
 RECT 7.59 0.885 7.72 1.015 ;
 RECT 7.585 2.015 7.715 2.145 ;
 RECT 3.93 0.21 4.06 0.34 ;
 RECT 7.315 2.64 7.445 2.77 ;
 RECT 7.93 0.915 8.06 1.045 ;
 RECT 8.53 2.525 8.66 2.655 ;
 RECT 8.635 1.815 8.765 1.945 ;
 RECT 13.23 1.24 13.36 1.37 ;
 RECT 13.52 0.68 13.65 0.81 ;
 RECT 12.95 0.77 13.08 0.9 ;
 RECT 9.41 1.22 9.54 1.35 ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 4.5 0.86 4.63 0.99 ;
 RECT 3.295 1.535 3.425 1.665 ;
 RECT 12.37 0.12 12.5 0.25 ;
 RECT 5.97 0.42 6.1 0.55 ;
 RECT 6.575 0.235 6.705 0.365 ;
 RECT 9.13 1.875 9.26 2.005 ;
 RECT 9.13 0.87 9.26 1 ;
 RECT 8.66 0.87 8.79 1 ;
 RECT 8.885 0.505 9.015 0.635 ;
 RECT 6.295 1.825 6.425 1.955 ;
 RECT 5.815 2.125 5.945 2.255 ;
 RECT 9.995 0.4 10.125 0.53 ;
 RECT 12.235 1.535 12.365 1.665 ;
 RECT 12.235 2.085 12.365 2.215 ;
 RECT 12.235 1.795 12.365 1.925 ;
 RECT 12.705 1.565 12.835 1.695 ;
 RECT 12.705 1.83 12.835 1.96 ;
 RECT 3.66 1.995 3.79 2.125 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 12.705 2.09 12.835 2.22 ;
 RECT 11.765 2.085 11.895 2.215 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 2.4 1.19 2.53 1.32 ;
 RECT 11.765 0.77 11.895 0.9 ;
 RECT 11.765 1.535 11.895 1.665 ;
 RECT 11.765 1.795 11.895 1.925 ;
 RECT 11.12 0.63 11.25 0.76 ;
 RECT 2.58 1.61 2.71 1.74 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 8.21 1.69 8.34 1.82 ;
 RECT 4.555 2.12 4.685 2.25 ;
 RECT 7.655 0.505 7.785 0.635 ;
 RECT 10.125 1.56 10.255 1.69 ;
 RECT 4.435 1.825 4.565 1.955 ;
 RECT 5.25 0.425 5.38 0.555 ;
 RECT 11.23 1.24 11.36 1.37 ;
 RECT 10.71 0.87 10.84 1 ;
 RECT 9.92 2.145 10.05 2.275 ;
 RECT 11.1 2.19 11.23 2.32 ;
 RECT 3.855 2.63 3.985 2.76 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.795 5.495 0.925 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.795 5.025 0.925 ;
 RECT 4.615 1.155 4.745 1.285 ;
 RECT 6.645 2.125 6.775 2.255 ;
 RECT 10.41 0.285 10.54 0.415 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 0.305 0.61 0.435 0.74 ;
 RECT 0.305 0.35 0.435 0.48 ;
 RECT 0.305 2.345 0.435 2.475 ;
 LAYER M1 ;
 RECT 5.745 2.12 6.845 2.26 ;
 RECT 5.18 0.42 5.825 0.56 ;
 RECT 5.685 0.56 5.825 0.79 ;
 RECT 7.18 0.5 7.855 0.64 ;
 RECT 7.18 0.64 7.32 0.79 ;
 RECT 5.685 0.79 7.32 0.93 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.365 2.11 2.995 2.25 ;
 RECT 4.89 0.67 5.03 2.035 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 3.46 0.53 5.03 0.67 ;
 RECT 4.845 2.035 5.03 2.17 ;
 RECT 4.845 2.17 4.985 2.305 ;
 RECT 9.405 1.24 9.545 1.41 ;
 RECT 11.395 0.58 11.535 0.955 ;
 RECT 10.705 0.955 11.535 1.095 ;
 RECT 10.705 1.095 10.845 1.1 ;
 RECT 10.705 1.24 10.845 1.395 ;
 RECT 9.405 1.1 10.845 1.24 ;
 RECT 10.705 0.815 10.845 0.955 ;
 RECT 10.535 1.535 10.675 2.35 ;
 RECT 10.535 1.395 10.845 1.535 ;
 RECT 13.225 0.58 13.365 1.45 ;
 RECT 11.395 0.44 13.365 0.58 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 8.14 1.685 8.795 1.81 ;
 RECT 8.655 1.005 8.795 1.685 ;
 RECT 8.14 1.81 8.835 1.825 ;
 RECT 8.565 1.825 8.835 1.95 ;
 RECT 8.585 0.865 8.865 1.005 ;
 RECT 6.305 1.07 7.72 1.21 ;
 RECT 7.52 0.875 8.13 1.05 ;
 RECT 7.52 1.05 7.72 1.07 ;
 RECT 7.58 1.21 7.72 2.215 ;
 RECT 6.305 1.21 6.445 1.315 ;
 RECT 5.575 1.315 6.445 1.455 ;
 RECT 4.495 1.075 4.75 1.365 ;
 RECT 4.495 1.365 4.69 1.82 ;
 RECT 4.495 0.81 4.635 1.075 ;
 RECT 4.365 1.82 4.69 1.96 ;
 RECT 4.545 1.96 4.69 2.3 ;
 RECT 9.125 1.695 9.335 1.87 ;
 RECT 9.125 0.805 9.265 1.555 ;
 RECT 9.055 1.87 9.335 2.01 ;
 RECT 10.815 1.92 10.955 2.52 ;
 RECT 10.25 2.52 10.955 2.66 ;
 RECT 9.125 1.555 10.39 1.695 ;
 RECT 10.25 1.695 10.39 2.52 ;
 RECT 11.05 1.375 11.19 1.78 ;
 RECT 11.05 1.235 11.43 1.375 ;
 RECT 10.815 1.78 11.19 1.92 ;
 RECT 5.185 1.82 7.39 1.96 ;
 RECT 5.185 1.005 5.5 1.145 ;
 RECT 5.36 0.705 5.5 1.005 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 7.25 1.38 7.39 1.82 ;
 RECT 5.185 1.145 5.325 1.82 ;
 RECT 3.635 1.775 3.84 1.99 ;
 RECT 3.7 1.63 3.84 1.775 ;
 RECT 3.7 1.475 4.045 1.63 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 4.18 2.48 4.32 2.51 ;
 RECT 3.635 2.34 4.32 2.48 ;
 RECT 3.59 1.99 3.84 2.13 ;
 RECT 3.635 2.13 3.775 2.34 ;
 RECT 4.18 2.51 7.125 2.65 ;
 RECT 6.985 2.495 7.125 2.51 ;
 RECT 7.86 1.21 8.44 1.35 ;
 RECT 8.46 2.24 8.6 2.52 ;
 RECT 7.86 1.35 8 2.1 ;
 RECT 7.86 2.24 8 2.355 ;
 RECT 7.86 2.1 8.6 2.24 ;
 RECT 6.985 2.355 8 2.495 ;
 RECT 8.58 0.5 9.09 0.58 ;
 RECT 8.3 0.58 9.09 0.64 ;
 RECT 8.3 0.64 8.76 0.72 ;
 RECT 8.3 0.72 8.44 1.21 ;
 RECT 8.46 2.52 8.715 2.66 ;
 END
END SDFFNARX2

MACRO SDFFNASRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 14.08 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 14.08 2.96 ;
 RECT 3.835 2.38 4.085 2.8 ;
 RECT 7.265 2.635 7.525 2.8 ;
 RECT 1.27 1.985 1.41 2.8 ;
 RECT 12.195 2.06 12.335 2.8 ;
 RECT 13.72 1.73 13.86 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 8.285 2.38 8.425 2.8 ;
 RECT 3.18 1.98 3.32 2.8 ;
 RECT 11.075 2.085 11.215 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 14.08 0.08 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 3.81 0.08 4.11 0.26 ;
 RECT 10.535 0.08 10.785 0.54 ;
 RECT 6.525 0.08 6.76 0.26 ;
 RECT 12.215 0.08 12.355 0.7 ;
 RECT 0.3 0.08 0.44 0.79 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 13.805 0.08 13.945 0.88 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.255 0.36 10.395 1.115 ;
 RECT 5.92 0.51 7.075 0.65 ;
 RECT 10.255 1.115 11.18 1.255 ;
 RECT 10.96 0.28 11.24 0.42 ;
 RECT 7.945 0.36 8.33 0.645 ;
 RECT 6.935 0.22 10.395 0.36 ;
 RECT 6.935 0.36 7.075 0.51 ;
 RECT 10.96 0.42 11.18 1.115 ;
 END
 ANTENNAGATEAREA 0.105 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.875 1.68 2.715 1.82 ;
 RECT 1.555 2.07 2.015 2.49 ;
 RECT 2.575 1.82 2.715 1.89 ;
 RECT 2.575 1.615 2.715 1.68 ;
 RECT 1.875 1.82 2.015 2.07 ;
 RECT 1.875 1.11 2.015 1.68 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.225 1.15 2.58 1.465 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.775 0.505 10.115 0.935 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.78 1.105 13.105 1.425 ;
 RECT 12.78 1.425 12.92 2.35 ;
 RECT 12.8 0.545 12.94 1.105 ;
 END
 ANTENNADIFFAREA 0.714 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.07 2.015 13.45 2.38 ;
 RECT 13.245 0.7 13.385 2.015 ;
 END
 ANTENNADIFFAREA 0.506 ;
 END Q

 OBS
 LAYER PO ;
 RECT 3.78 1.585 5.2 1.62 ;
 RECT 3.78 1.62 4.025 1.69 ;
 RECT 4.215 1.62 5.2 1.685 ;
 RECT 4.215 1.685 4.315 2.27 ;
 RECT 3.78 1.44 4.025 1.52 ;
 RECT 4.28 0.685 4.38 1.52 ;
 RECT 4.6 0.285 4.7 0.585 ;
 RECT 4.6 0.185 6.435 0.285 ;
 RECT 6.335 0.285 6.435 1.24 ;
 RECT 4.28 0.585 4.7 0.685 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 7.67 1.33 7.77 1.565 ;
 RECT 8.06 1.665 8.16 2.69 ;
 RECT 10.035 0.73 10.135 2.69 ;
 RECT 7.15 0.635 7.25 1.23 ;
 RECT 7.15 1.23 7.77 1.33 ;
 RECT 7.67 1.565 8.16 1.665 ;
 RECT 8.06 2.69 10.135 2.79 ;
 RECT 9.84 0.51 10.135 0.73 ;
 RECT 12.28 1.1 12.63 1.33 ;
 RECT 12.53 0.095 12.63 1.1 ;
 RECT 12.53 1.33 12.63 2.79 ;
 RECT 11.205 1.63 11.43 1.94 ;
 RECT 11.33 1.94 11.43 2.56 ;
 RECT 10.835 0.65 10.935 1.53 ;
 RECT 10.835 1.53 11.43 1.63 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 2.665 1.865 2.765 2.48 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 8.045 0.865 8.44 1.095 ;
 RECT 8.34 1.095 8.44 1.64 ;
 RECT 8.34 1.64 8.575 1.87 ;
 RECT 10.645 2.47 10.96 2.71 ;
 RECT 10.86 1.83 10.96 2.47 ;
 RECT 9.56 0.645 9.66 1.24 ;
 RECT 9.56 1.24 9.805 1.45 ;
 RECT 9.56 1.45 9.66 2.37 ;
 RECT 9.09 0.685 9.19 1.255 ;
 RECT 9.015 0.455 9.245 0.685 ;
 RECT 11.14 0.47 11.24 1.22 ;
 RECT 11.89 1.32 11.99 2.545 ;
 RECT 11.14 1.22 11.99 1.32 ;
 RECT 10.985 0.29 11.24 0.47 ;
 RECT 10.985 0.23 11.215 0.29 ;
 RECT 6.035 0.695 6.135 1.61 ;
 RECT 6.07 1.71 6.17 2.48 ;
 RECT 6.035 1.61 6.17 1.71 ;
 RECT 5.915 0.465 6.155 0.695 ;
 RECT 7.2 1.61 7.465 1.82 ;
 RECT 7.365 1.82 7.465 2.49 ;
 RECT 6.795 0.625 6.895 1.51 ;
 RECT 6.795 1.51 7.465 1.61 ;
 RECT 4.62 2.33 4.72 2.685 ;
 RECT 6.895 1.79 6.995 2.685 ;
 RECT 4.5 2.09 4.72 2.33 ;
 RECT 4.62 2.685 6.995 2.785 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.245 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 2.245 1.455 2.345 1.645 ;
 RECT 2.665 0.655 2.765 1.245 ;
 RECT 2.245 1.225 2.465 1.245 ;
 RECT 2.245 1.345 2.465 1.455 ;
 RECT 2.245 1.245 2.765 1.345 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.195 1.745 2.295 2.49 ;
 RECT 13.505 0.23 13.605 1.175 ;
 RECT 13.505 1.41 13.605 2.79 ;
 RECT 13.505 1.175 13.72 1.41 ;
 RECT 8.62 0.265 8.72 0.585 ;
 RECT 8.62 0.685 8.72 1.35 ;
 RECT 10.375 0.265 10.475 1.32 ;
 RECT 7.52 0.455 7.75 0.585 ;
 RECT 7.52 0.585 8.72 0.685 ;
 RECT 9.065 1.545 9.165 2.405 ;
 RECT 8.62 0.165 10.475 0.265 ;
 RECT 8.62 1.35 8.91 1.445 ;
 RECT 8.62 1.445 9.165 1.45 ;
 RECT 8.81 1.45 9.165 1.545 ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 5.595 1.33 5.735 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.635 0.65 5.735 1.33 ;
 RECT 5.595 1.475 5.825 1.71 ;
 RECT 5.145 0.705 5.245 1.21 ;
 RECT 4.575 1.16 4.82 1.21 ;
 RECT 4.575 1.21 5.245 1.31 ;
 RECT 4.575 1.31 4.82 1.405 ;
 RECT 5.145 0.47 5.43 0.705 ;
 RECT 5.1 1.685 5.2 2.495 ;
 RECT 3.78 1.52 4.38 1.585 ;
 LAYER CO ;
 RECT 13.25 1.91 13.38 2.04 ;
 RECT 13.25 2.17 13.38 2.3 ;
 RECT 13.725 2.32 13.855 2.45 ;
 RECT 13.25 0.75 13.38 0.88 ;
 RECT 12.33 1.15 12.46 1.28 ;
 RECT 13.725 1.8 13.855 1.93 ;
 RECT 13.725 2.06 13.855 2.19 ;
 RECT 11.035 0.285 11.165 0.415 ;
 RECT 12.805 0.615 12.935 0.745 ;
 RECT 12.785 1.65 12.915 1.78 ;
 RECT 12.785 1.91 12.915 2.04 ;
 RECT 9.31 1.9 9.44 2.03 ;
 RECT 9.31 0.87 9.44 1 ;
 RECT 10.26 1.92 10.39 2.05 ;
 RECT 9.78 1.965 9.91 2.095 ;
 RECT 8.84 0.87 8.97 1 ;
 RECT 9.065 0.505 9.195 0.635 ;
 RECT 9.62 1.28 9.75 1.41 ;
 RECT 11.08 2.17 11.21 2.3 ;
 RECT 10.61 2.135 10.74 2.265 ;
 RECT 8.115 0.915 8.245 1.045 ;
 RECT 11.64 2.13 11.77 2.26 ;
 RECT 11.255 1.76 11.385 1.89 ;
 RECT 5.97 0.515 6.1 0.645 ;
 RECT 6.575 0.12 6.705 0.25 ;
 RECT 7.57 0.505 7.7 0.635 ;
 RECT 6.295 1.825 6.425 1.955 ;
 RECT 5.815 2.105 5.945 2.235 ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 3.905 2.385 4.035 2.515 ;
 RECT 12.2 2.13 12.33 2.26 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 4.63 1.205 4.76 1.335 ;
 RECT 7.255 1.63 7.385 1.76 ;
 RECT 5.645 1.525 5.775 1.655 ;
 RECT 7.59 0.88 7.72 1.01 ;
 RECT 7.585 2.015 7.715 2.145 ;
 RECT 3.93 0.125 4.06 0.255 ;
 RECT 7.315 2.64 7.445 2.77 ;
 RECT 6.645 2.125 6.775 2.255 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 3.295 1.535 3.425 1.665 ;
 RECT 3.71 1.995 3.84 2.125 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 11.36 0.87 11.49 1 ;
 RECT 4.435 1.825 4.565 1.955 ;
 RECT 5.25 0.525 5.38 0.655 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 9.935 0.56 10.065 0.69 ;
 RECT 10.71 2.525 10.84 2.655 ;
 RECT 8.815 1.815 8.945 1.945 ;
 RECT 12.22 0.505 12.35 0.635 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 8.395 1.69 8.525 1.82 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 10.595 0.405 10.725 0.535 ;
 RECT 12.785 2.17 12.915 2.3 ;
 RECT 4.55 2.145 4.68 2.275 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 2.285 1.275 2.415 1.405 ;
 RECT 0.305 0.61 0.435 0.74 ;
 RECT 0.305 0.35 0.435 0.48 ;
 RECT 8.29 2.44 8.42 2.57 ;
 RECT 13.55 1.225 13.68 1.355 ;
 RECT 13.81 0.68 13.94 0.81 ;
 RECT 13.25 1.65 13.38 1.78 ;
 LAYER M1 ;
 RECT 5.745 2.1 6.845 2.26 ;
 RECT 5.18 0.52 5.78 0.66 ;
 RECT 5.64 0.66 5.78 0.79 ;
 RECT 7.215 0.5 7.795 0.64 ;
 RECT 5.64 0.79 7.355 0.93 ;
 RECT 7.215 0.64 7.355 0.79 ;
 RECT 7.52 0.875 8.315 1.05 ;
 RECT 6.97 1.185 7.72 1.325 ;
 RECT 7.52 1.05 7.72 1.185 ;
 RECT 7.58 1.325 7.72 2.01 ;
 RECT 5.575 1.52 7.11 1.66 ;
 RECT 6.97 1.325 7.11 1.52 ;
 RECT 7.53 2.01 7.785 2.15 ;
 RECT 9.615 1.395 11.775 1.535 ;
 RECT 11.635 1.535 11.775 2.33 ;
 RECT 11.635 1.105 11.775 1.395 ;
 RECT 11.355 0.76 11.495 0.855 ;
 RECT 11.355 0.995 11.775 1.105 ;
 RECT 9.615 1.21 9.755 1.395 ;
 RECT 11.355 0.855 12.64 0.995 ;
 RECT 12.5 0.36 12.64 0.855 ;
 RECT 12.5 0.22 13.665 0.36 ;
 RECT 13.525 0.36 13.665 1.175 ;
 RECT 13.525 1.175 13.72 1.455 ;
 RECT 4.365 1.82 4.685 1.96 ;
 RECT 4.495 1.385 4.685 1.82 ;
 RECT 4.545 1.96 4.685 2.345 ;
 RECT 4.495 0.84 4.685 1.155 ;
 RECT 4.495 1.155 4.765 1.385 ;
 RECT 7.925 1.35 8.065 2.1 ;
 RECT 7.925 2.24 8.065 2.295 ;
 RECT 6.985 2.295 8.065 2.435 ;
 RECT 4.225 2.515 7.125 2.655 ;
 RECT 6.985 2.435 7.125 2.515 ;
 RECT 3.705 1.475 4.045 2.1 ;
 RECT 4.225 2.24 4.365 2.515 ;
 RECT 3.775 0.825 4.045 1.475 ;
 RECT 3.705 2.1 4.365 2.24 ;
 RECT 9.425 2.32 9.565 2.52 ;
 RECT 7.925 2.18 9.495 2.185 ;
 RECT 7.925 2.185 9.565 2.24 ;
 RECT 8.48 0.5 9.27 0.64 ;
 RECT 8.78 2.24 9.565 2.32 ;
 RECT 7.925 2.1 8.92 2.18 ;
 RECT 8.48 0.64 8.62 1.21 ;
 RECT 7.925 1.21 8.62 1.35 ;
 RECT 9.425 2.52 10.92 2.66 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.27 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.365 2.11 2.995 2.25 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 3.46 0.53 4.41 0.67 ;
 RECT 4.27 0.22 5.03 0.36 ;
 RECT 4.89 0.36 5.03 0.875 ;
 RECT 4.845 2.035 5.045 2.305 ;
 RECT 4.905 1.015 5.045 2.035 ;
 RECT 4.27 0.36 4.41 0.53 ;
 RECT 4.825 0.875 5.1 1.015 ;
 RECT 5.185 1.82 7.39 1.96 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 5.36 0.805 5.5 1.22 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 7.25 1.56 7.39 1.82 ;
 RECT 5.185 1.36 5.325 1.82 ;
 RECT 9.775 2.1 9.96 2.22 ;
 RECT 10.605 2.065 10.745 2.22 ;
 RECT 9.73 1.96 9.96 2.1 ;
 RECT 9.775 2.22 10.745 2.36 ;
 RECT 8.765 0.865 9.045 1.685 ;
 RECT 8.765 1.825 9.045 1.95 ;
 RECT 8.325 1.685 9.045 1.825 ;
 RECT 9.305 1.675 11.495 1.815 ;
 RECT 11.915 1.92 12.055 2.505 ;
 RECT 11.195 1.815 11.495 1.935 ;
 RECT 11.355 1.935 11.495 2.505 ;
 RECT 11.355 2.505 12.055 2.645 ;
 RECT 9.305 0.805 9.445 1.675 ;
 RECT 9.305 1.815 9.515 1.895 ;
 RECT 9.235 1.895 9.515 2.035 ;
 RECT 10.21 1.815 10.44 2.055 ;
 RECT 12.15 1.285 12.29 1.78 ;
 RECT 12.15 1.145 12.53 1.285 ;
 RECT 11.915 1.78 12.29 1.92 ;
 END
END SDFFNASRX1

MACRO SDFFNASRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 14.72 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 14.72 2.96 ;
 RECT 7.265 2.635 7.525 2.8 ;
 RECT 3.75 2.7 4.025 2.8 ;
 RECT 14.195 1.485 14.335 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 3.18 1.93 3.32 2.8 ;
 RECT 13.25 1.485 13.39 2.8 ;
 RECT 1.27 1.985 1.41 2.8 ;
 RECT 8.285 2.38 8.425 2.8 ;
 RECT 11.075 2.21 11.215 2.8 ;
 RECT 12.195 2.06 12.335 2.8 ;
 RECT 3.755 2.635 4.025 2.7 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 14.72 0.08 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 3.88 0.08 4.11 0.39 ;
 RECT 10.545 0.08 10.8 0.845 ;
 RECT 6.525 0.08 6.76 0.37 ;
 RECT 13.38 0.08 13.615 0.46 ;
 RECT 12.215 0.08 12.355 0.74 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 14.475 0.08 14.615 0.86 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.935 0.22 9.745 0.36 ;
 RECT 5.92 0.51 7.075 0.65 ;
 RECT 10.195 1 11.485 1.14 ;
 RECT 6.935 0.36 7.075 0.51 ;
 RECT 9.395 0.36 9.745 0.635 ;
 RECT 9.605 0.635 9.745 0.83 ;
 RECT 9.605 0.83 10.335 0.97 ;
 RECT 10.195 0.97 10.335 1 ;
 END
 ANTENNAGATEAREA 0.172 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.202 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.615 2.04 2.015 2.415 ;
 RECT 2.575 1.51 2.715 1.72 ;
 RECT 1.875 1.72 2.715 1.86 ;
 RECT 1.875 1.86 2.015 2.04 ;
 RECT 1.875 1.11 2.015 1.72 ;
 END
 ANTENNAGATEAREA 0.101 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.2 0.96 2.715 1.37 ;
 END
 ANTENNAGATEAREA 0.101 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.885 0.31 10.285 0.685 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.78 1.44 12.92 2.575 ;
 RECT 12.78 1.105 13.09 1.44 ;
 RECT 12.78 0.5 12.92 1.105 ;
 END
 ANTENNADIFFAREA 0.544 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.72 2.015 14.05 2.4 ;
 RECT 13.72 0.6 14.21 0.74 ;
 RECT 13.72 2.4 13.86 2.58 ;
 RECT 13.72 0.74 13.86 2.015 ;
 END
 ANTENNADIFFAREA 0.568 ;
 END Q

 OBS
 LAYER PO ;
 RECT 9.56 1.24 9.805 1.45 ;
 RECT 9.56 1.45 9.66 2.51 ;
 RECT 9.09 0.685 9.19 1.19 ;
 RECT 9.015 0.455 9.245 0.685 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 2.965 0.405 3.065 2.79 ;
 RECT 12.28 1.17 13.135 1.2 ;
 RECT 12.53 0.12 12.63 1.1 ;
 RECT 12.53 1.1 13.135 1.17 ;
 RECT 12.28 1.2 12.63 1.4 ;
 RECT 13.035 0.1 13.135 1.1 ;
 RECT 13.035 1.2 13.135 2.775 ;
 RECT 12.53 1.4 12.63 2.775 ;
 RECT 13.505 1.3 13.605 2.775 ;
 RECT 13.345 1.2 13.605 1.3 ;
 RECT 13.79 0.35 13.89 1.1 ;
 RECT 14.26 0.35 14.36 1.1 ;
 RECT 13.345 1.1 14.36 1.2 ;
 RECT 13.345 1.065 13.6 1.1 ;
 RECT 13.98 1.2 14.08 2.775 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.79 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.79 ;
 RECT 8.06 1.515 8.16 2.69 ;
 RECT 10.035 0.685 10.135 2.69 ;
 RECT 7.15 0.635 7.25 1.13 ;
 RECT 7.15 1.13 7.77 1.23 ;
 RECT 7.67 1.23 7.77 1.415 ;
 RECT 7.67 1.415 8.16 1.515 ;
 RECT 8.06 2.69 10.135 2.79 ;
 RECT 9.965 0.475 10.195 0.685 ;
 RECT 10.645 2.47 10.96 2.71 ;
 RECT 10.86 1.635 10.96 2.47 ;
 RECT 11.33 1.79 11.43 2.79 ;
 RECT 10.87 0.65 10.97 1.355 ;
 RECT 11.205 1.455 11.43 1.79 ;
 RECT 10.87 1.355 11.43 1.455 ;
 RECT 8.045 0.835 8.44 1.065 ;
 RECT 8.34 1.065 8.44 1.415 ;
 RECT 8.34 1.415 8.575 1.645 ;
 RECT 11.325 0.495 11.425 0.935 ;
 RECT 11.89 1.175 11.99 2.79 ;
 RECT 11.255 0.935 11.485 1.075 ;
 RECT 11.255 1.075 11.99 1.175 ;
 RECT 6.035 0.695 6.135 1.445 ;
 RECT 6.07 1.545 6.17 2.495 ;
 RECT 6.035 1.445 6.17 1.545 ;
 RECT 5.915 0.465 6.155 0.695 ;
 RECT 7.2 1.51 7.465 1.64 ;
 RECT 7.365 1.64 7.465 2.52 ;
 RECT 6.795 0.625 6.895 1.41 ;
 RECT 6.795 1.41 7.465 1.51 ;
 RECT 5.635 0.65 5.735 1.295 ;
 RECT 5.595 1.53 5.695 2.495 ;
 RECT 5.595 1.295 5.825 1.53 ;
 RECT 2.47 1.11 2.765 1.24 ;
 RECT 2.665 0.655 2.765 1.11 ;
 RECT 2.195 1.71 2.295 2.79 ;
 RECT 2.245 1.34 2.345 1.61 ;
 RECT 2.195 1.61 2.345 1.71 ;
 RECT 2.245 1.24 2.765 1.34 ;
 RECT 4.465 2.09 4.71 2.675 ;
 RECT 6.895 1.735 6.995 2.675 ;
 RECT 4.465 2.675 6.995 2.775 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.255 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 4.28 0.285 4.38 1.44 ;
 RECT 4.185 1.69 4.285 2.28 ;
 RECT 5.1 1.5 5.2 1.545 ;
 RECT 5.1 1.645 5.2 2.495 ;
 RECT 6.335 0.285 6.435 1.24 ;
 RECT 4.28 0.185 6.435 0.285 ;
 RECT 3.78 1.44 4.38 1.545 ;
 RECT 3.78 1.645 4.38 1.69 ;
 RECT 3.78 1.545 5.2 1.645 ;
 RECT 8.62 0.635 8.72 1.125 ;
 RECT 10.375 0.265 10.475 1.22 ;
 RECT 8.62 0.265 8.72 0.535 ;
 RECT 7.645 0.46 7.875 0.535 ;
 RECT 7.645 0.535 8.72 0.635 ;
 RECT 7.645 0.635 7.875 0.69 ;
 RECT 9.065 1.5 9.165 2.51 ;
 RECT 8.62 0.165 10.475 0.265 ;
 RECT 8.62 1.125 8.91 1.225 ;
 RECT 8.81 1.225 8.91 1.4 ;
 RECT 8.81 1.4 9.165 1.5 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 2.665 1.76 2.765 2.79 ;
 RECT 2.525 1.52 2.765 1.76 ;
 RECT 4.56 1.15 5.245 1.31 ;
 RECT 5.145 0.705 5.245 1.15 ;
 RECT 4.56 1.31 4.805 1.365 ;
 RECT 5.145 0.47 5.43 0.705 ;
 RECT 9.56 0.645 9.66 1.24 ;
 LAYER CO ;
 RECT 3.305 1.535 3.435 1.665 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 1.995 3.315 2.125 ;
 RECT 10.71 2.525 10.84 2.655 ;
 RECT 8.815 1.815 8.945 1.945 ;
 RECT 8.29 2.44 8.42 2.57 ;
 RECT 14.48 0.68 14.61 0.81 ;
 RECT 13.385 1.115 13.515 1.245 ;
 RECT 14.01 0.605 14.14 0.735 ;
 RECT 12.33 1.22 12.46 1.35 ;
 RECT 12.785 0.55 12.915 0.68 ;
 RECT 12.785 1.825 12.915 1.955 ;
 RECT 12.785 2.085 12.915 2.215 ;
 RECT 12.22 0.54 12.35 0.67 ;
 RECT 2.58 1.56 2.71 1.69 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 8.395 1.465 8.525 1.595 ;
 RECT 8.115 0.885 8.245 1.015 ;
 RECT 11.305 1.005 11.435 1.135 ;
 RECT 10.62 0.695 10.75 0.825 ;
 RECT 5.97 0.515 6.1 0.645 ;
 RECT 6.575 0.23 6.705 0.36 ;
 RECT 7.695 0.51 7.825 0.64 ;
 RECT 14.2 1.555 14.33 1.685 ;
 RECT 9.78 2.02 9.91 2.15 ;
 RECT 8.84 0.805 8.97 0.935 ;
 RECT 9.065 0.505 9.195 0.635 ;
 RECT 13.725 1.555 13.855 1.685 ;
 RECT 13.725 2.35 13.855 2.48 ;
 RECT 13.725 1.825 13.855 1.955 ;
 RECT 11.64 0.715 11.77 0.845 ;
 RECT 11.08 2.28 11.21 2.41 ;
 RECT 10.61 2.19 10.74 2.32 ;
 RECT 12.785 1.555 12.915 1.685 ;
 RECT 12.785 2.35 12.915 2.48 ;
 RECT 7.255 1.45 7.385 1.58 ;
 RECT 6.295 1.825 6.425 1.955 ;
 RECT 5.815 2.105 5.945 2.235 ;
 RECT 7.585 2.015 7.715 2.145 ;
 RECT 3.93 0.255 4.06 0.385 ;
 RECT 3.825 2.64 3.955 2.77 ;
 RECT 6.645 2.105 6.775 2.235 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.615 1.195 4.745 1.325 ;
 RECT 3.66 1.995 3.79 2.125 ;
 RECT 9.31 1.85 9.44 1.98 ;
 RECT 9.31 0.845 9.44 0.975 ;
 RECT 10.26 1.92 10.39 2.05 ;
 RECT 5.25 0.525 5.38 0.655 ;
 RECT 9.62 1.28 9.75 1.41 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 2.53 1.165 2.66 1.295 ;
 RECT 12.2 2.13 12.33 2.26 ;
 RECT 11.64 2.13 11.77 2.26 ;
 RECT 11.255 1.61 11.385 1.74 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 5.645 1.345 5.775 1.475 ;
 RECT 7.59 0.88 7.72 1.01 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 7.315 2.64 7.445 2.77 ;
 RECT 10.015 0.515 10.145 0.645 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.58 2.35 0.71 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 4.52 2.15 4.65 2.28 ;
 RECT 13.43 0.325 13.56 0.455 ;
 RECT 13.255 1.555 13.385 1.685 ;
 RECT 13.255 2.35 13.385 2.48 ;
 RECT 13.255 1.825 13.385 1.955 ;
 RECT 13.255 2.085 13.385 2.215 ;
 RECT 4.5 1.835 4.63 1.965 ;
 RECT 14.2 2.35 14.33 2.48 ;
 RECT 14.2 1.825 14.33 1.955 ;
 RECT 14.2 2.085 14.33 2.215 ;
 RECT 13.725 2.085 13.855 2.215 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 4.5 0.905 4.63 1.035 ;
 LAYER M1 ;
 RECT 5.745 2.1 6.845 2.24 ;
 RECT 5.18 0.52 5.78 0.66 ;
 RECT 5.64 0.66 5.78 0.79 ;
 RECT 5.64 0.79 7.355 0.93 ;
 RECT 7.215 0.505 7.875 0.645 ;
 RECT 7.215 0.645 7.355 0.79 ;
 RECT 4.495 2.04 4.655 2.345 ;
 RECT 4.495 1.375 4.635 2.04 ;
 RECT 4.495 0.84 4.635 1.145 ;
 RECT 4.495 1.145 4.75 1.375 ;
 RECT 7.52 0.875 8.315 1.02 ;
 RECT 7.52 1.02 7.72 1.07 ;
 RECT 7.58 1.21 7.72 2.01 ;
 RECT 6.2 1.07 7.72 1.21 ;
 RECT 5.575 1.34 6.34 1.48 ;
 RECT 7.53 2.01 7.785 2.15 ;
 RECT 6.2 1.21 6.34 1.34 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 9.305 0.78 9.445 1.72 ;
 RECT 9.375 1.985 9.515 1.99 ;
 RECT 9.235 1.86 9.515 1.985 ;
 RECT 9.305 1.72 11.495 1.745 ;
 RECT 10.255 1.605 11.495 1.72 ;
 RECT 11.915 1.92 12.055 2.52 ;
 RECT 11.355 2.52 12.055 2.66 ;
 RECT 11.355 1.745 11.495 2.52 ;
 RECT 9.305 1.745 10.44 1.845 ;
 RECT 9.235 1.845 10.44 1.86 ;
 RECT 10.21 1.86 10.44 2.055 ;
 RECT 12.15 1.355 12.29 1.78 ;
 RECT 12.15 1.215 12.53 1.355 ;
 RECT 11.915 1.78 12.29 1.92 ;
 RECT 2.855 0.715 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.155 0.575 2.995 0.715 ;
 RECT 2.365 2.11 2.995 2.25 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 4.89 0.67 5.03 2.05 ;
 RECT 3.46 0.53 5.03 0.67 ;
 RECT 4.845 2.05 5.03 2.315 ;
 RECT 9.425 2.32 9.565 2.52 ;
 RECT 7.925 2.18 9.565 2.24 ;
 RECT 8.565 2.24 9.565 2.32 ;
 RECT 7.925 1.3 8.065 2.1 ;
 RECT 7.925 2.24 8.065 2.295 ;
 RECT 6.985 2.295 8.065 2.435 ;
 RECT 4.215 2.52 7.125 2.66 ;
 RECT 6.985 2.435 7.125 2.52 ;
 RECT 8.48 0.5 9.245 0.64 ;
 RECT 7.925 2.1 8.705 2.18 ;
 RECT 8.48 0.64 8.62 1.16 ;
 RECT 7.925 1.16 8.62 1.3 ;
 RECT 3.7 1.475 4.045 1.63 ;
 RECT 3.7 1.63 3.84 1.925 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.7 2.175 3.84 2.355 ;
 RECT 4.215 2.495 4.355 2.52 ;
 RECT 3.7 2.355 4.355 2.495 ;
 RECT 3.655 1.925 3.84 2.175 ;
 RECT 9.425 2.52 10.92 2.66 ;
 RECT 9.615 1.21 9.755 1.3 ;
 RECT 9.615 1.44 9.755 1.48 ;
 RECT 11.635 0.885 12.635 1.03 ;
 RECT 12.495 0.36 12.635 0.885 ;
 RECT 11.635 1.03 11.775 1.3 ;
 RECT 11.635 1.44 11.775 2.33 ;
 RECT 11.635 0.65 11.775 0.885 ;
 RECT 9.615 1.3 11.775 1.44 ;
 RECT 13.09 0.36 13.23 0.67 ;
 RECT 12.495 0.22 13.23 0.36 ;
 RECT 13.25 0.81 13.39 1.11 ;
 RECT 13.25 1.11 13.58 1.25 ;
 RECT 13.09 0.67 13.39 0.81 ;
 RECT 5.185 1.82 7.39 1.96 ;
 RECT 5.185 1.06 5.5 1.2 ;
 RECT 5.36 0.805 5.5 1.06 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 7.25 1.38 7.39 1.82 ;
 RECT 5.185 1.2 5.325 1.82 ;
 RECT 9.775 2.155 9.96 2.22 ;
 RECT 9.775 2 9.915 2.015 ;
 RECT 9.775 2.22 10.795 2.36 ;
 RECT 10.555 2.185 10.795 2.22 ;
 RECT 9.73 2.015 9.96 2.155 ;
 RECT 8.765 1.6 8.975 1.81 ;
 RECT 8.835 0.94 8.975 1.46 ;
 RECT 8.325 1.46 8.975 1.6 ;
 RECT 8.765 1.81 9.015 1.95 ;
 RECT 8.765 0.8 9.045 0.94 ;
 END
END SDFFNASRX2

MACRO SDFFNASX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 12.8 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 12.8 2.96 ;
 RECT 3.98 2.555 4.12 2.8 ;
 RECT 6.33 2.62 6.59 2.8 ;
 RECT 1.51 2.025 1.65 2.8 ;
 RECT 3.42 2 3.56 2.8 ;
 RECT 0.54 1.76 0.68 2.8 ;
 RECT 10.18 2.055 10.32 2.8 ;
 RECT 11.855 1.48 11.995 2.8 ;
 RECT 7.405 2.38 7.545 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 12.8 0.08 ;
 RECT 3.375 0.89 3.605 1.03 ;
 RECT 3.995 0.08 4.225 0.385 ;
 RECT 0.54 0.08 0.68 0.795 ;
 RECT 9.695 0.08 9.835 1.07 ;
 RECT 1.51 0.08 1.65 1.075 ;
 RECT 11.95 0.08 12.09 0.76 ;
 RECT 6.385 0.08 6.525 0.38 ;
 RECT 3.42 0.08 3.56 0.89 ;
 END
 END VSS

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.8 0.325 9.24 0.66 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.19 0.52 11.525 0.815 ;
 RECT 11.3 0.815 11.44 2.51 ;
 END
 ANTENNADIFFAREA 0.553 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.145 2.065 12.475 2.385 ;
 RECT 12.335 0.85 12.56 0.99 ;
 RECT 12.42 0.535 12.56 0.85 ;
 RECT 12.335 2.385 12.475 2.52 ;
 RECT 12.335 0.99 12.475 2.065 ;
 END
 ANTENNADIFFAREA 0.46 ;
 END Q

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.445 1.495 1.925 1.77 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.9 2.125 2.255 2.385 ;
 RECT 2.115 1.13 2.255 2.125 ;
 RECT 2.815 2.625 2.955 2.66 ;
 RECT 2.115 2.455 2.955 2.625 ;
 RECT 2.815 2.41 2.955 2.455 ;
 RECT 2.115 2.385 2.255 2.455 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.525 1.245 2.86 1.605 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.485 1.48 3.885 1.805 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 OBS
 LAYER PO ;
 RECT 4.455 1.255 4.62 1.355 ;
 RECT 7.075 0.575 7.825 0.675 ;
 RECT 7.725 0.675 7.825 1.35 ;
 RECT 9.48 0.19 9.58 1.175 ;
 RECT 7.725 0.19 7.825 0.575 ;
 RECT 7.075 0.455 7.305 0.575 ;
 RECT 7.075 0.675 7.305 0.685 ;
 RECT 8.17 1.545 8.27 2.51 ;
 RECT 7.725 0.09 9.58 0.19 ;
 RECT 7.725 1.35 8.015 1.445 ;
 RECT 7.725 1.445 8.27 1.45 ;
 RECT 7.915 1.45 8.27 1.545 ;
 RECT 7.445 1.095 7.545 1.64 ;
 RECT 7.445 1.64 7.76 1.87 ;
 RECT 7.275 0.865 7.545 1.095 ;
 RECT 12.205 0.215 12.305 1.035 ;
 RECT 12.115 1.27 12.215 2.79 ;
 RECT 11.955 1.035 12.305 1.27 ;
 RECT 10.435 1.285 10.535 1.72 ;
 RECT 10.31 1.17 10.535 1.285 ;
 RECT 10.435 1.94 10.535 2.75 ;
 RECT 9.95 0.6 10.05 1.07 ;
 RECT 9.95 1.07 10.535 1.17 ;
 RECT 10.345 1.72 10.575 1.94 ;
 RECT 5.385 0.705 5.485 1.255 ;
 RECT 5.385 0.47 5.67 0.705 ;
 RECT 4.8 1.19 5.045 1.255 ;
 RECT 4.8 1.355 5.045 1.44 ;
 RECT 4.8 1.255 5.485 1.355 ;
 RECT 1.295 1.495 1.865 1.77 ;
 RECT 1.765 0.675 1.865 1.495 ;
 RECT 1.765 1.77 1.865 2.485 ;
 RECT 1.295 0.655 1.395 1.495 ;
 RECT 1.295 1.77 1.395 2.485 ;
 RECT 2.1 0.66 2.2 1.165 ;
 RECT 2.06 1.165 2.305 1.405 ;
 RECT 3 0.195 3.305 0.425 ;
 RECT 3.205 0.425 3.305 2.485 ;
 RECT 8.665 0.6 8.765 1.24 ;
 RECT 8.665 1.24 8.91 1.45 ;
 RECT 8.665 1.45 8.765 2.505 ;
 RECT 8.195 0.6 8.295 1.175 ;
 RECT 8.12 0.37 8.35 0.6 ;
 RECT 6.495 0.625 6.595 1.58 ;
 RECT 6.625 1.82 6.725 2.69 ;
 RECT 6.495 1.58 6.735 1.82 ;
 RECT 5.835 1.43 5.935 1.475 ;
 RECT 5.835 1.71 5.935 2.505 ;
 RECT 5.855 0.65 5.955 1.33 ;
 RECT 5.835 1.33 5.955 1.43 ;
 RECT 5.705 1.475 5.935 1.71 ;
 RECT 6.14 1.795 6.24 2.685 ;
 RECT 4.735 2.11 4.965 2.685 ;
 RECT 4.735 2.685 6.24 2.785 ;
 RECT 3.68 0.675 3.78 1.5 ;
 RECT 3.485 1.5 3.78 1.74 ;
 RECT 3.68 1.74 3.78 2.39 ;
 RECT 2.905 1.655 3.005 2.43 ;
 RECT 2.765 2.43 3.005 2.66 ;
 RECT 10.985 1.28 11.195 1.415 ;
 RECT 10.985 1.18 11.665 1.28 ;
 RECT 11.565 0.145 11.665 1.18 ;
 RECT 11.565 1.28 11.665 2.79 ;
 RECT 2.485 1.475 2.585 1.665 ;
 RECT 2.905 0.675 3.005 1.245 ;
 RECT 2.435 1.765 2.535 2.49 ;
 RECT 2.435 1.665 2.585 1.765 ;
 RECT 2.485 1.245 3.005 1.475 ;
 RECT 9.965 1.505 10.065 2.545 ;
 RECT 9.42 2.47 9.67 2.545 ;
 RECT 9.42 2.645 9.67 2.71 ;
 RECT 9.42 2.545 10.065 2.645 ;
 RECT 7.115 1.375 7.215 2.69 ;
 RECT 6.795 1.275 7.215 1.375 ;
 RECT 7.115 2.69 9.24 2.79 ;
 RECT 9.14 0.655 9.24 2.69 ;
 RECT 6.795 0.635 6.895 1.275 ;
 RECT 8.965 0.435 9.24 0.655 ;
 RECT 4.205 1.44 4.555 1.635 ;
 RECT 4.455 1.355 4.555 1.44 ;
 RECT 4.205 1.635 5.44 1.69 ;
 RECT 4.455 1.735 4.555 2.31 ;
 RECT 4.455 1.69 5.44 1.735 ;
 RECT 6.17 0.285 6.27 1.24 ;
 RECT 4.52 0.185 6.27 0.285 ;
 RECT 4.52 0.285 4.62 1.255 ;
 RECT 5.34 1.735 5.44 2.495 ;
 LAYER CO ;
 RECT 9.365 1.965 9.495 2.095 ;
 RECT 8.885 1.965 9.015 2.095 ;
 RECT 7.945 0.82 8.075 0.95 ;
 RECT 8.17 0.415 8.3 0.545 ;
 RECT 7.92 1.815 8.05 1.945 ;
 RECT 7.41 2.44 7.54 2.57 ;
 RECT 11.995 1.085 12.125 1.215 ;
 RECT 10.395 1.76 10.525 1.89 ;
 RECT 6.565 1.63 6.695 1.76 ;
 RECT 5.755 1.525 5.885 1.655 ;
 RECT 6.85 2.015 6.98 2.145 ;
 RECT 4.045 0.25 4.175 0.38 ;
 RECT 7.34 0.915 7.47 1.045 ;
 RECT 7.125 0.505 7.255 0.635 ;
 RECT 4.785 2.15 4.915 2.28 ;
 RECT 0.545 0.61 0.675 0.74 ;
 RECT 2.12 1.215 2.25 1.345 ;
 RECT 0.545 0.35 0.675 0.48 ;
 RECT 3.425 0.895 3.555 1.025 ;
 RECT 11.025 1.23 11.155 1.36 ;
 RECT 12.34 1.53 12.47 1.66 ;
 RECT 12.34 1.79 12.47 1.92 ;
 RECT 12.34 2.05 12.47 2.18 ;
 RECT 12.34 2.31 12.47 2.44 ;
 RECT 11.86 1.53 11.99 1.66 ;
 RECT 2.655 2.135 2.785 2.265 ;
 RECT 2.64 1.295 2.77 1.425 ;
 RECT 0.545 2.365 0.675 2.495 ;
 RECT 3.9 2.015 4.03 2.145 ;
 RECT 1.515 0.895 1.645 1.025 ;
 RECT 4.87 1.245 5 1.375 ;
 RECT 1.515 2.075 1.645 2.205 ;
 RECT 1.52 1.57 1.65 1.7 ;
 RECT 2.82 2.48 2.95 2.61 ;
 RECT 3.425 2.07 3.555 2.2 ;
 RECT 4.275 1.495 4.405 1.625 ;
 RECT 5.135 0.88 5.265 1.01 ;
 RECT 0.545 2.105 0.675 2.235 ;
 RECT 4.03 0.895 4.16 1.025 ;
 RECT 6.39 0.2 6.52 0.33 ;
 RECT 4.675 1.86 4.805 1.99 ;
 RECT 5.49 0.525 5.62 0.655 ;
 RECT 9.485 2.525 9.615 2.655 ;
 RECT 4.74 0.905 4.87 1.035 ;
 RECT 11.305 0.585 11.435 0.715 ;
 RECT 7.015 0.88 7.145 1.01 ;
 RECT 11.305 1.53 11.435 1.66 ;
 RECT 9.025 0.485 9.155 0.615 ;
 RECT 11.955 0.56 12.085 0.69 ;
 RECT 7.58 1.69 7.71 1.82 ;
 RECT 8.415 1.9 8.545 2.03 ;
 RECT 8.415 0.82 8.545 0.95 ;
 RECT 9.7 0.82 9.83 0.95 ;
 RECT 8.725 1.28 8.855 1.41 ;
 RECT 10.17 0.82 10.3 0.95 ;
 RECT 10.185 2.115 10.315 2.245 ;
 RECT 9.715 2.11 9.845 2.24 ;
 RECT 11.305 1.79 11.435 1.92 ;
 RECT 10.745 2.13 10.875 2.26 ;
 RECT 11.86 1.79 11.99 1.92 ;
 RECT 11.86 2.05 11.99 2.18 ;
 RECT 11.86 2.31 11.99 2.44 ;
 RECT 11.305 2.05 11.435 2.18 ;
 RECT 11.305 2.31 11.435 2.44 ;
 RECT 6.38 2.64 6.51 2.77 ;
 RECT 12.425 0.605 12.555 0.735 ;
 RECT 1.045 2.075 1.175 2.205 ;
 RECT 1.045 0.895 1.175 1.025 ;
 RECT 0.545 1.845 0.675 1.975 ;
 RECT 3.05 0.245 3.18 0.375 ;
 RECT 3.535 1.555 3.665 1.685 ;
 RECT 2.46 0.895 2.59 1.025 ;
 RECT 3.985 2.64 4.115 2.77 ;
 RECT 5.585 2.07 5.715 2.2 ;
 RECT 5.605 0.88 5.735 1.01 ;
 RECT 5.09 2.105 5.22 2.235 ;
 LAYER M1 ;
 RECT 7.125 1.36 7.265 2.1 ;
 RECT 7.125 2.24 7.265 2.34 ;
 RECT 6.05 2.34 7.265 2.48 ;
 RECT 4.27 2.15 4.41 2.52 ;
 RECT 4.27 2.52 6.19 2.66 ;
 RECT 4.025 0.845 4.165 1.125 ;
 RECT 6.05 2.48 6.19 2.52 ;
 RECT 4.025 1.125 4.41 1.265 ;
 RECT 4.27 1.265 4.41 2.01 ;
 RECT 3.83 2.01 4.41 2.15 ;
 RECT 7.66 0.415 8.375 0.55 ;
 RECT 7.66 0.55 8.12 0.555 ;
 RECT 7.87 0.41 8.375 0.415 ;
 RECT 8.53 2.32 8.67 2.52 ;
 RECT 7.66 0.555 7.8 1.22 ;
 RECT 7.125 2.1 8.025 2.18 ;
 RECT 7.125 2.18 8.67 2.24 ;
 RECT 7.885 2.24 8.67 2.32 ;
 RECT 7.125 1.22 7.8 1.36 ;
 RECT 8.53 2.52 9.685 2.66 ;
 RECT 5.425 1.805 6.7 1.945 ;
 RECT 5.425 1.945 5.79 1.96 ;
 RECT 5.425 1.22 5.74 1.36 ;
 RECT 5.6 0.805 5.74 1.22 ;
 RECT 5.51 1.96 5.79 2.215 ;
 RECT 5.425 1.36 5.565 1.805 ;
 RECT 6.56 1.56 6.7 1.805 ;
 RECT 1.825 0.38 1.965 1.215 ;
 RECT 1.04 1.215 1.965 1.355 ;
 RECT 1.04 0.82 1.18 1.215 ;
 RECT 1.04 1.355 1.18 2.325 ;
 RECT 1.825 0.24 3.25 0.38 ;
 RECT 8.88 2.1 9.065 2.24 ;
 RECT 9.71 2.03 9.85 2.24 ;
 RECT 8.835 1.96 9.065 2.1 ;
 RECT 8.88 2.24 9.85 2.38 ;
 RECT 6.845 1.04 7.52 1.05 ;
 RECT 6.28 0.91 7.52 1.04 ;
 RECT 6.28 0.9 7.15 0.91 ;
 RECT 6.845 1.08 6.985 2.2 ;
 RECT 6.845 1.05 7.15 1.08 ;
 RECT 5.705 1.52 6.42 1.66 ;
 RECT 7.01 0.81 7.15 0.9 ;
 RECT 6.28 1.04 6.42 1.52 ;
 RECT 5.42 0.52 7.33 0.66 ;
 RECT 7.045 0.47 7.33 0.52 ;
 RECT 8.41 1.815 8.62 1.895 ;
 RECT 8.41 0.77 8.55 1.675 ;
 RECT 9.315 1.815 9.545 2.1 ;
 RECT 8.34 1.895 8.62 2.035 ;
 RECT 8.41 1.675 10.6 1.815 ;
 RECT 11.02 1.18 11.16 2.505 ;
 RECT 10.3 1.815 10.6 1.915 ;
 RECT 10.46 1.915 10.6 2.505 ;
 RECT 10.46 2.505 11.16 2.645 ;
 RECT 7.57 1.685 8.08 1.81 ;
 RECT 7.57 1.81 8.12 1.825 ;
 RECT 7.94 0.77 8.08 1.685 ;
 RECT 7.57 1.615 7.71 1.685 ;
 RECT 7.57 1.825 7.71 1.895 ;
 RECT 7.85 1.825 8.12 1.95 ;
 RECT 3.095 1.03 3.235 1.17 ;
 RECT 3.095 1.31 3.235 2.13 ;
 RECT 2.395 0.89 3.235 1.03 ;
 RECT 2.585 2.13 3.235 2.27 ;
 RECT 5.13 0.665 5.27 0.875 ;
 RECT 3.095 1.17 3.885 1.31 ;
 RECT 3.745 0.69 3.885 1.17 ;
 RECT 3.7 0.665 3.885 0.69 ;
 RECT 3.7 0.525 5.27 0.665 ;
 RECT 5.145 1.015 5.285 2.035 ;
 RECT 5.085 0.875 5.34 1.015 ;
 RECT 5.085 2.035 5.285 2.305 ;
 RECT 4.67 1.995 4.92 2.355 ;
 RECT 4.6 1.98 4.92 1.995 ;
 RECT 4.6 1.855 4.875 1.98 ;
 RECT 4.735 0.815 4.875 1.155 ;
 RECT 4.735 1.155 5.005 1.475 ;
 RECT 4.735 1.475 4.875 1.855 ;
 RECT 10.74 0.38 10.88 0.815 ;
 RECT 10.12 0.815 10.88 0.955 ;
 RECT 10.74 0.955 10.88 1.395 ;
 RECT 8.72 1.395 10.88 1.535 ;
 RECT 10.74 1.535 10.88 2.32 ;
 RECT 8.72 1.21 8.86 1.395 ;
 RECT 11.67 0.38 11.81 1.15 ;
 RECT 10.74 0.24 11.81 0.38 ;
 RECT 11.99 1.02 12.13 1.15 ;
 RECT 11.67 1.15 12.13 1.29 ;
 END
END SDFFNASX1

MACRO SDFFNASX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 13.76 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 13.76 2.96 ;
 RECT 1.51 2.025 1.65 2.8 ;
 RECT 3.975 2.62 4.275 2.8 ;
 RECT 6.395 2.635 6.675 2.8 ;
 RECT 3.42 2 3.56 2.8 ;
 RECT 0.54 1.76 0.68 2.8 ;
 RECT 10.18 1.99 10.32 2.8 ;
 RECT 11.305 1.48 11.445 2.8 ;
 RECT 7.405 2.38 7.545 2.8 ;
 RECT 12.25 1.48 12.39 2.8 ;
 RECT 13.22 1.435 13.36 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 13.76 0.08 ;
 RECT 1.465 0.89 1.695 1.03 ;
 RECT 3.995 0.08 4.225 0.385 ;
 RECT 3.42 0.08 3.56 0.52 ;
 RECT 11.185 0.08 11.455 0.245 ;
 RECT 12.2 0.08 12.47 0.245 ;
 RECT 6.385 0.08 6.525 0.38 ;
 RECT 0.54 0.08 0.68 0.795 ;
 RECT 9.695 0.08 9.835 1.07 ;
 RECT 13.215 0.08 13.355 0.825 ;
 RECT 1.51 0.08 1.65 0.89 ;
 END
 END VSS

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.72 2.255 8.145 2.66 ;
 END
 ANTENNAGATEAREA 0.2115 ;
 END SETB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.43 1.48 1.925 1.77 ;
 END
 ANTENNAGATEAREA 0.172 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.9 2.12 2.255 2.385 ;
 RECT 2.815 1.655 2.955 1.74 ;
 RECT 2.115 1.74 2.955 1.91 ;
 RECT 2.115 1.91 2.255 2.12 ;
 RECT 2.115 1.13 2.255 1.74 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.405 1.435 2.68 1.56 ;
 RECT 2.405 1.175 2.88 1.435 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END D

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.52 1.43 3.885 1.805 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.675 2.08 11.995 2.375 ;
 RECT 11.78 2.375 11.92 2.51 ;
 RECT 11.78 0.665 11.92 2.08 ;
 END
 ANTENNADIFFAREA 0.506 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.65 1.765 12.955 2.06 ;
 RECT 12.745 2.06 12.885 2.145 ;
 RECT 12.745 0.595 12.885 1.765 ;
 END
 ANTENNADIFFAREA 0.448 ;
 END Q

 OBS
 LAYER PO ;
 RECT 9.48 0.19 9.58 1.32 ;
 RECT 7.075 0.265 7.305 0.385 ;
 RECT 7.075 0.485 7.305 0.495 ;
 RECT 7.725 1.28 8.27 1.38 ;
 RECT 7.725 0.09 9.58 0.19 ;
 RECT 12.415 1.1 12.63 1.18 ;
 RECT 12.53 0.145 12.63 1.1 ;
 RECT 12.53 1.335 12.63 2.335 ;
 RECT 12.415 1.28 12.63 1.335 ;
 RECT 12.415 1.18 13.1 1.28 ;
 RECT 13 0.145 13.1 1.18 ;
 RECT 13 1.28 13.1 2.335 ;
 RECT 8.665 0.475 8.765 1.24 ;
 RECT 8.665 1.24 8.91 1.45 ;
 RECT 8.665 1.45 8.765 2.465 ;
 RECT 8.195 0.62 8.295 1.1 ;
 RECT 8.12 0.39 8.35 0.62 ;
 RECT 11.565 0.445 11.665 1.145 ;
 RECT 11.565 1.245 11.665 2.79 ;
 RECT 10.985 1.095 11.195 1.145 ;
 RECT 10.985 1.145 12.135 1.245 ;
 RECT 10.985 1.245 11.195 1.33 ;
 RECT 12.035 0.45 12.135 1.145 ;
 RECT 12.035 1.245 12.135 2.79 ;
 RECT 6.14 1.425 6.24 2.685 ;
 RECT 4.735 2.06 4.965 2.685 ;
 RECT 4.735 2.685 6.24 2.785 ;
 RECT 4.8 1.155 5.485 1.355 ;
 RECT 5.385 0.61 5.485 1.155 ;
 RECT 5.385 0.375 5.65 0.61 ;
 RECT 4.8 1.355 5.045 1.375 ;
 RECT 4.8 1.125 5.045 1.155 ;
 RECT 10.31 1.24 10.535 1.77 ;
 RECT 10.435 1.77 10.535 2.79 ;
 RECT 9.95 1.14 10.535 1.24 ;
 RECT 9.95 0.65 10.05 1.14 ;
 RECT 7.445 0.905 7.545 1.56 ;
 RECT 7.445 1.56 7.76 1.79 ;
 RECT 7.275 0.675 7.545 0.905 ;
 RECT 6.425 1.365 6.73 1.56 ;
 RECT 6.495 0.515 6.595 1.32 ;
 RECT 6.425 1.32 6.64 1.365 ;
 RECT 6.625 1.56 6.725 2.46 ;
 RECT 5.835 1.33 5.955 1.355 ;
 RECT 5.835 1.59 5.935 2.5 ;
 RECT 5.855 0.625 5.955 1.33 ;
 RECT 5.725 1.355 5.955 1.59 ;
 RECT 3.68 0.675 3.78 1.5 ;
 RECT 3.485 1.5 3.78 1.74 ;
 RECT 3.68 1.74 3.78 2.39 ;
 RECT 2.905 1.885 3.005 2.79 ;
 RECT 2.765 1.655 3.005 1.885 ;
 RECT 2.905 0.675 3.005 1.2 ;
 RECT 2.485 1.43 2.585 1.665 ;
 RECT 2.435 1.765 2.535 2.79 ;
 RECT 2.435 1.665 2.585 1.765 ;
 RECT 2.485 1.2 3.005 1.43 ;
 RECT 2.1 0.66 2.2 1.165 ;
 RECT 2.06 1.165 2.305 1.405 ;
 RECT 4.205 1.555 5.44 1.655 ;
 RECT 4.205 1.44 4.555 1.555 ;
 RECT 4.455 1.355 4.555 1.44 ;
 RECT 4.205 1.655 4.555 1.69 ;
 RECT 4.455 1.69 4.555 2.215 ;
 RECT 6.17 0.19 6.27 1.2 ;
 RECT 4.52 0.09 6.27 0.19 ;
 RECT 4.52 0.19 4.62 1.255 ;
 RECT 5.34 1.655 5.44 2.505 ;
 RECT 4.455 1.255 4.62 1.355 ;
 RECT 7.115 1.185 7.215 2.69 ;
 RECT 7.735 2.46 7.965 2.69 ;
 RECT 9.14 0.37 9.24 2.69 ;
 RECT 7.115 2.69 9.24 2.79 ;
 RECT 6.795 0.51 6.895 1.085 ;
 RECT 6.795 1.085 7.215 1.185 ;
 RECT 3.205 0.425 3.305 2.79 ;
 RECT 3 0.195 3.305 0.425 ;
 RECT 1.295 1.495 1.865 1.77 ;
 RECT 1.295 0.655 1.395 1.495 ;
 RECT 1.295 1.77 1.395 2.78 ;
 RECT 1.765 0.675 1.865 1.495 ;
 RECT 1.765 1.77 1.865 2.66 ;
 RECT 9.75 2.375 10.065 2.615 ;
 RECT 9.965 1.42 10.065 2.375 ;
 RECT 7.725 0.19 7.825 0.385 ;
 RECT 7.075 0.385 7.825 0.485 ;
 RECT 7.725 0.485 7.825 1.28 ;
 RECT 8.17 1.38 8.27 2.405 ;
 LAYER CO ;
 RECT 7.945 0.75 8.075 0.88 ;
 RECT 8.17 0.45 8.3 0.58 ;
 RECT 10.745 2.01 10.875 2.14 ;
 RECT 10.36 1.555 10.49 1.685 ;
 RECT 6.47 1.37 6.6 1.5 ;
 RECT 13.22 0.625 13.35 0.755 ;
 RECT 13.225 1.53 13.355 1.66 ;
 RECT 13.225 1.79 13.355 1.92 ;
 RECT 12.75 1.79 12.88 1.92 ;
 RECT 12.75 1.53 12.88 1.66 ;
 RECT 12.75 0.645 12.88 0.775 ;
 RECT 12.28 0.11 12.41 0.24 ;
 RECT 4.87 1.195 5 1.325 ;
 RECT 1.045 2.075 1.175 2.205 ;
 RECT 11.785 1.53 11.915 1.66 ;
 RECT 11.785 2.05 11.915 2.18 ;
 RECT 9.7 0.87 9.83 1 ;
 RECT 3.05 0.245 3.18 0.375 ;
 RECT 3.535 1.555 3.665 1.685 ;
 RECT 2.46 0.895 2.59 1.025 ;
 RECT 11.31 1.53 11.44 1.66 ;
 RECT 11.31 1.79 11.44 1.92 ;
 RECT 11.31 2.05 11.44 2.18 ;
 RECT 11.31 2.31 11.44 2.44 ;
 RECT 0.545 2.365 0.675 2.495 ;
 RECT 3.9 2.015 4.03 2.145 ;
 RECT 1.515 0.895 1.645 1.025 ;
 RECT 0.545 0.61 0.675 0.74 ;
 RECT 2.12 1.215 2.25 1.345 ;
 RECT 0.545 0.35 0.675 0.48 ;
 RECT 3.425 0.32 3.555 0.45 ;
 RECT 1.045 0.895 1.175 1.025 ;
 RECT 2.655 2.135 2.785 2.265 ;
 RECT 2.64 1.25 2.77 1.38 ;
 RECT 3.425 2.07 3.555 2.2 ;
 RECT 4.275 1.495 4.405 1.625 ;
 RECT 4.06 2.625 4.19 2.755 ;
 RECT 0.545 2.105 0.675 2.235 ;
 RECT 4.03 0.895 4.16 1.025 ;
 RECT 0.545 1.845 0.675 1.975 ;
 RECT 1.515 2.075 1.645 2.205 ;
 RECT 1.52 1.57 1.65 1.7 ;
 RECT 2.82 1.705 2.95 1.835 ;
 RECT 5.585 2.07 5.715 2.2 ;
 RECT 5.605 0.85 5.735 0.98 ;
 RECT 5.09 2.105 5.22 2.235 ;
 RECT 5.135 0.85 5.265 0.98 ;
 RECT 4.74 0.905 4.87 1.035 ;
 RECT 7.015 0.82 7.145 0.95 ;
 RECT 6.39 0.2 6.52 0.33 ;
 RECT 7.785 2.505 7.915 2.635 ;
 RECT 9.815 2.43 9.945 2.56 ;
 RECT 7.92 1.68 8.05 1.81 ;
 RECT 7.34 0.725 7.47 0.855 ;
 RECT 7.125 0.315 7.255 0.445 ;
 RECT 8.415 1.68 8.545 1.81 ;
 RECT 8.415 0.75 8.545 0.88 ;
 RECT 9.365 1.69 9.495 1.82 ;
 RECT 8.725 1.28 8.855 1.41 ;
 RECT 10.17 0.87 10.3 1 ;
 RECT 10.185 2.085 10.315 2.215 ;
 RECT 9.715 1.98 9.845 2.11 ;
 RECT 5.775 1.405 5.905 1.535 ;
 RECT 6.85 2.015 6.98 2.145 ;
 RECT 4.045 0.25 4.175 0.38 ;
 RECT 6.465 2.64 6.595 2.77 ;
 RECT 12.255 1.53 12.385 1.66 ;
 RECT 12.255 1.79 12.385 1.92 ;
 RECT 11.255 0.11 11.385 0.24 ;
 RECT 11.785 0.715 11.915 0.845 ;
 RECT 11.785 2.31 11.915 2.44 ;
 RECT 11.785 1.79 11.915 1.92 ;
 RECT 4.79 2.115 4.92 2.245 ;
 RECT 12.455 1.15 12.585 1.28 ;
 RECT 11.025 1.145 11.155 1.275 ;
 RECT 4.675 1.805 4.805 1.935 ;
 RECT 5.47 0.43 5.6 0.56 ;
 RECT 7.41 2.44 7.54 2.57 ;
 RECT 7.58 1.615 7.71 1.745 ;
 RECT 8.885 1.98 9.015 2.11 ;
 LAYER M1 ;
 RECT 8.81 1.975 9.915 2.115 ;
 RECT 10.74 0.745 11.63 0.865 ;
 RECT 10.12 0.865 11.63 0.885 ;
 RECT 11.49 0.525 11.63 0.745 ;
 RECT 11.49 0.885 11.63 0.89 ;
 RECT 10.12 0.885 10.88 1.005 ;
 RECT 10.74 1.005 10.88 1.22 ;
 RECT 8.72 1.22 10.88 1.36 ;
 RECT 10.74 1.36 10.88 2.2 ;
 RECT 8.72 1.21 8.86 1.22 ;
 RECT 8.72 1.36 8.86 1.48 ;
 RECT 11.49 0.385 12.59 0.525 ;
 RECT 12.45 0.525 12.59 1.34 ;
 RECT 7.94 0.885 8.08 1.535 ;
 RECT 7.575 1.675 7.715 1.825 ;
 RECT 7.895 0.745 8.145 0.885 ;
 RECT 7.515 1.535 8.15 1.675 ;
 RECT 7.865 1.675 8.15 1.815 ;
 RECT 5.425 1.805 6.605 1.945 ;
 RECT 5.425 1.945 5.79 1.96 ;
 RECT 5.425 1.115 5.74 1.255 ;
 RECT 5.6 0.8 5.74 1.115 ;
 RECT 5.425 1.255 5.565 1.805 ;
 RECT 5.51 1.96 5.79 2.215 ;
 RECT 6.465 1.295 6.605 1.805 ;
 RECT 7.125 2.11 7.265 2.355 ;
 RECT 7.125 1.36 7.265 1.97 ;
 RECT 6.05 2.355 7.265 2.495 ;
 RECT 4.505 2.52 6.19 2.655 ;
 RECT 4.785 2.515 6.19 2.52 ;
 RECT 4.505 2.655 5.065 2.66 ;
 RECT 4.025 0.845 4.165 1.125 ;
 RECT 4.27 2.15 4.41 2.335 ;
 RECT 6.05 2.495 6.19 2.515 ;
 RECT 4.505 2.475 4.645 2.52 ;
 RECT 4.27 2.335 4.645 2.475 ;
 RECT 4.025 1.125 4.41 1.265 ;
 RECT 4.27 1.265 4.41 2.01 ;
 RECT 3.83 2.01 4.41 2.15 ;
 RECT 7.125 1.97 8.67 2.11 ;
 RECT 7.615 0.405 8.12 0.445 ;
 RECT 8.53 2.11 8.67 2.425 ;
 RECT 7.615 0.445 8.365 0.585 ;
 RECT 7.615 0.585 7.755 1.22 ;
 RECT 7.125 1.22 7.755 1.36 ;
 RECT 8.53 2.425 10.025 2.565 ;
 RECT 1.04 0.82 1.18 1.18 ;
 RECT 1.04 1.32 1.18 2.325 ;
 RECT 1.835 0.38 1.975 1.18 ;
 RECT 1.04 1.18 1.975 1.32 ;
 RECT 1.835 0.24 3.25 0.38 ;
 RECT 8.41 0.885 8.55 1.675 ;
 RECT 8.34 0.745 8.615 0.885 ;
 RECT 8.335 1.685 9.545 1.825 ;
 RECT 8.34 1.675 10.6 1.685 ;
 RECT 9.36 1.545 10.6 1.675 ;
 RECT 10.305 1.505 10.535 1.545 ;
 RECT 11.02 1.095 11.16 2.375 ;
 RECT 10.305 1.685 10.6 1.745 ;
 RECT 10.46 1.745 10.6 2.375 ;
 RECT 10.46 2.375 11.16 2.515 ;
 RECT 4.735 0.835 4.875 1.13 ;
 RECT 4.735 1.41 4.875 1.495 ;
 RECT 4.735 1.13 5.005 1.41 ;
 RECT 4.67 1.635 4.81 2.045 ;
 RECT 4.785 2.185 4.925 2.315 ;
 RECT 4.67 2.045 4.925 2.185 ;
 RECT 4.67 1.495 4.875 1.635 ;
 RECT 3.095 1.03 3.235 2.13 ;
 RECT 2.585 2.13 3.235 2.27 ;
 RECT 5.13 0.665 5.27 0.845 ;
 RECT 2.395 0.89 3.84 1.03 ;
 RECT 3.7 0.665 3.84 0.89 ;
 RECT 3.7 0.525 5.27 0.665 ;
 RECT 5.145 0.985 5.285 2.005 ;
 RECT 5.085 0.845 5.34 0.985 ;
 RECT 5.085 2.005 5.285 2.305 ;
 RECT 5.42 0.375 5.79 0.425 ;
 RECT 5.42 0.425 5.795 0.52 ;
 RECT 5.42 0.535 6.83 0.66 ;
 RECT 5.42 0.52 7.305 0.535 ;
 RECT 6.69 0.395 7.305 0.52 ;
 RECT 7.075 0.245 7.305 0.395 ;
 RECT 6.845 1.025 7.15 1.08 ;
 RECT 6.845 1.08 6.985 2.2 ;
 RECT 5.975 0.94 7.15 1.025 ;
 RECT 6.975 0.68 7.475 0.885 ;
 RECT 5.725 1.4 6.115 1.54 ;
 RECT 5.975 0.885 7.475 0.94 ;
 RECT 6.98 0.675 7.475 0.68 ;
 RECT 5.975 1.025 6.115 1.4 ;
 END
END SDFFNASX2

MACRO SDFFNX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.84 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.84 2.96 ;
 RECT 1.27 2.005 1.41 2.8 ;
 RECT 3.835 2.635 4.085 2.8 ;
 RECT 6.195 2.635 6.455 2.8 ;
 RECT 9.105 1.955 9.245 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 10.745 1.7 10.885 2.8 ;
 RECT 3.18 1.98 3.32 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.84 0.08 ;
 RECT 3.81 0.08 4.11 0.26 ;
 RECT 9.11 0.08 9.365 0.285 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 6.13 0.08 6.27 0.58 ;
 RECT 10.795 0.08 10.935 0.815 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.84 1.48 2.205 1.72 ;
 RECT 2.575 1.86 2.715 1.89 ;
 RECT 1.84 1.72 2.715 1.86 ;
 RECT 2.575 1.615 2.715 1.72 ;
 RECT 1.875 1.11 2.015 1.48 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.205 2.395 2.56 2.66 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.23 2.085 10.57 2.39 ;
 RECT 10.23 0.56 10.37 2.085 ;
 END
 ANTENNADIFFAREA 0.492 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.22 2.125 11.51 2.385 ;
 RECT 11.275 2.385 11.415 2.52 ;
 RECT 11.275 0.61 11.415 2.125 ;
 END
 ANTENNADIFFAREA 0.406 ;
 END Q

 OBS
 LAYER PO ;
 RECT 9.285 1.48 9.515 1.72 ;
 RECT 6.355 0.635 6.455 1.495 ;
 RECT 6.355 1.495 6.675 1.725 ;
 RECT 6.355 1.725 6.455 2.49 ;
 RECT 3.78 1.52 4.38 1.585 ;
 RECT 5.1 1.685 5.2 2.495 ;
 RECT 4.28 0.685 4.38 1.52 ;
 RECT 3.78 1.585 5.2 1.62 ;
 RECT 4.215 1.62 5.2 1.685 ;
 RECT 4.6 0.185 6.015 0.285 ;
 RECT 4.6 0.285 4.7 0.585 ;
 RECT 4.215 1.685 4.315 2.27 ;
 RECT 3.78 1.44 4.025 1.52 ;
 RECT 3.78 1.62 4.025 1.69 ;
 RECT 5.915 0.285 6.015 1.26 ;
 RECT 4.28 0.585 4.7 0.685 ;
 RECT 5.145 0.705 5.245 1.21 ;
 RECT 4.575 1.16 4.82 1.21 ;
 RECT 4.575 1.21 5.245 1.31 ;
 RECT 4.575 1.31 4.82 1.405 ;
 RECT 5.145 0.47 5.43 0.705 ;
 RECT 7.63 0.265 7.73 0.575 ;
 RECT 7.63 0.675 7.73 1.35 ;
 RECT 6.825 0.575 7.73 0.675 ;
 RECT 8.075 1.545 8.175 2.405 ;
 RECT 8.965 0.265 9.065 1.32 ;
 RECT 6.825 0.46 7.055 0.575 ;
 RECT 6.825 0.675 7.055 0.69 ;
 RECT 7.82 1.45 8.175 1.545 ;
 RECT 7.63 0.165 9.065 0.265 ;
 RECT 7.63 1.35 7.92 1.445 ;
 RECT 7.63 1.445 8.175 1.45 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 8.89 1.64 8.99 2.585 ;
 RECT 7.67 2.47 7.89 2.585 ;
 RECT 7.67 2.685 7.89 2.71 ;
 RECT 7.67 2.585 8.99 2.685 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 8.57 0.645 8.67 1.24 ;
 RECT 8.57 1.45 8.67 2.37 ;
 RECT 8.55 1.24 8.785 1.45 ;
 RECT 8.1 0.685 8.2 1.255 ;
 RECT 8.025 0.455 8.255 0.685 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.245 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 9.905 1.225 10.585 1.455 ;
 RECT 10.485 0.14 10.585 1.225 ;
 RECT 10.485 1.455 10.585 2.775 ;
 RECT 11.06 0.33 11.16 1.225 ;
 RECT 11.06 1.46 11.16 2.775 ;
 RECT 10.86 1.225 11.16 1.46 ;
 RECT 2.195 1.745 2.295 2.44 ;
 RECT 2.195 2.44 2.445 2.67 ;
 RECT 2.245 1.345 2.345 1.645 ;
 RECT 2.665 0.655 2.765 1.245 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.245 1.245 2.765 1.345 ;
 RECT 4.62 2.33 4.72 2.685 ;
 RECT 4.62 2.685 6.015 2.785 ;
 RECT 5.915 1.7 6.015 2.685 ;
 RECT 4.5 2.09 4.72 2.33 ;
 RECT 5.595 1.37 5.735 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.595 1.33 5.715 1.37 ;
 RECT 5.48 1.475 5.735 1.5 ;
 RECT 5.48 1.5 5.71 1.71 ;
 RECT 5.615 0.65 5.715 1.33 ;
 RECT 7.05 0.875 7.38 1.105 ;
 RECT 7.28 1.105 7.38 1.64 ;
 RECT 7.28 1.64 7.515 1.87 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 2.665 1.865 2.765 2.48 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 9.38 0.65 9.48 1.48 ;
 RECT 9.38 1.72 9.48 2.56 ;
 LAYER CO ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 6.865 0.51 6.995 0.64 ;
 RECT 9.34 1.535 9.47 1.665 ;
 RECT 10.235 2.13 10.365 2.26 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 2.265 2.49 2.395 2.62 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 4.63 1.205 4.76 1.335 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 5.53 1.525 5.66 1.655 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 10.75 2.29 10.88 2.42 ;
 RECT 11.28 2.32 11.41 2.45 ;
 RECT 9.955 1.275 10.085 1.405 ;
 RECT 7.335 1.69 7.465 1.82 ;
 RECT 7.12 0.915 7.25 1.045 ;
 RECT 9.185 0.15 9.315 0.28 ;
 RECT 3.84 1.495 3.97 1.625 ;
 RECT 3.905 2.64 4.035 2.77 ;
 RECT 8.075 0.505 8.205 0.635 ;
 RECT 8.6 1.28 8.73 1.41 ;
 RECT 9.6 0.87 9.73 1 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 3.295 1.535 3.425 1.665 ;
 RECT 6.78 0.88 6.91 1.01 ;
 RECT 6.775 2.015 6.905 2.145 ;
 RECT 3.93 0.125 4.06 0.255 ;
 RECT 6.245 2.64 6.375 2.77 ;
 RECT 7.72 2.525 7.85 2.655 ;
 RECT 7.825 1.815 7.955 1.945 ;
 RECT 10.9 1.275 11.03 1.405 ;
 RECT 11.28 0.68 11.41 0.81 ;
 RECT 10.75 1.77 10.88 1.9 ;
 RECT 10.75 2.03 10.88 2.16 ;
 RECT 4.55 2.145 4.68 2.275 ;
 RECT 10.235 0.63 10.365 0.76 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 9.11 2.01 9.24 2.14 ;
 RECT 9.67 2.13 9.8 2.26 ;
 RECT 6.49 1.535 6.62 1.665 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 3.71 1.995 3.84 2.125 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 11.28 1.8 11.41 1.93 ;
 RECT 11.28 2.06 11.41 2.19 ;
 RECT 10.8 0.615 10.93 0.745 ;
 RECT 10.235 1.87 10.365 2 ;
 RECT 4.435 1.825 4.565 1.955 ;
 RECT 5.25 0.525 5.38 0.655 ;
 RECT 6.135 0.38 6.265 0.51 ;
 RECT 8.32 1.9 8.45 2.03 ;
 RECT 8.32 0.87 8.45 1 ;
 RECT 7.85 0.87 7.98 1 ;
 LAYER M1 ;
 RECT 6.77 1.05 6.91 1.185 ;
 RECT 6.77 1.325 6.91 2.215 ;
 RECT 5.985 1.185 6.91 1.325 ;
 RECT 5.465 1.52 6.125 1.66 ;
 RECT 6.71 0.91 7.32 1.015 ;
 RECT 6.71 0.875 6.98 0.91 ;
 RECT 6.77 1.015 7.32 1.05 ;
 RECT 5.985 1.325 6.125 1.52 ;
 RECT 5.18 0.52 5.78 0.66 ;
 RECT 5.64 0.66 5.78 0.79 ;
 RECT 5.64 0.79 6.55 0.93 ;
 RECT 6.41 0.505 7.045 0.645 ;
 RECT 6.41 0.645 6.55 0.79 ;
 RECT 9.595 0.36 9.735 0.965 ;
 RECT 9.665 1.105 9.805 1.245 ;
 RECT 9.665 1.385 9.805 2.33 ;
 RECT 8.595 1.245 9.81 1.385 ;
 RECT 9.595 0.965 9.805 1.105 ;
 RECT 8.595 1.21 8.735 1.245 ;
 RECT 8.595 1.385 8.735 1.465 ;
 RECT 10.515 0.36 10.655 1.27 ;
 RECT 9.595 0.22 10.655 0.36 ;
 RECT 10.895 1.2 11.035 1.27 ;
 RECT 10.895 1.41 11.035 1.48 ;
 RECT 10.515 1.27 11.035 1.41 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.365 2.11 2.995 2.195 ;
 RECT 2.365 2.195 2.99 2.25 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 3.46 0.53 4.41 0.67 ;
 RECT 4.27 0.22 5.03 0.36 ;
 RECT 4.89 0.36 5.03 0.875 ;
 RECT 4.905 1.015 5.045 2.035 ;
 RECT 4.845 2.035 5.045 2.17 ;
 RECT 4.845 2.17 4.985 2.305 ;
 RECT 4.27 0.36 4.41 0.53 ;
 RECT 4.825 0.875 5.1 1.015 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 8.315 1.815 8.525 1.895 ;
 RECT 8.315 0.805 8.455 1.675 ;
 RECT 8.245 1.895 8.525 2.035 ;
 RECT 8.315 1.675 9.175 1.815 ;
 RECT 9.035 1.67 9.175 1.675 ;
 RECT 9.95 1.205 10.09 2.505 ;
 RECT 9.035 1.53 9.525 1.67 ;
 RECT 9.385 2.505 10.09 2.645 ;
 RECT 9.385 1.67 9.525 2.505 ;
 RECT 4.495 1.385 4.635 1.82 ;
 RECT 4.365 1.825 4.685 1.96 ;
 RECT 4.365 1.82 4.635 1.825 ;
 RECT 4.545 1.96 4.685 2.345 ;
 RECT 4.495 0.84 4.635 1.155 ;
 RECT 4.495 1.155 4.765 1.385 ;
 RECT 4.225 2.515 5.76 2.65 ;
 RECT 4.225 2.65 5.515 2.655 ;
 RECT 5.08 2.51 5.76 2.515 ;
 RECT 4.225 2.49 4.365 2.515 ;
 RECT 3.705 1.63 3.845 2.35 ;
 RECT 3.705 1.475 4.045 1.63 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 5.62 2.495 5.76 2.51 ;
 RECT 3.705 2.35 4.365 2.49 ;
 RECT 7.49 0.58 8.28 0.64 ;
 RECT 7.49 0.64 7.95 0.72 ;
 RECT 7.77 0.5 8.28 0.58 ;
 RECT 7.05 1.21 7.63 1.35 ;
 RECT 7.05 1.35 7.19 2.1 ;
 RECT 7.05 2.1 7.79 2.24 ;
 RECT 7.05 2.24 7.19 2.355 ;
 RECT 7.65 2.24 7.79 2.52 ;
 RECT 5.62 2.355 7.19 2.495 ;
 RECT 7.65 2.52 7.92 2.66 ;
 RECT 7.49 0.72 7.63 1.21 ;
 RECT 7.33 1.685 7.985 1.81 ;
 RECT 7.845 1.005 7.985 1.685 ;
 RECT 7.33 1.81 8.025 1.825 ;
 RECT 7.33 1.825 7.47 1.89 ;
 RECT 7.33 1.62 7.47 1.685 ;
 RECT 7.755 1.825 8.025 1.95 ;
 RECT 7.775 0.865 8.055 1.005 ;
 RECT 5.185 1.82 6.625 1.955 ;
 RECT 5.185 1.955 6.12 1.96 ;
 RECT 6.485 1.465 6.625 1.815 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 5.36 0.805 5.5 1.22 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 5.95 1.815 6.625 1.82 ;
 RECT 5.185 1.36 5.325 1.82 ;
 END
END SDFFNX1

MACRO SDFFNX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 12.8 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 12.8 2.96 ;
 RECT 6.195 2.635 6.455 2.8 ;
 RECT 1.27 2.005 1.41 2.8 ;
 RECT 3.835 2.625 4.085 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 10.385 1.51 10.525 2.8 ;
 RECT 11.335 1.51 11.475 2.8 ;
 RECT 12.275 1.51 12.415 2.8 ;
 RECT 3.18 1.98 3.32 2.8 ;
 RECT 9.105 1.955 9.245 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 12.8 0.08 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 3.81 0.08 4.11 0.26 ;
 RECT 11.255 0.08 11.51 0.285 ;
 RECT 9.11 0.08 9.365 0.285 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 6.13 0.08 6.27 0.58 ;
 RECT 10.295 0.08 10.435 0.695 ;
 RECT 12.28 0.08 12.42 0.86 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.162 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.595 2.075 2.015 2.45 ;
 RECT 2.575 1.86 2.715 1.89 ;
 RECT 1.875 1.72 2.715 1.86 ;
 RECT 2.575 1.615 2.715 1.72 ;
 RECT 1.875 1.86 2.015 2.075 ;
 RECT 1.875 1.11 2.015 1.72 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.225 1.18 2.58 1.445 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.855 2.085 11.195 2.39 ;
 RECT 10.855 2.39 10.995 2.575 ;
 RECT 10.855 0.72 10.995 2.085 ;
 END
 ANTENNADIFFAREA 0.58 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.7 2.08 12.005 2.385 ;
 RECT 11.805 2.385 11.945 2.575 ;
 RECT 11.805 0.61 11.945 2.08 ;
 END
 ANTENNADIFFAREA 0.562 ;
 END Q

 OBS
 LAYER PO ;
 RECT 5.145 0.705 5.245 1.155 ;
 RECT 4.565 1.255 4.82 1.395 ;
 RECT 4.565 1.155 5.245 1.255 ;
 RECT 6.355 0.635 6.455 1.465 ;
 RECT 6.355 1.465 6.675 1.695 ;
 RECT 6.355 1.695 6.455 2.54 ;
 RECT 5.595 1.66 5.695 2.505 ;
 RECT 5.595 1.33 5.715 1.425 ;
 RECT 5.48 1.425 5.715 1.66 ;
 RECT 5.615 0.65 5.715 1.33 ;
 RECT 2.665 0.655 2.765 1.245 ;
 RECT 2.245 1.225 2.465 1.245 ;
 RECT 2.245 1.345 2.465 1.455 ;
 RECT 2.245 1.455 2.345 1.645 ;
 RECT 2.245 1.245 2.765 1.345 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.195 1.745 2.295 2.74 ;
 RECT 7.63 0.265 7.73 0.575 ;
 RECT 6.805 0.575 7.73 0.675 ;
 RECT 7.63 0.675 7.73 1.35 ;
 RECT 8.075 1.545 8.175 2.505 ;
 RECT 6.805 0.405 7.075 0.575 ;
 RECT 8.965 0.265 9.065 1.32 ;
 RECT 7.82 1.45 8.175 1.545 ;
 RECT 7.63 1.35 7.92 1.445 ;
 RECT 7.63 1.445 8.175 1.45 ;
 RECT 7.63 0.165 9.065 0.265 ;
 RECT 9.905 1.075 10.74 1.105 ;
 RECT 9.905 1.205 10.74 1.305 ;
 RECT 11.11 0.19 11.21 1.105 ;
 RECT 11.11 1.205 11.21 2.79 ;
 RECT 9.905 1.105 11.21 1.205 ;
 RECT 10.64 0.195 10.74 1.075 ;
 RECT 10.64 1.305 10.74 2.79 ;
 RECT 11.39 1.035 11.69 1.105 ;
 RECT 11.39 1.205 11.69 1.27 ;
 RECT 11.39 1.105 12.16 1.205 ;
 RECT 12.06 0.25 12.16 1.105 ;
 RECT 12.06 1.205 12.16 2.79 ;
 RECT 11.59 0.285 11.69 1.035 ;
 RECT 11.59 1.27 11.69 2.79 ;
 RECT 9.38 0.65 9.48 1.48 ;
 RECT 9.38 1.745 9.48 2.79 ;
 RECT 9.34 1.48 9.57 1.745 ;
 RECT 4.07 1.49 4.38 1.575 ;
 RECT 4.07 1.575 5.2 1.675 ;
 RECT 5.1 1.675 5.2 2.505 ;
 RECT 5.1 1.535 5.2 1.575 ;
 RECT 4.28 0.285 4.38 1.49 ;
 RECT 4.07 1.675 4.315 1.735 ;
 RECT 4.215 1.735 4.315 2.295 ;
 RECT 4.28 0.185 6.015 0.285 ;
 RECT 5.915 0.285 6.015 1.26 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.245 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 2.965 0.405 3.065 2.73 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 5.915 1.535 6.015 2.685 ;
 RECT 4.495 2.075 4.71 2.685 ;
 RECT 4.495 2.685 6.015 2.785 ;
 RECT 8.89 1.545 8.99 2.69 ;
 RECT 7.67 2.46 7.89 2.69 ;
 RECT 7.67 2.69 8.99 2.79 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.605 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.73 ;
 RECT 7.05 0.875 7.38 1.105 ;
 RECT 7.28 1.105 7.38 1.64 ;
 RECT 7.28 1.64 7.515 1.87 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 2.665 1.865 2.765 2.73 ;
 RECT 8.57 0.645 8.67 1.155 ;
 RECT 8.57 1.365 8.67 2.505 ;
 RECT 8.55 1.155 8.785 1.365 ;
 RECT 8.1 0.685 8.2 1.255 ;
 RECT 8.025 0.455 8.255 0.685 ;
 RECT 5.145 0.47 5.435 0.705 ;
 LAYER CO ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 11.81 2.115 11.94 2.245 ;
 RECT 11.81 2.375 11.94 2.505 ;
 RECT 11.81 1.59 11.94 1.72 ;
 RECT 10.39 1.59 10.52 1.72 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 4.125 1.535 4.255 1.665 ;
 RECT 7.72 2.515 7.85 2.645 ;
 RECT 7.825 1.815 7.955 1.945 ;
 RECT 8.6 1.195 8.73 1.325 ;
 RECT 9.6 0.87 9.73 1 ;
 RECT 9.11 2.01 9.24 2.14 ;
 RECT 10.86 2.115 10.99 2.245 ;
 RECT 10.86 2.375 10.99 2.505 ;
 RECT 10.86 0.77 10.99 0.9 ;
 RECT 5.53 1.475 5.66 1.605 ;
 RECT 6.775 0.88 6.905 1.01 ;
 RECT 6.775 2.015 6.905 2.145 ;
 RECT 3.93 0.125 4.06 0.255 ;
 RECT 7.335 1.69 7.465 1.82 ;
 RECT 7.12 0.915 7.25 1.045 ;
 RECT 9.185 0.15 9.315 0.28 ;
 RECT 3.905 2.63 4.035 2.76 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 3.295 1.535 3.425 1.665 ;
 RECT 3.71 1.985 3.84 2.115 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 12.28 1.85 12.41 1.98 ;
 RECT 12.28 2.115 12.41 2.245 ;
 RECT 12.28 2.375 12.41 2.505 ;
 RECT 12.28 1.59 12.41 1.72 ;
 RECT 11.33 0.15 11.46 0.28 ;
 RECT 10.3 0.495 10.43 0.625 ;
 RECT 4.54 2.125 4.67 2.255 ;
 RECT 12.285 0.68 12.415 0.81 ;
 RECT 11.34 2.375 11.47 2.505 ;
 RECT 11.34 1.59 11.47 1.72 ;
 RECT 11.34 1.85 11.47 1.98 ;
 RECT 11.34 2.115 11.47 2.245 ;
 RECT 11.81 1.85 11.94 1.98 ;
 RECT 10.39 1.85 10.52 1.98 ;
 RECT 10.39 2.115 10.52 2.245 ;
 RECT 10.39 2.375 10.52 2.505 ;
 RECT 10.86 1.59 10.99 1.72 ;
 RECT 10.86 1.85 10.99 1.98 ;
 RECT 5.255 0.525 5.385 0.655 ;
 RECT 6.865 0.45 6.995 0.58 ;
 RECT 9.39 1.55 9.52 1.68 ;
 RECT 4.435 1.825 4.565 1.955 ;
 RECT 11.43 1.085 11.56 1.215 ;
 RECT 11.81 0.68 11.94 0.81 ;
 RECT 10.105 1.125 10.235 1.255 ;
 RECT 2.285 1.275 2.415 1.405 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 6.135 0.38 6.265 0.51 ;
 RECT 8.32 1.9 8.45 2.03 ;
 RECT 8.32 0.87 8.45 1 ;
 RECT 7.85 0.87 7.98 1 ;
 RECT 8.075 0.505 8.205 0.635 ;
 RECT 4.615 1.22 4.745 1.35 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 9.67 2.13 9.8 2.26 ;
 RECT 6.49 1.505 6.62 1.635 ;
 RECT 6.245 2.64 6.375 2.77 ;
 LAYER M1 ;
 RECT 5.18 0.52 5.85 0.66 ;
 RECT 5.71 0.66 5.85 0.79 ;
 RECT 6.41 0.445 7.045 0.585 ;
 RECT 5.71 0.79 6.55 0.93 ;
 RECT 6.41 0.585 6.55 0.79 ;
 RECT 5.465 1.47 6.125 1.61 ;
 RECT 6.77 0.875 7.32 1.05 ;
 RECT 6.77 0.805 6.91 0.875 ;
 RECT 6.77 1.05 6.91 1.075 ;
 RECT 6.77 1.215 6.91 2.215 ;
 RECT 5.985 1.075 6.91 1.215 ;
 RECT 5.95 1.61 6.125 1.66 ;
 RECT 5.985 1.215 6.125 1.47 ;
 RECT 8.315 1.815 8.525 1.895 ;
 RECT 8.315 0.805 8.455 1.675 ;
 RECT 8.245 1.895 8.525 2.035 ;
 RECT 9.95 1.26 10.09 2.505 ;
 RECT 9.035 1.545 9.525 1.675 ;
 RECT 8.315 1.675 9.525 1.685 ;
 RECT 9.385 1.475 9.525 1.545 ;
 RECT 9.385 1.685 9.525 2.52 ;
 RECT 8.315 1.685 9.175 1.815 ;
 RECT 9.87 2.505 10.09 2.52 ;
 RECT 9.95 1.12 10.305 1.26 ;
 RECT 9.385 2.52 10.09 2.66 ;
 RECT 7.33 1.685 7.985 1.81 ;
 RECT 7.845 1.005 7.985 1.685 ;
 RECT 7.33 1.81 8.025 1.825 ;
 RECT 7.33 1.825 7.47 1.89 ;
 RECT 7.33 1.62 7.47 1.685 ;
 RECT 7.755 1.825 8.025 1.95 ;
 RECT 7.775 0.865 8.055 1.005 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 10.575 0.58 10.715 0.835 ;
 RECT 9.595 0.835 10.715 0.975 ;
 RECT 9.595 0.975 9.805 1.19 ;
 RECT 9.665 1.33 9.805 2.33 ;
 RECT 9.595 0.785 9.735 0.835 ;
 RECT 8.595 1.19 9.805 1.33 ;
 RECT 8.595 1.125 8.735 1.19 ;
 RECT 8.595 1.33 8.735 1.38 ;
 RECT 11.425 0.58 11.565 1.29 ;
 RECT 10.575 0.44 11.565 0.58 ;
 RECT 3.705 1.53 4.325 1.67 ;
 RECT 3.705 1.475 3.925 1.53 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.705 1.67 3.845 2.345 ;
 RECT 4.225 2.51 5.76 2.65 ;
 RECT 3.705 2.345 4.365 2.485 ;
 RECT 4.225 2.485 4.365 2.51 ;
 RECT 5.62 2.495 5.76 2.51 ;
 RECT 5.62 2.355 7.19 2.495 ;
 RECT 7.65 2.24 7.79 2.51 ;
 RECT 7.05 2.24 7.19 2.355 ;
 RECT 7.05 1.35 7.19 2.1 ;
 RECT 7.05 2.1 7.79 2.24 ;
 RECT 7.05 1.21 7.63 1.35 ;
 RECT 7.65 2.51 7.92 2.65 ;
 RECT 7.77 0.5 8.28 0.58 ;
 RECT 7.49 0.58 8.28 0.64 ;
 RECT 7.49 0.64 7.95 0.72 ;
 RECT 7.49 0.72 7.63 1.21 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.365 2.11 2.995 2.25 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 3.46 0.53 5.03 0.67 ;
 RECT 4.89 0.67 5.03 0.8 ;
 RECT 4.89 0.8 5.045 1.095 ;
 RECT 4.905 1.095 5.045 2.035 ;
 RECT 4.845 2.035 5.045 2.305 ;
 RECT 4.495 1.44 4.675 1.82 ;
 RECT 4.535 1.96 4.675 2.325 ;
 RECT 4.365 1.82 4.675 1.96 ;
 RECT 4.495 0.825 4.75 1.44 ;
 RECT 5.185 1.82 6.625 1.96 ;
 RECT 6.485 1.435 6.625 1.82 ;
 RECT 5.185 0.875 5.57 1.015 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 5.185 1.015 5.325 1.82 ;
 END
END SDFFNX2

MACRO SDFFSSRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 13.76 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 13.76 2.96 ;
 RECT 6.645 2.275 6.895 2.8 ;
 RECT 9.005 2.63 9.265 2.8 ;
 RECT 2.845 1.955 2.985 2.8 ;
 RECT 12.595 1.505 12.735 2.8 ;
 RECT 0.94 1.975 1.08 2.8 ;
 RECT 11.12 1.95 11.26 2.8 ;
 RECT 6.045 1.945 6.185 2.8 ;
 RECT 4.13 1.96 4.27 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 13.76 0.08 ;
 RECT 10.875 0.08 11.13 0.28 ;
 RECT 0.835 0.08 1.135 0.26 ;
 RECT 6.62 0.08 6.92 0.255 ;
 RECT 3.165 0.08 3.305 0.77 ;
 RECT 8.94 0.08 9.08 0.575 ;
 RECT 12.645 0.08 12.785 0.81 ;
 RECT 4.13 0.08 4.27 0.65 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.325 1.47 6.715 1.78 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.08 2.08 12.455 2.385 ;
 RECT 12.08 2.385 12.22 2.57 ;
 RECT 12.08 0.555 12.22 2.08 ;
 END
 ANTENNADIFFAREA 0.527 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.08 2.075 13.455 2.38 ;
 RECT 13.125 2.38 13.265 2.57 ;
 RECT 13.125 0.605 13.265 2.075 ;
 END
 ANTENNADIFFAREA 0.47 ;
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.55 1.455 1.93 1.735 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.655 1.48 0.97 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SETB

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.92 1.16 3.285 1.44 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.53 0.22 3.99 0.635 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4 1.15 4.535 1.41 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 OBS
 LAYER PO ;
 RECT 11.395 1.435 11.495 2.69 ;
 RECT 12.335 0.19 12.435 1.13 ;
 RECT 12.335 1.36 12.435 2.785 ;
 RECT 12.91 0.255 13.01 1.03 ;
 RECT 12.91 1.265 13.01 2.785 ;
 RECT 12.71 1.03 13.01 1.265 ;
 RECT 6.88 1.485 7.19 1.615 ;
 RECT 7.025 1.73 7.125 2.68 ;
 RECT 7.09 1.25 7.19 1.485 ;
 RECT 7.955 0.465 8.245 0.7 ;
 RECT 7.955 0.7 8.055 1.15 ;
 RECT 8.725 1.775 8.825 2.68 ;
 RECT 7.09 0.68 7.19 1.15 ;
 RECT 6.88 1.615 7.125 1.73 ;
 RECT 7.025 2.68 8.825 2.78 ;
 RECT 7.09 1.15 8.055 1.25 ;
 RECT 9.935 1.5 10.035 2.265 ;
 RECT 9.935 2.265 10.455 2.505 ;
 RECT 2.83 1.42 2.93 1.71 ;
 RECT 2.135 1.81 2.235 2.465 ;
 RECT 2.83 0.565 2.93 1.185 ;
 RECT 1.195 0.565 1.295 1.325 ;
 RECT 2.83 1.185 3.235 1.42 ;
 RECT 2.135 1.71 2.93 1.81 ;
 RECT 1.195 0.465 2.93 0.565 ;
 RECT 10.255 0.44 10.53 0.65 ;
 RECT 10.43 0.65 10.53 2.085 ;
 RECT 9.96 0.68 10.06 1.25 ;
 RECT 9.825 0.45 10.06 0.68 ;
 RECT 5.415 0.41 5.515 1.215 ;
 RECT 5.34 0.175 5.57 0.41 ;
 RECT 4.945 1.685 5.045 2.565 ;
 RECT 3.4 2.565 5.045 2.665 ;
 RECT 3.4 1.965 3.63 2.565 ;
 RECT 7.91 1.67 8.01 2.49 ;
 RECT 7.385 1.485 7.63 1.57 ;
 RECT 7.385 1.67 7.63 1.73 ;
 RECT 7.385 1.57 8.01 1.67 ;
 RECT 10.905 1.635 11.005 2.685 ;
 RECT 9.53 2.38 9.75 2.685 ;
 RECT 9.53 2.685 11.005 2.785 ;
 RECT 0.725 0.565 0.825 1.485 ;
 RECT 0.725 1.72 0.825 2.465 ;
 RECT 0.69 1.485 0.92 1.72 ;
 RECT 1.195 1.775 1.295 2.675 ;
 RECT 0.28 2.375 0.51 2.675 ;
 RECT 0.28 2.675 1.295 2.775 ;
 RECT 2.135 0.745 2.235 1.28 ;
 RECT 2.135 1.28 2.645 1.515 ;
 RECT 7.41 0.18 8.825 0.28 ;
 RECT 7.41 0.28 7.51 0.52 ;
 RECT 8.725 0.28 8.825 1.255 ;
 RECT 7.37 0.52 7.6 0.755 ;
 RECT 1.665 0.745 1.765 1.475 ;
 RECT 1.665 1.71 1.765 2.465 ;
 RECT 1.62 1.475 1.85 1.71 ;
 RECT 3.705 0.315 4.015 0.45 ;
 RECT 3.915 0.45 4.015 2.385 ;
 RECT 4.945 0.315 5.045 1.395 ;
 RECT 4.94 1.395 5.515 1.495 ;
 RECT 5.415 1.495 5.515 2.395 ;
 RECT 3.705 0.215 5.045 0.315 ;
 RECT 4.475 0.64 4.575 1.155 ;
 RECT 4.475 1.39 4.575 2.385 ;
 RECT 4.195 1.155 4.575 1.39 ;
 RECT 10.73 0.26 10.83 1.155 ;
 RECT 9.2 0.26 9.505 0.43 ;
 RECT 10.73 1.155 10.965 1.365 ;
 RECT 9.2 0.16 10.83 0.26 ;
 RECT 9.165 0.655 9.265 1.585 ;
 RECT 9.165 1.815 9.265 2.485 ;
 RECT 9.115 1.585 9.355 1.815 ;
 RECT 8.405 1.325 8.525 1.475 ;
 RECT 8.405 1.71 8.505 2.47 ;
 RECT 8.425 0.645 8.525 1.325 ;
 RECT 8.325 1.475 8.555 1.71 ;
 RECT 6.485 1.295 6.585 1.475 ;
 RECT 6.485 1.195 6.87 1.295 ;
 RECT 6.77 0.635 6.87 1.195 ;
 RECT 6.3 1.715 6.4 2.365 ;
 RECT 6.3 1.475 6.595 1.715 ;
 RECT 11.145 1.2 12.435 1.36 ;
 RECT 11.575 1.13 12.435 1.2 ;
 RECT 11.145 1.36 12.07 1.435 ;
 RECT 11.185 0.5 11.285 1.2 ;
 LAYER CO ;
 RECT 9.055 2.635 9.185 2.765 ;
 RECT 9.58 2.43 9.71 2.56 ;
 RECT 9.585 1.75 9.715 1.88 ;
 RECT 12.75 1.08 12.88 1.21 ;
 RECT 5.39 0.23 5.52 0.36 ;
 RECT 3.46 2.025 3.59 2.155 ;
 RECT 6.715 2.38 6.845 2.51 ;
 RECT 7.705 0.875 7.835 1.005 ;
 RECT 7.44 1.53 7.57 1.66 ;
 RECT 7.31 0.9 7.44 1.03 ;
 RECT 6.425 1.53 6.555 1.66 ;
 RECT 3.575 1.685 3.705 1.815 ;
 RECT 4.135 0.435 4.265 0.565 ;
 RECT 4.135 2.03 4.265 2.16 ;
 RECT 4.695 0.865 4.825 0.995 ;
 RECT 4.695 1.995 4.825 2.125 ;
 RECT 5.165 0.865 5.295 0.995 ;
 RECT 5.165 1.995 5.295 2.125 ;
 RECT 2.465 1.335 2.595 1.465 ;
 RECT 2.355 2.05 2.485 2.18 ;
 RECT 2.355 0.97 2.485 1.1 ;
 RECT 1.885 2.05 2.015 2.18 ;
 RECT 1.885 0.97 2.015 1.1 ;
 RECT 0.475 2.05 0.605 2.18 ;
 RECT 0.475 0.79 0.605 0.92 ;
 RECT 6.52 0.9 6.65 1.03 ;
 RECT 6.05 1.995 6.18 2.125 ;
 RECT 10.285 2.325 10.415 2.455 ;
 RECT 10.78 1.195 10.91 1.325 ;
 RECT 0.955 0.125 1.085 0.255 ;
 RECT 0.74 1.54 0.87 1.67 ;
 RECT 12.6 2.37 12.73 2.5 ;
 RECT 12.085 1.585 12.215 1.715 ;
 RECT 12.085 1.845 12.215 1.975 ;
 RECT 6.935 1.53 7.065 1.66 ;
 RECT 8.065 0.52 8.195 0.65 ;
 RECT 0.33 2.43 0.46 2.56 ;
 RECT 0.945 2.05 1.075 2.18 ;
 RECT 1.415 2.05 1.545 2.18 ;
 RECT 1.415 0.97 1.545 1.1 ;
 RECT 7.245 1.82 7.375 1.95 ;
 RECT 7.42 0.575 7.55 0.705 ;
 RECT 1.67 1.53 1.8 1.66 ;
 RECT 2.85 2.34 2.98 2.47 ;
 RECT 2.85 2.08 2.98 2.21 ;
 RECT 13.13 1.845 13.26 1.975 ;
 RECT 13.13 2.11 13.26 2.24 ;
 RECT 13.13 2.37 13.26 2.5 ;
 RECT 13.13 1.585 13.26 1.715 ;
 RECT 12.6 1.585 12.73 1.715 ;
 RECT 13.13 0.675 13.26 0.805 ;
 RECT 4.32 1.21 4.45 1.34 ;
 RECT 8.945 0.375 9.075 0.505 ;
 RECT 10.18 1.895 10.31 2.025 ;
 RECT 10.18 0.865 10.31 0.995 ;
 RECT 9.875 0.5 10.005 0.63 ;
 RECT 8.155 2.065 8.285 2.195 ;
 RECT 8.175 0.875 8.305 1.005 ;
 RECT 7.66 2.1 7.79 2.23 ;
 RECT 11.615 1.96 11.745 2.09 ;
 RECT 9.17 1.625 9.3 1.755 ;
 RECT 6.52 1.995 6.65 2.125 ;
 RECT 3.775 0.255 3.905 0.385 ;
 RECT 3.665 0.865 3.795 0.995 ;
 RECT 5.635 0.865 5.765 0.995 ;
 RECT 5.635 1.995 5.765 2.125 ;
 RECT 3.055 1.24 3.185 1.37 ;
 RECT 12.6 1.845 12.73 1.975 ;
 RECT 12.6 2.11 12.73 2.24 ;
 RECT 12.65 0.61 12.78 0.74 ;
 RECT 12.085 2.11 12.215 2.24 ;
 RECT 12.085 2.37 12.215 2.5 ;
 RECT 12.085 0.625 12.215 0.755 ;
 RECT 10.95 0.145 11.08 0.275 ;
 RECT 9.315 0.25 9.445 0.38 ;
 RECT 11.2 1.245 11.33 1.375 ;
 RECT 10.305 0.48 10.435 0.61 ;
 RECT 11.41 0.865 11.54 0.995 ;
 RECT 11.125 2.005 11.255 2.135 ;
 RECT 3.17 0.585 3.3 0.715 ;
 RECT 3.17 0.325 3.3 0.455 ;
 RECT 8.375 1.525 8.505 1.655 ;
 RECT 9.585 0.875 9.715 1.005 ;
 RECT 9.585 2.01 9.715 2.14 ;
 RECT 6.74 0.12 6.87 0.25 ;
 LAYER M1 ;
 RECT 4.69 0.675 4.83 2.175 ;
 RECT 1.41 2.465 2.49 2.605 ;
 RECT 2.35 1.98 2.49 2.465 ;
 RECT 1.41 1.98 1.55 2.465 ;
 RECT 1.41 0.825 1.55 0.965 ;
 RECT 1.41 0.685 2.49 0.825 ;
 RECT 2.35 0.825 2.49 1.16 ;
 RECT 1.335 0.965 1.62 1.105 ;
 RECT 10.585 1.19 10.98 1.33 ;
 RECT 10.585 1.33 10.725 2.32 ;
 RECT 10.195 2.32 10.725 2.46 ;
 RECT 7.99 0.515 8.8 0.655 ;
 RECT 8.66 0.655 8.8 0.785 ;
 RECT 8.66 0.785 9.36 0.925 ;
 RECT 9.22 0.245 9.515 0.385 ;
 RECT 9.22 0.385 9.36 0.785 ;
 RECT 8.275 1.52 8.935 1.655 ;
 RECT 8.76 1.515 8.935 1.52 ;
 RECT 8.275 1.655 8.93 1.66 ;
 RECT 8.795 1.18 9.72 1.32 ;
 RECT 9.58 0.805 9.72 1.18 ;
 RECT 9.58 1.32 9.72 2.21 ;
 RECT 8.795 1.32 8.935 1.515 ;
 RECT 3.455 1.96 3.71 2.26 ;
 RECT 3.57 1 3.71 1.96 ;
 RECT 4.41 0.365 4.55 0.86 ;
 RECT 3.57 0.86 4.55 1 ;
 RECT 4.41 1 4.55 1.005 ;
 RECT 4.41 0.225 5.6 0.365 ;
 RECT 2.07 1.67 3.3 1.81 ;
 RECT 3.16 1.81 3.3 2.515 ;
 RECT 3.85 1.82 3.99 2.515 ;
 RECT 3.16 2.515 3.99 2.655 ;
 RECT 2.07 1.81 2.21 1.9 ;
 RECT 1.88 2.04 2.02 2.255 ;
 RECT 1.805 0.965 2.21 1.105 ;
 RECT 2.07 1.105 2.21 1.67 ;
 RECT 1.88 1.9 2.21 2.04 ;
 RECT 4.41 1.82 4.55 2.315 ;
 RECT 5.63 0.785 5.77 2.315 ;
 RECT 3.85 1.68 4.55 1.82 ;
 RECT 4.41 2.315 5.77 2.455 ;
 RECT 0.325 0.925 0.465 2.045 ;
 RECT 0.325 0.54 0.465 0.785 ;
 RECT 0.325 2.185 0.465 2.63 ;
 RECT 0.325 2.045 0.665 2.185 ;
 RECT 0.325 0.785 0.675 0.925 ;
 RECT 2.35 1.33 2.77 1.47 ;
 RECT 2.63 0.54 2.77 1.33 ;
 RECT 0.325 0.4 2.77 0.54 ;
 RECT 5.155 0.645 5.3 0.67 ;
 RECT 5.16 0.67 5.3 2.175 ;
 RECT 5.155 0.505 7.23 0.645 ;
 RECT 7.7 0.36 7.84 0.795 ;
 RECT 7.09 0.36 7.23 0.505 ;
 RECT 7.09 0.22 7.84 0.36 ;
 RECT 7.7 0.795 7.855 1.09 ;
 RECT 7.715 1.09 7.855 2.03 ;
 RECT 7.655 2.03 7.855 2.3 ;
 RECT 7.175 1.815 7.495 1.955 ;
 RECT 7.355 1.955 7.495 2.505 ;
 RECT 7.355 2.505 8.57 2.645 ;
 RECT 7.305 1.71 7.495 1.815 ;
 RECT 8.43 2.49 8.57 2.505 ;
 RECT 7.415 0.505 7.555 0.835 ;
 RECT 7.305 0.835 7.555 1.03 ;
 RECT 7.305 1.03 7.445 1.48 ;
 RECT 7.305 1.48 7.575 1.71 ;
 RECT 9.405 2.49 10.01 2.565 ;
 RECT 8.43 2.35 9.545 2.425 ;
 RECT 8.43 2.425 10.01 2.49 ;
 RECT 9.87 0.445 10.01 2.425 ;
 RECT 7.995 1.815 9.305 1.955 ;
 RECT 8.17 1.01 8.31 1.215 ;
 RECT 9.165 1.555 9.305 1.815 ;
 RECT 7.995 1.215 8.31 1.355 ;
 RECT 8.08 1.955 8.36 2.21 ;
 RECT 8.1 0.87 8.38 1.01 ;
 RECT 7.995 1.355 8.135 1.815 ;
 RECT 6.515 0.83 6.655 1.145 ;
 RECT 6.92 1.285 7.06 1.525 ;
 RECT 6.895 1.67 7.035 1.99 ;
 RECT 6.515 1.145 7.06 1.285 ;
 RECT 6.45 1.99 7.035 2.13 ;
 RECT 6.885 1.525 7.115 1.67 ;
 RECT 11.405 0.96 11.75 1.1 ;
 RECT 11.405 0.625 11.545 0.96 ;
 RECT 11.405 0.365 11.545 0.485 ;
 RECT 10.3 0.485 11.545 0.625 ;
 RECT 11.61 1.1 11.75 2.16 ;
 RECT 10.3 0.42 10.445 0.485 ;
 RECT 10.3 0.625 10.445 0.67 ;
 RECT 12.365 0.365 12.505 1.075 ;
 RECT 11.405 0.225 12.505 0.365 ;
 RECT 12.745 1.005 12.885 1.075 ;
 RECT 12.745 1.215 12.885 1.285 ;
 RECT 12.365 1.075 12.885 1.215 ;
 RECT 10.175 0.815 10.315 0.855 ;
 RECT 10.175 0.995 10.315 2.105 ;
 RECT 10.175 0.855 11.265 0.995 ;
 RECT 11.125 1.24 11.4 1.38 ;
 RECT 11.125 0.995 11.265 1.24 ;
 END
END SDFFSSRX1

MACRO SDFFSSRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 15.04 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 15.04 2.96 ;
 RECT 6.645 2.28 6.895 2.8 ;
 RECT 9.005 2.635 9.265 2.8 ;
 RECT 12.595 1.51 12.735 2.8 ;
 RECT 0.94 1.98 1.08 2.8 ;
 RECT 14.11 1.51 14.25 2.8 ;
 RECT 11.12 1.955 11.26 2.8 ;
 RECT 6.045 1.95 6.185 2.8 ;
 RECT 4.13 1.965 4.27 2.8 ;
 RECT 2.845 1.96 2.985 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 15.04 0.08 ;
 RECT 6.62 0.08 6.92 0.26 ;
 RECT 10.875 0.08 11.13 0.285 ;
 RECT 0.835 0.08 1.135 0.265 ;
 RECT 12.59 0.08 12.865 0.33 ;
 RECT 4.13 0.08 4.27 0.655 ;
 RECT 14.16 0.08 14.3 0.9 ;
 RECT 3.165 0.08 3.305 0.775 ;
 RECT 8.94 0.08 9.08 0.58 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.255 1.475 6.64 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.08 2.085 12.455 2.39 ;
 RECT 12.01 0.76 12.29 0.9 ;
 RECT 13.04 0.76 13.335 0.9 ;
 RECT 12.08 2.39 12.22 2.575 ;
 RECT 13.125 1.18 13.265 2.575 ;
 RECT 12.08 1.18 12.22 2.085 ;
 RECT 12.08 1.04 13.265 1.18 ;
 RECT 12.08 0.9 12.22 1.04 ;
 RECT 13.125 0.9 13.265 1.04 ;
 RECT 13.125 0.755 13.265 0.76 ;
 END
 ANTENNADIFFAREA 1.007 ;
 END QN

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.55 1.46 1.93 1.74 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.655 1.485 0.97 1.745 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SETB

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.91 1.125 3.285 1.445 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END RSTB

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.515 0.22 3.99 0.635 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4 1.145 4.535 1.445 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.64 1.43 14.78 2.575 ;
 RECT 13.64 1.18 13.78 2.575 ;
 RECT 13.64 1.04 14.78 1.18 ;
 RECT 13.64 0.615 13.78 1.04 ;
 RECT 14.415 1.18 14.78 1.43 ;
 RECT 14.64 0.47 14.78 1.04 ;
 END
 ANTENNADIFFAREA 0.999 ;
 END Q

 OBS
 LAYER PO ;
 RECT 7.025 1.735 7.125 2.685 ;
 RECT 7.09 1.255 7.19 1.49 ;
 RECT 7.955 0.47 8.245 0.705 ;
 RECT 7.955 0.705 8.055 1.155 ;
 RECT 8.725 1.78 8.825 2.685 ;
 RECT 7.09 0.685 7.19 1.155 ;
 RECT 6.88 1.62 7.125 1.735 ;
 RECT 7.025 2.685 8.825 2.785 ;
 RECT 7.09 1.155 8.055 1.255 ;
 RECT 9.935 1.505 10.035 2.27 ;
 RECT 9.935 2.27 10.455 2.51 ;
 RECT 1.665 0.75 1.765 1.48 ;
 RECT 1.665 1.715 1.765 2.47 ;
 RECT 1.62 1.48 1.85 1.715 ;
 RECT 11.145 1.325 13.01 1.365 ;
 RECT 11.145 1.365 12.07 1.44 ;
 RECT 11.145 1.205 12.435 1.325 ;
 RECT 11.575 1.135 12.435 1.205 ;
 RECT 12.335 1.425 12.435 2.79 ;
 RECT 12.335 1.365 13.01 1.425 ;
 RECT 11.185 0.5 11.285 1.205 ;
 RECT 11.395 1.44 11.495 2.695 ;
 RECT 12.335 0.195 12.435 1.135 ;
 RECT 12.91 0.195 13.01 1.325 ;
 RECT 12.91 1.425 13.01 2.79 ;
 RECT 2.135 0.75 2.235 1.285 ;
 RECT 2.135 1.285 2.645 1.52 ;
 RECT 0.725 0.485 0.825 1.49 ;
 RECT 0.725 1.725 0.825 2.47 ;
 RECT 0.69 1.49 0.92 1.725 ;
 RECT 7.41 0.185 8.825 0.285 ;
 RECT 7.41 0.285 7.51 0.525 ;
 RECT 8.725 0.285 8.825 1.26 ;
 RECT 7.37 0.525 7.6 0.76 ;
 RECT 10.255 0.445 10.53 0.655 ;
 RECT 10.43 0.655 10.53 2.09 ;
 RECT 3.705 0.22 5.045 0.32 ;
 RECT 3.705 0.32 4.015 0.455 ;
 RECT 4.945 0.32 5.045 1.4 ;
 RECT 5.415 1.5 5.515 2.4 ;
 RECT 3.915 0.455 4.015 2.39 ;
 RECT 4.94 1.4 5.53 1.5 ;
 RECT 4.475 0.645 4.575 1.16 ;
 RECT 4.475 1.395 4.575 2.39 ;
 RECT 4.225 1.16 4.575 1.395 ;
 RECT 5.415 0.415 5.515 1.22 ;
 RECT 5.34 0.18 5.57 0.415 ;
 RECT 4.945 1.69 5.045 2.57 ;
 RECT 3.4 2.57 5.045 2.67 ;
 RECT 3.4 1.97 3.63 2.57 ;
 RECT 6.485 1.3 6.585 1.48 ;
 RECT 6.485 1.2 6.87 1.3 ;
 RECT 6.77 0.64 6.87 1.2 ;
 RECT 6.3 1.72 6.4 2.37 ;
 RECT 6.3 1.48 6.595 1.72 ;
 RECT 13.895 0.29 13.995 1.325 ;
 RECT 13.895 1.325 14.525 1.425 ;
 RECT 13.895 1.425 13.995 2.79 ;
 RECT 13.255 0.29 13.49 0.45 ;
 RECT 13.255 0.195 13.995 0.29 ;
 RECT 13.255 0.19 13.99 0.195 ;
 RECT 14.425 0.26 14.525 1.325 ;
 RECT 14.425 1.425 14.525 2.79 ;
 RECT 2.83 0.57 2.93 1.19 ;
 RECT 1.195 0.57 1.295 1.33 ;
 RECT 2.83 1.425 2.93 1.715 ;
 RECT 2.135 1.815 2.235 2.47 ;
 RECT 2.83 1.19 3.235 1.425 ;
 RECT 1.195 0.47 2.93 0.57 ;
 RECT 2.135 1.715 2.93 1.815 ;
 RECT 1.195 1.78 1.295 2.68 ;
 RECT 0.28 2.38 0.51 2.68 ;
 RECT 0.28 2.68 1.295 2.78 ;
 RECT 7.91 1.675 8.01 2.495 ;
 RECT 7.385 1.49 7.63 1.575 ;
 RECT 7.385 1.575 8.01 1.675 ;
 RECT 7.385 1.675 7.63 1.735 ;
 RECT 10.73 0.265 10.83 1.16 ;
 RECT 9.165 0.265 9.505 0.435 ;
 RECT 9.165 0.165 10.83 0.265 ;
 RECT 10.73 1.16 10.965 1.37 ;
 RECT 10.905 1.64 11.005 2.69 ;
 RECT 9.53 2.385 9.75 2.69 ;
 RECT 9.53 2.69 11.005 2.79 ;
 RECT 9.96 0.685 10.06 1.255 ;
 RECT 9.825 0.455 10.06 0.685 ;
 RECT 9.165 0.66 9.265 1.59 ;
 RECT 9.165 1.82 9.265 2.49 ;
 RECT 9.115 1.59 9.355 1.82 ;
 RECT 8.425 0.65 8.525 1.48 ;
 RECT 8.405 1.715 8.505 2.475 ;
 RECT 8.325 1.48 8.555 1.715 ;
 RECT 6.88 1.49 7.19 1.62 ;
 LAYER CO ;
 RECT 5.635 2 5.765 2.13 ;
 RECT 3.055 1.245 3.185 1.375 ;
 RECT 3.665 0.87 3.795 1 ;
 RECT 3.575 1.69 3.705 1.82 ;
 RECT 4.135 0.44 4.265 0.57 ;
 RECT 4.135 2.035 4.265 2.165 ;
 RECT 4.695 0.87 4.825 1 ;
 RECT 4.695 2 4.825 2.13 ;
 RECT 5.165 0.87 5.295 1 ;
 RECT 5.165 2 5.295 2.13 ;
 RECT 5.635 0.87 5.765 1 ;
 RECT 1.885 0.975 2.015 1.105 ;
 RECT 0.33 2.435 0.46 2.565 ;
 RECT 0.945 2.055 1.075 2.185 ;
 RECT 1.415 2.055 1.545 2.185 ;
 RECT 2.465 1.34 2.595 1.47 ;
 RECT 0.955 0.13 1.085 0.26 ;
 RECT 0.74 1.545 0.87 1.675 ;
 RECT 2.355 2.055 2.485 2.185 ;
 RECT 2.355 0.975 2.485 1.105 ;
 RECT 1.885 2.055 2.015 2.185 ;
 RECT 1.415 0.975 1.545 1.105 ;
 RECT 0.475 2.055 0.605 2.185 ;
 RECT 0.475 0.705 0.605 0.835 ;
 RECT 6.52 0.905 6.65 1.035 ;
 RECT 6.05 2 6.18 2.13 ;
 RECT 1.67 1.535 1.8 1.665 ;
 RECT 13.13 1.59 13.26 1.72 ;
 RECT 12.6 1.59 12.73 1.72 ;
 RECT 12.6 1.85 12.73 1.98 ;
 RECT 12.6 2.115 12.73 2.245 ;
 RECT 12.6 2.375 12.73 2.505 ;
 RECT 10.285 2.33 10.415 2.46 ;
 RECT 10.78 1.2 10.91 1.33 ;
 RECT 13.13 1.85 13.26 1.98 ;
 RECT 13.13 2.115 13.26 2.245 ;
 RECT 13.13 2.375 13.26 2.505 ;
 RECT 11.2 1.25 11.33 1.38 ;
 RECT 12.085 1.59 12.215 1.72 ;
 RECT 12.085 1.85 12.215 1.98 ;
 RECT 6.935 1.535 7.065 1.665 ;
 RECT 3.17 0.59 3.3 0.72 ;
 RECT 3.17 0.33 3.3 0.46 ;
 RECT 10.95 0.15 11.08 0.28 ;
 RECT 8.945 0.38 9.075 0.51 ;
 RECT 9.58 2.435 9.71 2.565 ;
 RECT 9.585 1.755 9.715 1.885 ;
 RECT 10.305 0.485 10.435 0.615 ;
 RECT 11.41 0.87 11.54 1 ;
 RECT 11.125 2.01 11.255 2.14 ;
 RECT 11.615 1.965 11.745 2.095 ;
 RECT 9.17 1.63 9.3 1.76 ;
 RECT 8.375 1.53 8.505 1.66 ;
 RECT 14.115 1.59 14.245 1.72 ;
 RECT 14.115 1.85 14.245 1.98 ;
 RECT 14.115 2.115 14.245 2.245 ;
 RECT 14.165 0.6 14.295 0.73 ;
 RECT 9.055 2.64 9.185 2.77 ;
 RECT 6.715 2.385 6.845 2.515 ;
 RECT 13.645 2.115 13.775 2.245 ;
 RECT 13.645 1.59 13.775 1.72 ;
 RECT 13.645 2.375 13.775 2.505 ;
 RECT 13.645 0.765 13.775 0.895 ;
 RECT 14.645 1.85 14.775 1.98 ;
 RECT 8.065 0.525 8.195 0.655 ;
 RECT 9.315 0.255 9.445 0.385 ;
 RECT 2.85 2.345 2.98 2.475 ;
 RECT 2.85 2.085 2.98 2.215 ;
 RECT 7.245 1.825 7.375 1.955 ;
 RECT 7.42 0.58 7.55 0.71 ;
 RECT 12.65 0.15 12.78 0.28 ;
 RECT 12.085 2.115 12.215 2.245 ;
 RECT 12.085 2.375 12.215 2.505 ;
 RECT 12.085 0.765 12.215 0.895 ;
 RECT 13.13 0.765 13.26 0.895 ;
 RECT 13.305 0.28 13.435 0.41 ;
 RECT 10.18 1.9 10.31 2.03 ;
 RECT 10.18 0.87 10.31 1 ;
 RECT 9.875 0.505 10.005 0.635 ;
 RECT 14.115 2.375 14.245 2.505 ;
 RECT 4.32 1.215 4.45 1.345 ;
 RECT 5.39 0.235 5.52 0.365 ;
 RECT 3.46 2.03 3.59 2.16 ;
 RECT 9.585 0.88 9.715 1.01 ;
 RECT 9.585 2.015 9.715 2.145 ;
 RECT 6.74 0.125 6.87 0.255 ;
 RECT 8.155 2.07 8.285 2.2 ;
 RECT 8.175 0.88 8.305 1.01 ;
 RECT 7.66 2.105 7.79 2.235 ;
 RECT 7.705 0.88 7.835 1.01 ;
 RECT 7.44 1.535 7.57 1.665 ;
 RECT 7.31 0.905 7.44 1.035 ;
 RECT 6.425 1.535 6.555 1.665 ;
 RECT 6.52 2 6.65 2.13 ;
 RECT 13.645 1.85 13.775 1.98 ;
 RECT 14.645 2.115 14.775 2.245 ;
 RECT 14.645 2.375 14.775 2.505 ;
 RECT 14.645 1.59 14.775 1.72 ;
 RECT 14.645 0.625 14.775 0.755 ;
 RECT 3.775 0.26 3.905 0.39 ;
 LAYER M1 ;
 RECT 3.57 1.005 3.71 1.965 ;
 RECT 3.455 1.965 3.71 2.265 ;
 RECT 3.57 0.865 4.55 1.005 ;
 RECT 4.41 0.37 4.55 0.865 ;
 RECT 4.41 0.23 5.6 0.37 ;
 RECT 4.69 0.795 4.83 2.18 ;
 RECT 1.41 2.47 2.49 2.61 ;
 RECT 2.35 1.985 2.49 2.47 ;
 RECT 1.41 1.985 1.55 2.47 ;
 RECT 0.325 0.545 0.465 0.7 ;
 RECT 0.325 0.84 0.465 2.05 ;
 RECT 0.325 2.19 0.465 2.635 ;
 RECT 0.325 2.05 0.665 2.19 ;
 RECT 0.325 0.7 0.675 0.84 ;
 RECT 2.35 1.335 2.77 1.475 ;
 RECT 2.63 0.545 2.77 1.335 ;
 RECT 0.325 0.405 2.77 0.545 ;
 RECT 2.07 1.11 2.21 1.675 ;
 RECT 2.07 1.815 2.21 1.905 ;
 RECT 1.88 2.045 2.02 2.26 ;
 RECT 1.805 0.97 2.21 1.11 ;
 RECT 1.88 1.905 2.21 2.045 ;
 RECT 2.07 1.675 3.3 1.815 ;
 RECT 3.85 1.825 3.99 2.52 ;
 RECT 3.16 1.815 3.3 2.52 ;
 RECT 3.16 2.52 3.99 2.66 ;
 RECT 4.41 1.825 4.55 2.32 ;
 RECT 5.63 0.79 5.77 2.32 ;
 RECT 3.85 1.685 4.55 1.825 ;
 RECT 4.41 2.32 5.77 2.46 ;
 RECT 1.41 0.83 1.55 0.97 ;
 RECT 1.41 0.69 2.49 0.83 ;
 RECT 2.35 0.83 2.49 1.165 ;
 RECT 1.335 0.97 1.62 1.11 ;
 RECT 10.585 1.195 10.98 1.335 ;
 RECT 10.585 1.335 10.725 2.325 ;
 RECT 10.195 2.325 10.725 2.465 ;
 RECT 7.99 0.52 8.8 0.66 ;
 RECT 8.66 0.66 8.8 0.79 ;
 RECT 8.66 0.79 9.36 0.93 ;
 RECT 9.22 0.25 9.515 0.39 ;
 RECT 9.22 0.39 9.36 0.79 ;
 RECT 9.58 0.81 9.72 1.185 ;
 RECT 9.58 1.325 9.72 2.215 ;
 RECT 8.795 1.185 9.72 1.325 ;
 RECT 8.275 1.525 8.935 1.66 ;
 RECT 8.76 1.52 8.935 1.525 ;
 RECT 8.275 1.66 8.93 1.665 ;
 RECT 8.795 1.325 8.935 1.52 ;
 RECT 8.08 1.96 8.36 2.215 ;
 RECT 8.17 1.015 8.31 1.22 ;
 RECT 7.995 1.22 8.31 1.36 ;
 RECT 7.995 1.82 9.305 1.96 ;
 RECT 9.165 1.56 9.305 1.82 ;
 RECT 8.1 0.875 8.38 1.015 ;
 RECT 7.995 1.36 8.135 1.82 ;
 RECT 7.175 1.82 7.495 1.96 ;
 RECT 7.355 1.96 7.495 2.51 ;
 RECT 7.355 2.51 8.57 2.65 ;
 RECT 7.305 1.715 7.495 1.82 ;
 RECT 8.43 2.495 8.57 2.51 ;
 RECT 7.415 0.5 7.555 0.84 ;
 RECT 7.305 0.84 7.555 1.035 ;
 RECT 7.305 1.035 7.445 1.485 ;
 RECT 7.305 1.485 7.575 1.715 ;
 RECT 9.405 2.495 10.01 2.57 ;
 RECT 8.43 2.355 9.545 2.43 ;
 RECT 8.43 2.43 10.01 2.495 ;
 RECT 9.87 0.45 10.01 2.43 ;
 RECT 5.155 0.65 5.3 0.675 ;
 RECT 5.16 0.675 5.3 2.18 ;
 RECT 7.7 0.36 7.84 0.8 ;
 RECT 5.155 0.51 7.22 0.65 ;
 RECT 7.08 0.36 7.22 0.51 ;
 RECT 7.08 0.22 7.84 0.36 ;
 RECT 7.7 0.8 7.855 1.095 ;
 RECT 7.715 1.095 7.855 2.035 ;
 RECT 7.655 2.035 7.855 2.305 ;
 RECT 6.515 0.835 6.655 1.15 ;
 RECT 6.92 1.29 7.06 1.53 ;
 RECT 6.895 1.675 7.035 1.995 ;
 RECT 6.515 1.15 7.06 1.29 ;
 RECT 6.45 1.995 7.035 2.135 ;
 RECT 6.885 1.53 7.115 1.675 ;
 RECT 11.405 0.965 11.75 1.105 ;
 RECT 11.405 0.615 11.545 0.965 ;
 RECT 11.61 1.105 11.75 2.165 ;
 RECT 10.3 0.425 10.445 0.475 ;
 RECT 10.3 0.615 10.445 0.675 ;
 RECT 10.3 0.475 13.335 0.615 ;
 RECT 13.195 0.22 13.445 0.47 ;
 RECT 13.195 0.47 13.335 0.475 ;
 RECT 10.175 0.82 10.315 0.86 ;
 RECT 10.175 1 10.315 2.11 ;
 RECT 10.175 0.86 11.265 1 ;
 RECT 11.125 1.245 11.4 1.385 ;
 RECT 11.125 1 11.265 1.245 ;
 END
END SDFFSSRX2

MACRO SDFFX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.56 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.56 2.96 ;
 RECT 6.195 2.635 6.455 2.8 ;
 RECT 1.27 2.005 1.41 2.8 ;
 RECT 3.835 2.38 4.085 2.8 ;
 RECT 3.18 1.98 3.32 2.8 ;
 RECT 8.31 1.955 8.45 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 9.785 1.51 9.925 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.56 0.08 ;
 RECT 3.81 0.08 4.11 0.26 ;
 RECT 8.065 0.08 8.32 0.285 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 1.055 ;
 RECT 6.13 0.08 6.27 0.58 ;
 RECT 9.835 0.08 9.975 0.815 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.49 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.595 2.075 2.015 2.45 ;
 RECT 2.575 1.86 2.715 1.89 ;
 RECT 1.875 1.72 2.715 1.86 ;
 RECT 2.575 1.615 2.715 1.72 ;
 RECT 1.875 1.86 2.015 2.075 ;
 RECT 1.875 1.11 2.015 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.225 1.16 2.58 1.455 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.27 2.085 9.56 2.39 ;
 RECT 9.27 2.39 9.41 2.575 ;
 RECT 9.27 0.56 9.41 2.085 ;
 END
 ANTENNADIFFAREA 0.527 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.085 2.08 10.49 2.385 ;
 RECT 10.315 2.385 10.455 2.575 ;
 RECT 10.315 0.61 10.455 2.08 ;
 END
 ANTENNADIFFAREA 0.467 ;
 END Q

 OBS
 LAYER PO ;
 RECT 7.125 2.27 7.645 2.51 ;
 RECT 6.595 0.165 8.02 0.205 ;
 RECT 6.355 0.205 8.02 0.265 ;
 RECT 6.355 0.265 6.695 0.435 ;
 RECT 7.92 0.265 8.02 1.16 ;
 RECT 7.92 1.16 8.155 1.37 ;
 RECT 10.1 0.27 10.2 1.035 ;
 RECT 10.1 1.27 10.2 2.79 ;
 RECT 9.9 1.035 10.2 1.27 ;
 RECT 2.245 1.455 2.345 1.645 ;
 RECT 2.665 0.655 2.765 1.245 ;
 RECT 2.245 1.225 2.465 1.245 ;
 RECT 2.245 1.345 2.465 1.455 ;
 RECT 2.195 1.745 2.295 2.67 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.245 1.245 2.765 1.345 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 2.665 1.865 2.765 2.48 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 4.07 1.49 4.38 1.62 ;
 RECT 4.28 1.255 4.38 1.49 ;
 RECT 4.215 1.735 4.315 2.685 ;
 RECT 5.915 1.78 6.015 2.685 ;
 RECT 4.07 1.62 4.315 1.735 ;
 RECT 5.145 0.705 5.245 1.155 ;
 RECT 4.28 0.685 4.38 1.155 ;
 RECT 5.145 0.47 5.435 0.705 ;
 RECT 4.215 2.685 6.015 2.785 ;
 RECT 4.28 1.155 5.245 1.255 ;
 RECT 4.6 0.185 6.015 0.285 ;
 RECT 4.6 0.285 4.7 0.525 ;
 RECT 5.915 0.285 6.015 1.26 ;
 RECT 4.56 0.525 4.79 0.76 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 5.1 1.675 5.2 2.495 ;
 RECT 4.575 1.49 4.82 1.575 ;
 RECT 4.575 1.675 4.82 1.735 ;
 RECT 4.575 1.575 5.2 1.675 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 8.585 1.44 8.685 2.51 ;
 RECT 8.335 1.205 9.625 1.365 ;
 RECT 9.525 1.365 9.625 2.79 ;
 RECT 8.375 0.65 8.475 1.205 ;
 RECT 8.335 1.365 9.26 1.44 ;
 RECT 9.525 0.195 9.625 1.135 ;
 RECT 8.765 1.135 9.625 1.205 ;
 RECT 8.095 1.64 8.195 2.69 ;
 RECT 6.72 2.385 6.94 2.69 ;
 RECT 6.72 2.69 8.195 2.79 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.245 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 7.445 0.445 7.72 0.655 ;
 RECT 7.62 0.655 7.72 2.09 ;
 RECT 7.15 0.685 7.25 1.255 ;
 RECT 7.015 0.455 7.25 0.685 ;
 RECT 5.595 1.33 5.715 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.48 1.475 5.715 1.71 ;
 RECT 5.615 0.65 5.715 1.33 ;
 RECT 6.355 0.66 6.455 1.59 ;
 RECT 6.355 1.82 6.455 2.49 ;
 RECT 6.305 1.59 6.545 1.82 ;
 RECT 7.125 1.465 7.225 2.27 ;
 LAYER CO ;
 RECT 3.295 1.535 3.425 1.665 ;
 RECT 3.71 1.995 3.84 2.125 ;
 RECT 7.065 0.505 7.195 0.635 ;
 RECT 7.495 0.485 7.625 0.615 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 9.94 1.085 10.07 1.215 ;
 RECT 10.32 0.68 10.45 0.81 ;
 RECT 9.84 0.615 9.97 0.745 ;
 RECT 3.905 2.385 4.035 2.515 ;
 RECT 9.275 0.63 9.405 0.76 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 8.14 0.15 8.27 0.28 ;
 RECT 10.32 2.115 10.45 2.245 ;
 RECT 10.32 2.375 10.45 2.505 ;
 RECT 10.32 1.59 10.45 1.72 ;
 RECT 9.79 2.375 9.92 2.505 ;
 RECT 9.275 1.59 9.405 1.72 ;
 RECT 9.275 1.85 9.405 1.98 ;
 RECT 4.125 1.535 4.255 1.665 ;
 RECT 5.255 0.525 5.385 0.655 ;
 RECT 6.36 1.63 6.49 1.76 ;
 RECT 5.53 1.525 5.66 1.655 ;
 RECT 6.775 0.88 6.905 1.01 ;
 RECT 6.245 2.64 6.375 2.77 ;
 RECT 2.285 1.275 2.415 1.405 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 4.435 1.825 4.565 1.955 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 4.63 1.535 4.76 1.665 ;
 RECT 6.135 0.38 6.265 0.51 ;
 RECT 7.37 1.9 7.5 2.03 ;
 RECT 7.37 0.87 7.5 1 ;
 RECT 9.79 1.59 9.92 1.72 ;
 RECT 9.79 1.85 9.92 1.98 ;
 RECT 9.79 2.115 9.92 2.245 ;
 RECT 8.6 0.87 8.73 1 ;
 RECT 8.315 2.01 8.445 2.14 ;
 RECT 8.805 1.965 8.935 2.095 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 0.805 0.875 0.935 1.005 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 9.275 2.115 9.405 2.245 ;
 RECT 9.275 2.375 9.405 2.505 ;
 RECT 7.475 2.33 7.605 2.46 ;
 RECT 7.97 1.2 8.1 1.33 ;
 RECT 10.32 1.85 10.45 1.98 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 6.505 0.255 6.635 0.385 ;
 RECT 8.39 1.25 8.52 1.38 ;
 RECT 6.775 2.015 6.905 2.145 ;
 RECT 3.93 0.125 4.06 0.255 ;
 RECT 4.61 0.58 4.74 0.71 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 6.77 2.435 6.9 2.565 ;
 RECT 6.775 1.755 6.905 1.885 ;
 LAYER M1 ;
 RECT 5.465 1.52 6.125 1.66 ;
 RECT 5.985 1.185 6.91 1.325 ;
 RECT 6.77 0.81 6.91 1.185 ;
 RECT 6.77 1.325 6.91 2.215 ;
 RECT 5.985 1.325 6.125 1.52 ;
 RECT 5.18 0.52 5.99 0.66 ;
 RECT 5.85 0.66 5.99 0.79 ;
 RECT 5.85 0.79 6.55 0.93 ;
 RECT 6.41 0.25 6.705 0.39 ;
 RECT 6.41 0.39 6.55 0.79 ;
 RECT 7.775 1.195 8.17 1.335 ;
 RECT 7.775 1.335 7.915 2.325 ;
 RECT 7.385 2.325 7.915 2.465 ;
 RECT 7.365 0.82 7.505 0.86 ;
 RECT 7.365 1 7.505 2.11 ;
 RECT 7.365 0.86 8.455 1 ;
 RECT 8.315 1.245 8.59 1.385 ;
 RECT 8.315 1 8.455 1.245 ;
 RECT 4.365 1.82 4.685 1.96 ;
 RECT 4.545 1.96 4.685 2.51 ;
 RECT 4.545 2.51 5.76 2.65 ;
 RECT 4.495 1.715 4.685 1.82 ;
 RECT 5.62 2.495 5.76 2.51 ;
 RECT 4.605 0.5 4.745 0.84 ;
 RECT 4.495 0.84 4.745 1.035 ;
 RECT 4.495 1.035 4.635 1.485 ;
 RECT 4.495 1.485 4.765 1.715 ;
 RECT 5.62 2.355 6.735 2.43 ;
 RECT 5.62 2.43 7.2 2.495 ;
 RECT 6.595 2.495 7.2 2.57 ;
 RECT 7.06 0.45 7.2 2.43 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.365 2.11 2.995 2.25 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 3.46 0.53 4.41 0.67 ;
 RECT 4.89 0.36 5.03 0.8 ;
 RECT 4.27 0.36 4.41 0.53 ;
 RECT 4.27 0.22 5.03 0.36 ;
 RECT 4.89 0.8 5.045 1.095 ;
 RECT 4.905 1.095 5.045 2.035 ;
 RECT 4.845 2.035 5.045 2.305 ;
 RECT 8.595 0.965 8.94 1.105 ;
 RECT 8.595 0.63 8.735 0.965 ;
 RECT 8.595 0.36 8.735 0.49 ;
 RECT 7.49 0.49 8.735 0.63 ;
 RECT 8.8 1.105 8.94 2.165 ;
 RECT 9.555 0.36 9.695 1.08 ;
 RECT 8.595 0.22 9.695 0.36 ;
 RECT 7.49 0.425 7.635 0.49 ;
 RECT 7.49 0.63 7.635 0.675 ;
 RECT 9.935 1.01 10.075 1.08 ;
 RECT 9.935 1.22 10.075 1.29 ;
 RECT 9.555 1.08 10.075 1.22 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.705 1.475 3.925 1.53 ;
 RECT 3.705 1.53 4.325 1.67 ;
 RECT 3.705 1.67 3.845 2.175 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 5.36 1.015 5.5 1.22 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 5.185 1.82 6.495 1.96 ;
 RECT 6.355 1.56 6.495 1.82 ;
 RECT 5.29 0.875 5.57 1.015 ;
 RECT 5.185 1.36 5.325 1.82 ;
 END
END SDFFX1

MACRO SDFFX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 11.52 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 11.52 2.96 ;
 RECT 3.835 2.38 4.085 2.8 ;
 RECT 1.27 2.005 1.41 2.8 ;
 RECT 6.195 2.635 6.455 2.8 ;
 RECT 9.26 1.515 9.4 2.8 ;
 RECT 10.315 1.51 10.455 2.8 ;
 RECT 11.255 1.51 11.395 2.8 ;
 RECT 3.18 1.98 3.32 2.8 ;
 RECT 8.31 1.955 8.45 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 11.52 0.08 ;
 RECT 3.18 0.08 3.32 1.055 ;
 RECT 8.065 0.08 8.32 0.285 ;
 RECT 10.245 0.08 10.5 0.245 ;
 RECT 3.81 0.08 4.11 0.26 ;
 RECT 6.13 0.08 6.27 0.58 ;
 RECT 9.18 0.08 9.32 0.63 ;
 RECT 11.255 0.08 11.395 0.7 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.27 0.08 1.41 1.055 ;
 END
 END VSS

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.475 3.505 1.785 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.09 1.475 1.615 1.75 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.595 2.075 2.015 2.45 ;
 RECT 2.575 1.86 2.715 1.89 ;
 RECT 1.875 1.72 2.715 1.86 ;
 RECT 2.575 1.615 2.715 1.72 ;
 RECT 1.875 1.86 2.015 2.075 ;
 RECT 1.875 1.11 2.015 1.72 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.225 1.16 2.58 1.445 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.635 2.085 9.945 2.39 ;
 RECT 9.74 2.39 9.88 2.575 ;
 RECT 9.74 0.72 9.88 2.085 ;
 END
 ANTENNADIFFAREA 0.788 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.785 2.39 10.925 2.575 ;
 RECT 10.6 2.085 10.925 2.39 ;
 RECT 10.785 0.72 10.925 2.085 ;
 END
 ANTENNADIFFAREA 0.622 ;
 END Q

 OBS
 LAYER PO ;
 RECT 2.965 0.405 3.065 2.465 ;
 RECT 2.76 0.175 3.065 0.405 ;
 RECT 1.86 0.64 1.96 1.145 ;
 RECT 1.82 1.145 2.065 1.385 ;
 RECT 2.665 1.865 2.765 2.48 ;
 RECT 2.525 1.635 2.765 1.865 ;
 RECT 10.57 0.2 10.67 1.035 ;
 RECT 10.46 1.035 10.67 1.2 ;
 RECT 10.57 1.3 10.67 2.79 ;
 RECT 11.04 0.2 11.14 1.2 ;
 RECT 11.04 1.3 11.14 2.79 ;
 RECT 10.46 1.2 11.14 1.3 ;
 RECT 7.125 1.4 7.225 2.27 ;
 RECT 7.125 2.27 7.645 2.51 ;
 RECT 6.355 0.205 8.02 0.265 ;
 RECT 7.92 0.265 8.02 1.16 ;
 RECT 6.595 0.165 8.02 0.205 ;
 RECT 6.355 0.265 6.695 0.435 ;
 RECT 7.92 1.16 8.155 1.37 ;
 RECT 7.445 0.445 7.72 0.655 ;
 RECT 7.62 0.655 7.72 2.03 ;
 RECT 7.15 0.685 7.25 1.22 ;
 RECT 7.015 0.455 7.25 0.685 ;
 RECT 8.765 1.2 10.2 1.205 ;
 RECT 8.335 1.205 10.2 1.3 ;
 RECT 8.335 1.365 9.26 1.44 ;
 RECT 8.335 1.3 9.625 1.365 ;
 RECT 8.765 1.135 9.625 1.2 ;
 RECT 10.1 0.2 10.2 1.2 ;
 RECT 10.1 1.3 10.2 2.79 ;
 RECT 8.375 0.65 8.475 1.205 ;
 RECT 8.585 1.44 8.685 2.46 ;
 RECT 9.525 0.195 9.625 1.135 ;
 RECT 9.525 1.365 9.625 2.79 ;
 RECT 6.355 0.66 6.455 1.59 ;
 RECT 6.355 1.82 6.455 2.49 ;
 RECT 6.305 1.59 6.545 1.82 ;
 RECT 5.595 1.33 5.715 1.475 ;
 RECT 5.595 1.71 5.695 2.475 ;
 RECT 5.48 1.475 5.715 1.71 ;
 RECT 5.615 0.65 5.715 1.33 ;
 RECT 4.6 0.185 6.015 0.285 ;
 RECT 4.6 0.285 4.7 0.525 ;
 RECT 5.915 0.285 6.015 1.26 ;
 RECT 4.56 0.525 4.79 0.76 ;
 RECT 2.245 1.455 2.345 1.645 ;
 RECT 2.665 0.655 2.765 1.245 ;
 RECT 2.245 1.225 2.465 1.245 ;
 RECT 2.245 1.345 2.465 1.455 ;
 RECT 2.195 1.745 2.295 2.67 ;
 RECT 2.195 1.645 2.345 1.745 ;
 RECT 2.245 1.245 2.765 1.345 ;
 RECT 1.055 1.475 1.625 1.75 ;
 RECT 1.525 0.655 1.625 1.475 ;
 RECT 1.525 1.75 1.625 2.465 ;
 RECT 1.055 0.635 1.155 1.475 ;
 RECT 1.055 1.75 1.155 2.465 ;
 RECT 3.44 0.655 3.54 1.48 ;
 RECT 3.245 1.48 3.54 1.72 ;
 RECT 3.44 1.72 3.54 2.37 ;
 RECT 8.095 1.64 8.195 2.69 ;
 RECT 6.72 2.385 6.94 2.69 ;
 RECT 6.72 2.69 8.195 2.79 ;
 RECT 5.1 1.675 5.2 2.495 ;
 RECT 4.575 1.49 4.82 1.575 ;
 RECT 4.575 1.575 5.2 1.675 ;
 RECT 4.575 1.675 4.82 1.735 ;
 RECT 4.07 1.49 4.38 1.62 ;
 RECT 4.215 1.735 4.315 2.685 ;
 RECT 4.28 1.255 4.38 1.49 ;
 RECT 5.145 0.47 5.435 0.705 ;
 RECT 5.145 0.705 5.245 1.155 ;
 RECT 5.915 1.78 6.015 2.685 ;
 RECT 4.28 0.685 4.38 1.155 ;
 RECT 4.07 1.62 4.315 1.735 ;
 RECT 4.215 2.685 6.015 2.785 ;
 RECT 4.28 1.155 5.245 1.255 ;
 LAYER CO ;
 RECT 7.475 2.33 7.605 2.46 ;
 RECT 7.97 1.2 8.1 1.33 ;
 RECT 9.265 1.59 9.395 1.72 ;
 RECT 9.265 1.85 9.395 1.98 ;
 RECT 9.265 2.115 9.395 2.245 ;
 RECT 9.265 2.375 9.395 2.505 ;
 RECT 4.125 1.535 4.255 1.665 ;
 RECT 5.255 0.525 5.385 0.655 ;
 RECT 6.505 0.255 6.635 0.385 ;
 RECT 8.39 1.25 8.52 1.38 ;
 RECT 4.435 1.825 4.565 1.955 ;
 RECT 4.61 0.58 4.74 0.71 ;
 RECT 1.275 0.875 1.405 1.005 ;
 RECT 6.245 2.64 6.375 2.77 ;
 RECT 2.285 1.275 2.415 1.405 ;
 RECT 11.26 1.85 11.39 1.98 ;
 RECT 11.26 2.115 11.39 2.245 ;
 RECT 11.26 2.375 11.39 2.505 ;
 RECT 10.5 1.085 10.63 1.215 ;
 RECT 10.79 0.77 10.92 0.9 ;
 RECT 10.79 1.85 10.92 1.98 ;
 RECT 10.79 2.115 10.92 2.245 ;
 RECT 10.79 2.375 10.92 2.505 ;
 RECT 10.79 1.59 10.92 1.72 ;
 RECT 10.32 0.11 10.45 0.24 ;
 RECT 10.32 1.59 10.45 1.72 ;
 RECT 10.32 1.85 10.45 1.98 ;
 RECT 10.32 2.115 10.45 2.245 ;
 RECT 10.32 2.375 10.45 2.505 ;
 RECT 9.745 2.115 9.875 2.245 ;
 RECT 9.185 0.43 9.315 0.56 ;
 RECT 9.745 1.85 9.875 1.98 ;
 RECT 5.365 0.88 5.495 1.01 ;
 RECT 4.85 2.105 4.98 2.235 ;
 RECT 4.895 0.88 5.025 1.01 ;
 RECT 4.63 1.535 4.76 1.665 ;
 RECT 4.5 0.905 4.63 1.035 ;
 RECT 3.295 1.535 3.425 1.665 ;
 RECT 3.71 1.995 3.84 2.125 ;
 RECT 3.79 0.875 3.92 1.005 ;
 RECT 3.185 2.05 3.315 2.18 ;
 RECT 3.185 0.875 3.315 1.005 ;
 RECT 2.22 0.875 2.35 1.005 ;
 RECT 2.415 2.115 2.545 2.245 ;
 RECT 6.775 2.015 6.905 2.145 ;
 RECT 3.93 0.125 4.06 0.255 ;
 RECT 1.275 2.055 1.405 2.185 ;
 RECT 0.805 2.055 0.935 2.185 ;
 RECT 1.28 1.55 1.41 1.68 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 6.77 2.435 6.9 2.565 ;
 RECT 6.775 1.755 6.905 1.885 ;
 RECT 11.26 0.5 11.39 0.63 ;
 RECT 9.745 0.77 9.875 0.9 ;
 RECT 2.58 1.685 2.71 1.815 ;
 RECT 1.88 1.195 2.01 1.325 ;
 RECT 5.345 2.07 5.475 2.2 ;
 RECT 2.81 0.225 2.94 0.355 ;
 RECT 9.745 2.375 9.875 2.505 ;
 RECT 9.745 1.59 9.875 1.72 ;
 RECT 11.26 1.59 11.39 1.72 ;
 RECT 3.905 2.385 4.035 2.515 ;
 RECT 8.14 0.15 8.27 0.28 ;
 RECT 6.135 0.38 6.265 0.51 ;
 RECT 7.37 1.9 7.5 2.03 ;
 RECT 7.37 0.87 7.5 1 ;
 RECT 7.065 0.505 7.195 0.635 ;
 RECT 7.495 0.485 7.625 0.615 ;
 RECT 8.6 0.87 8.73 1 ;
 RECT 8.315 2.01 8.445 2.14 ;
 RECT 8.805 1.965 8.935 2.095 ;
 RECT 6.36 1.63 6.49 1.76 ;
 RECT 5.53 1.525 5.66 1.655 ;
 RECT 6.775 0.88 6.905 1.01 ;
 RECT 0.805 0.875 0.935 1.005 ;
 LAYER M1 ;
 RECT 7.775 1.195 8.17 1.335 ;
 RECT 7.775 1.335 7.915 2.325 ;
 RECT 7.385 2.325 7.915 2.465 ;
 RECT 6.77 0.81 6.91 1.185 ;
 RECT 6.77 1.325 6.91 2.215 ;
 RECT 5.985 1.185 6.91 1.325 ;
 RECT 5.465 1.52 6.125 1.66 ;
 RECT 5.985 1.325 6.125 1.52 ;
 RECT 5.18 0.52 5.99 0.66 ;
 RECT 5.85 0.66 5.99 0.79 ;
 RECT 5.85 0.79 6.55 0.93 ;
 RECT 6.41 0.25 6.705 0.39 ;
 RECT 6.41 0.39 6.55 0.79 ;
 RECT 8.595 0.965 9.6 1.105 ;
 RECT 9.46 0.535 9.6 0.965 ;
 RECT 8.595 0.63 8.735 0.965 ;
 RECT 7.49 0.49 8.735 0.63 ;
 RECT 8.8 1.105 8.94 2.165 ;
 RECT 7.49 0.425 7.635 0.49 ;
 RECT 7.49 0.63 7.635 0.675 ;
 RECT 10.385 0.535 10.525 1.01 ;
 RECT 9.46 0.395 10.525 0.535 ;
 RECT 10.385 1.01 10.635 1.29 ;
 RECT 4.365 1.82 4.685 1.96 ;
 RECT 4.545 1.96 4.685 2.51 ;
 RECT 4.545 2.51 5.76 2.65 ;
 RECT 4.495 1.715 4.685 1.82 ;
 RECT 5.62 2.495 5.76 2.51 ;
 RECT 4.605 0.5 4.745 0.84 ;
 RECT 4.495 0.84 4.745 1.035 ;
 RECT 4.495 1.035 4.635 1.485 ;
 RECT 4.495 1.485 4.765 1.715 ;
 RECT 6.595 2.495 7.2 2.57 ;
 RECT 5.62 2.355 6.735 2.43 ;
 RECT 5.62 2.43 7.2 2.495 ;
 RECT 7.06 0.45 7.2 2.43 ;
 RECT 2.855 1.01 2.995 1.195 ;
 RECT 2.855 1.335 2.995 2.11 ;
 RECT 2.155 0.87 2.995 1.01 ;
 RECT 2.365 2.11 2.995 2.25 ;
 RECT 2.855 1.195 3.6 1.335 ;
 RECT 3.46 0.67 3.6 1.195 ;
 RECT 3.46 0.53 4.41 0.67 ;
 RECT 4.89 0.36 5.03 0.8 ;
 RECT 4.27 0.36 4.41 0.53 ;
 RECT 4.27 0.22 5.03 0.36 ;
 RECT 4.89 0.8 5.045 1.095 ;
 RECT 4.905 1.095 5.045 2.035 ;
 RECT 4.845 2.035 5.045 2.305 ;
 RECT 5.185 1.82 6.495 1.96 ;
 RECT 5.36 1.015 5.5 1.22 ;
 RECT 5.185 1.22 5.5 1.36 ;
 RECT 6.355 1.56 6.495 1.82 ;
 RECT 5.27 1.96 5.55 2.215 ;
 RECT 5.29 0.875 5.57 1.015 ;
 RECT 5.185 1.36 5.325 1.82 ;
 RECT 0.8 0.8 0.94 1.195 ;
 RECT 0.8 1.335 0.94 2.305 ;
 RECT 1.585 0.36 1.725 1.195 ;
 RECT 0.8 1.195 1.725 1.335 ;
 RECT 1.585 0.22 3.01 0.36 ;
 RECT 7.365 0.82 7.505 0.86 ;
 RECT 7.365 1 7.505 2.11 ;
 RECT 7.365 0.86 8.455 1 ;
 RECT 8.315 1.245 8.59 1.385 ;
 RECT 8.315 1 8.455 1.245 ;
 RECT 3.785 0.825 3.925 1.475 ;
 RECT 3.705 1.475 3.925 1.53 ;
 RECT 3.705 1.53 4.325 1.67 ;
 RECT 3.705 1.67 3.845 2.175 ;
 END
END SDFFX2

MACRO AODFFARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8 BY 5.76 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8 2.96 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.945 1.475 2.27 1.835 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.8 0.505 1.06 0.775 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.92 4.32 7.16 4.64 ;
 RECT 5.07 4.985 5.21 5.4 ;
 RECT 4.235 4.845 5.21 4.985 ;
 RECT 4.165 5.35 4.44 5.49 ;
 RECT 7.01 4.64 7.15 5.4 ;
 RECT 7.01 3.11 7.42 3.25 ;
 RECT 7.01 3.25 7.15 4.32 ;
 RECT 4.235 4.985 4.375 5.35 ;
 RECT 5.07 5.4 7.15 5.54 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8 0.08 ;
 RECT 1.91 0.08 2.05 1.055 ;
 RECT 5.255 0.08 5.49 0.55 ;
 RECT 0.345 0.08 0.485 0.775 ;
 RECT 2.655 0.08 2.795 0.39 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 8 5.84 ;
 RECT 4.63 5.17 4.77 5.68 ;
 RECT 1.935 4.89 2.075 5.68 ;
 RECT 1.15 4.96 1.29 5.68 ;
 RECT 3.525 5.1 3.665 5.68 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.445 4.04 2.685 4.28 ;
 RECT 2.495 4.28 2.635 5.07 ;
 RECT 2.495 3.475 2.635 4.04 ;
 END
 ANTENNADIFFAREA 0.483 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.88 3.96 3.02 5.22 ;
 RECT 2.88 3.72 3.32 3.96 ;
 RECT 2.88 3.485 3.02 3.72 ;
 END
 ANTENNADIFFAREA 0.498 ;
 END QN

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.265 3.12 4.865 3.26 ;
 RECT 1.61 4.02 1.75 4.22 ;
 RECT 1.295 3.635 1.75 4.02 ;
 RECT 2.02 3.26 2.16 4.04 ;
 RECT 3.465 3.26 3.605 3.655 ;
 RECT 4.725 3.26 4.865 3.815 ;
 RECT 1.61 3.26 1.75 3.635 ;
 END
 END VDDG

 OBS
 LAYER PO ;
 RECT 3.29 1.595 3.535 1.69 ;
 RECT 6.495 2.67 6.595 3.085 ;
 RECT 4.98 3.185 5.08 4.195 ;
 RECT 4.98 3.085 6.595 3.185 ;
 RECT 5.32 3.06 5.54 3.085 ;
 RECT 5.32 3.185 5.54 3.3 ;
 RECT 6.375 2.43 6.595 2.67 ;
 RECT 4.765 0.695 4.865 1.61 ;
 RECT 4.8 1.71 4.9 2.345 ;
 RECT 4.765 1.61 4.9 1.71 ;
 RECT 4.645 0.465 4.885 0.695 ;
 RECT 5.93 1.61 6.195 1.74 ;
 RECT 6.095 1.74 6.195 2.31 ;
 RECT 5.905 0.635 6.005 1.51 ;
 RECT 5.905 1.51 6.195 1.61 ;
 RECT 0.81 0.52 1.055 0.54 ;
 RECT 0.81 0.64 1.055 0.77 ;
 RECT 1.695 0.64 1.795 2.465 ;
 RECT 0.81 0.54 1.795 0.64 ;
 RECT 7.18 2.415 7.4 3.305 ;
 RECT 2.17 0.655 2.27 1.495 ;
 RECT 1.975 1.495 2.27 1.745 ;
 RECT 2.17 1.745 2.27 2.37 ;
 RECT 5.065 0.285 5.165 1.24 ;
 RECT 3.33 0.185 5.165 0.285 ;
 RECT 3.33 0.285 3.43 0.51 ;
 RECT 3.29 0.51 3.535 0.755 ;
 RECT 3.01 1.265 3.11 1.52 ;
 RECT 2.51 1.52 3.11 1.62 ;
 RECT 2.945 1.62 3.045 2.68 ;
 RECT 5.625 1.61 5.725 2.68 ;
 RECT 2.51 1.44 2.755 1.52 ;
 RECT 2.51 1.62 2.755 1.69 ;
 RECT 3.875 0.705 3.975 1.165 ;
 RECT 3.01 0.585 3.11 1.165 ;
 RECT 3.875 0.47 4.16 0.705 ;
 RECT 2.945 2.68 5.725 2.78 ;
 RECT 3.01 1.165 3.975 1.265 ;
 RECT 2.275 2.98 2.375 4.44 ;
 RECT 2.275 4.675 2.375 5.455 ;
 RECT 2.18 4.44 2.39 4.675 ;
 RECT 3.135 2.98 3.235 4.49 ;
 RECT 3.135 4.72 3.235 5.635 ;
 RECT 3.135 4.49 3.6 4.72 ;
 RECT 4.365 0.65 4.465 1.215 ;
 RECT 4.325 1.45 4.425 2.345 ;
 RECT 4.325 1.215 4.555 1.45 ;
 RECT 5.77 4.54 5.87 5.075 ;
 RECT 5.715 5.075 5.945 5.305 ;
 RECT 1.02 2.475 1.51 3.315 ;
 RECT 6.375 1.32 7.68 1.42 ;
 RECT 7.58 1.42 7.68 3.76 ;
 RECT 6.6 3.76 7.68 3.86 ;
 RECT 6.6 3.86 6.82 4 ;
 RECT 6.375 1.205 6.595 1.32 ;
 RECT 6.375 1.42 6.595 1.445 ;
 RECT 5.815 3.465 5.915 4.225 ;
 RECT 5.815 4.225 6.45 4.325 ;
 RECT 4.905 4.45 5.005 5.505 ;
 RECT 4.905 5.505 6.45 5.605 ;
 RECT 6.35 4.325 6.45 5.505 ;
 RECT 6.85 2.5 6.95 3.365 ;
 RECT 5.815 3.365 6.95 3.465 ;
 RECT 6.78 2.26 7 2.5 ;
 RECT 4.49 3.07 4.59 3.82 ;
 RECT 4.345 3.82 4.59 4.06 ;
 RECT 4.49 4.06 4.59 5.12 ;
 RECT 3.89 3.07 3.99 4.45 ;
 RECT 4.19 4.55 4.29 5.3 ;
 RECT 3.89 4.45 4.29 4.55 ;
 RECT 4.19 5.3 4.42 5.54 ;
 RECT 5.3 3.485 5.4 4.38 ;
 RECT 5.3 4.59 5.4 5.125 ;
 RECT 5.185 4.38 5.42 4.59 ;
 RECT 3.83 1.595 3.93 2.35 ;
 RECT 3.29 1.445 3.535 1.495 ;
 RECT 3.29 1.495 3.93 1.595 ;
 LAYER CO ;
 RECT 5.375 1.95 5.505 2.08 ;
 RECT 1.335 3.125 1.465 3.255 ;
 RECT 1.155 5.015 1.285 5.145 ;
 RECT 1.155 5.275 1.285 5.405 ;
 RECT 6.645 3.81 6.775 3.94 ;
 RECT 6.42 1.26 6.55 1.39 ;
 RECT 6.42 2.48 6.55 2.61 ;
 RECT 2.5 4.89 2.63 5.02 ;
 RECT 2.885 3.845 3.015 3.975 ;
 RECT 5.025 1.63 5.155 1.76 ;
 RECT 4.545 1.95 4.675 2.08 ;
 RECT 2.57 1.495 2.7 1.625 ;
 RECT 4.39 3.875 4.52 4.005 ;
 RECT 2.885 5.025 3.015 5.155 ;
 RECT 6.1 4.77 6.23 4.9 ;
 RECT 4.075 1.925 4.205 2.055 ;
 RECT 4.095 0.88 4.225 1.01 ;
 RECT 3.58 1.94 3.71 2.07 ;
 RECT 3.625 0.88 3.755 1.01 ;
 RECT 3.345 1.49 3.475 1.62 ;
 RECT 3.23 0.905 3.36 1.035 ;
 RECT 2.025 3.58 2.155 3.71 ;
 RECT 2.5 4.075 2.63 4.205 ;
 RECT 1.445 0.875 1.575 1.005 ;
 RECT 1.445 2.115 1.575 2.245 ;
 RECT 0.87 0.575 1 0.705 ;
 RECT 3.42 4.54 3.55 4.67 ;
 RECT 1.94 4.96 2.07 5.09 ;
 RECT 3.47 3.45 3.6 3.58 ;
 RECT 3.53 5.155 3.66 5.285 ;
 RECT 2.22 4.495 2.35 4.625 ;
 RECT 0.35 0.59 0.48 0.72 ;
 RECT 0.35 0.33 0.48 0.46 ;
 RECT 4.7 0.515 4.83 0.645 ;
 RECT 5.305 0.41 5.435 0.54 ;
 RECT 2.655 2.345 2.785 2.475 ;
 RECT 2.39 1.995 2.52 2.125 ;
 RECT 2.52 0.875 2.65 1.005 ;
 RECT 1.915 2.05 2.045 2.18 ;
 RECT 1.915 0.875 2.045 1.005 ;
 RECT 7.225 3.115 7.355 3.245 ;
 RECT 7.225 2.465 7.355 2.595 ;
 RECT 6.825 2.31 6.955 2.44 ;
 RECT 2.035 1.55 2.165 1.68 ;
 RECT 3.345 0.555 3.475 0.685 ;
 RECT 3.165 1.825 3.295 1.955 ;
 RECT 3.98 0.525 4.11 0.655 ;
 RECT 4.24 5.355 4.37 5.485 ;
 RECT 2.885 4.105 3.015 4.235 ;
 RECT 5.765 5.125 5.895 5.255 ;
 RECT 2.885 3.555 3.015 3.685 ;
 RECT 5.36 3.115 5.49 3.245 ;
 RECT 1.615 4.025 1.745 4.155 ;
 RECT 1.615 3.765 1.745 3.895 ;
 RECT 1.615 3.505 1.745 3.635 ;
 RECT 6.1 3.825 6.23 3.955 ;
 RECT 4.73 3.63 4.86 3.76 ;
 RECT 5.52 4.77 5.65 4.9 ;
 RECT 4.09 3.81 4.22 3.94 ;
 RECT 5.985 1.55 6.115 1.68 ;
 RECT 4.375 1.26 4.505 1.39 ;
 RECT 6.32 0.88 6.45 1.01 ;
 RECT 6.315 1.84 6.445 1.97 ;
 RECT 2.66 0.21 2.79 0.34 ;
 RECT 6.045 2.465 6.175 2.595 ;
 RECT 3.94 4.77 4.07 4.9 ;
 RECT 5.52 3.765 5.65 3.895 ;
 RECT 5.24 4.42 5.37 4.55 ;
 RECT 2.5 3.55 2.63 3.68 ;
 RECT 1.335 2.525 1.465 2.655 ;
 RECT 4.635 5.24 4.765 5.37 ;
 RECT 2.025 3.84 2.155 3.97 ;
 RECT 2.5 3.81 2.63 3.94 ;
 RECT 2.025 3.32 2.155 3.45 ;
 LAYER M1 ;
 RECT 4.475 1.945 5.575 2.085 ;
 RECT 3.91 0.52 4.555 0.66 ;
 RECT 4.415 0.66 4.555 0.97 ;
 RECT 6.82 0.645 6.96 2.51 ;
 RECT 5.91 0.505 6.96 0.645 ;
 RECT 4.415 0.97 6.05 1.11 ;
 RECT 5.91 0.645 6.05 0.97 ;
 RECT 4.695 0.445 4.835 0.69 ;
 RECT 5.63 0.22 7.36 0.36 ;
 RECT 7.22 0.36 7.36 2.66 ;
 RECT 5.63 0.36 5.77 0.69 ;
 RECT 4.695 0.69 5.77 0.83 ;
 RECT 6.31 1.015 6.45 1.255 ;
 RECT 6.31 1.395 6.45 2.035 ;
 RECT 4.325 1.255 6.62 1.395 ;
 RECT 6.25 0.875 6.52 1.015 ;
 RECT 5.805 3.25 5.945 5.12 ;
 RECT 5.295 3.11 5.945 3.25 ;
 RECT 5.695 5.12 5.96 5.26 ;
 RECT 4.085 3.74 4.225 4.235 ;
 RECT 3.935 4.375 4.075 4.815 ;
 RECT 3.245 4.815 4.075 4.955 ;
 RECT 2.215 4.42 2.355 5.4 ;
 RECT 2.215 5.4 3.385 5.54 ;
 RECT 3.245 4.955 3.385 5.4 ;
 RECT 3.935 4.235 5.375 4.375 ;
 RECT 5.235 4.375 5.375 4.6 ;
 RECT 1.2 1.195 2.33 1.335 ;
 RECT 2.19 0.67 2.33 1.195 ;
 RECT 1.2 1.01 1.34 1.195 ;
 RECT 1.2 1.335 1.34 2.11 ;
 RECT 1.2 2.11 1.645 2.25 ;
 RECT 1.2 2.25 1.34 2.255 ;
 RECT 1.2 0.875 1.645 1.01 ;
 RECT 1.22 0.87 1.645 0.875 ;
 RECT 3.62 0.36 3.76 1.935 ;
 RECT 2.19 0.53 3.075 0.67 ;
 RECT 2.935 0.22 3.76 0.36 ;
 RECT 2.935 0.36 3.075 0.53 ;
 RECT 3.51 1.935 3.78 2.075 ;
 RECT 3.225 0.5 3.48 0.965 ;
 RECT 3.225 1.96 3.365 2.225 ;
 RECT 3.225 1.67 3.365 1.82 ;
 RECT 3.225 0.965 3.365 1.44 ;
 RECT 3.225 1.44 3.48 1.67 ;
 RECT 3.095 1.82 3.365 1.96 ;
 RECT 3.225 2.225 6.555 2.32 ;
 RECT 6.415 2.32 6.555 2.66 ;
 RECT 5.715 2.18 6.555 2.225 ;
 RECT 3.225 2.32 5.855 2.365 ;
 RECT 3.745 3.55 3.885 3.85 ;
 RECT 3.59 3.99 3.73 4.535 ;
 RECT 3.35 4.535 3.73 4.675 ;
 RECT 3.59 3.85 3.885 3.99 ;
 RECT 3.745 3.41 4.525 3.55 ;
 RECT 4.385 3.55 4.525 3.955 ;
 RECT 4.385 3.955 5.655 4.095 ;
 RECT 5.515 3.71 5.655 3.955 ;
 RECT 5.515 4.095 5.655 4.965 ;
 RECT 1.265 2.52 6.245 2.66 ;
 RECT 1.91 1.98 2.05 2.52 ;
 RECT 5.995 2.46 6.245 2.52 ;
 RECT 2.585 2.34 2.835 2.52 ;
 RECT 2.43 1.63 2.57 1.99 ;
 RECT 2.43 1.475 2.775 1.63 ;
 RECT 2.515 0.825 2.655 1.475 ;
 RECT 2.32 1.99 2.57 2.13 ;
 RECT 3.915 1.625 6.17 1.765 ;
 RECT 5.93 1.545 6.17 1.625 ;
 RECT 3.915 0.975 4.23 1.115 ;
 RECT 4.09 0.805 4.23 0.975 ;
 RECT 4.07 1.765 4.21 1.92 ;
 RECT 3.915 1.115 4.055 1.625 ;
 RECT 4 1.92 4.28 2.06 ;
 RECT 6.095 3.775 6.235 3.805 ;
 RECT 6.095 3.945 6.235 4.95 ;
 RECT 6.095 3.805 6.845 3.945 ;
 END
END AODFFARX1

MACRO RDFFSRASX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.84 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.93 0.515 21.3 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.16 1.435 26.5 1.8 ;
 RECT 24.48 1.99 26.345 2.13 ;
 RECT 22.25 2.22 24.62 2.36 ;
 RECT 26.205 1.8 26.345 1.99 ;
 RECT 24.48 1.435 24.62 1.99 ;
 RECT 22.25 1.39 22.39 2.22 ;
 RECT 23.635 1.37 23.775 2.22 ;
 RECT 24.48 2.13 24.62 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.175 1.14 0.445 1.42 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.86 0.08 2.14 0.295 ;
 RECT 24.6 0.08 24.84 0.26 ;
 RECT 5.79 0.31 6.08 0.45 ;
 RECT 9.475 0.615 9.745 0.755 ;
 RECT 13.4 0.275 14.425 0.415 ;
 RECT 17.76 0.335 18.025 0.495 ;
 RECT 14.285 0.75 15.23 0.89 ;
 RECT 0 -0.08 27.84 0.08 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.275 0.08 1.415 0.97 ;
 RECT 4.685 0.08 4.92 0.46 ;
 RECT 19.405 0.08 19.545 0.82 ;
 RECT 22.25 0.08 22.39 0.36 ;
 RECT 23.465 0.08 23.605 0.35 ;
 RECT 5.87 0.08 6.01 0.31 ;
 RECT 9.54 0.08 9.68 0.615 ;
 RECT 13.4 0.415 13.54 0.945 ;
 RECT 13.4 0.08 13.54 0.275 ;
 RECT 17.815 0.08 17.955 0.335 ;
 RECT 15.09 0.89 15.23 1.11 ;
 RECT 14.285 0.415 14.425 0.75 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.155 1.475 17.465 1.7 ;
 RECT 17.155 1.7 18.47 1.765 ;
 RECT 17.325 1.765 18.47 1.84 ;
 RECT 17.325 1.84 17.465 1.885 ;
 RECT 18.33 0.915 18.47 1.7 ;
 RECT 17.325 0.915 17.465 1.475 ;
 RECT 18.33 1.84 18.47 1.885 ;
 END
 ANTENNADIFFAREA 0.7 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 17.67 2.6 17.935 2.8 ;
 RECT 19.26 2.6 19.525 2.8 ;
 RECT 4.215 2.28 4.445 2.49 ;
 RECT 9.285 2.215 9.56 2.355 ;
 RECT 0 2.8 27.84 2.96 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 2.015 2.34 2.265 2.8 ;
 RECT 1.275 1.98 1.415 2.8 ;
 RECT 5.87 1.98 6.01 2.8 ;
 RECT 6.9 2 7.04 2.8 ;
 RECT 5.39 2.07 5.53 2.8 ;
 RECT 12.31 2.335 12.58 2.8 ;
 RECT 4.26 2.49 4.4 2.8 ;
 RECT 9.35 2.355 9.49 2.8 ;
 RECT 9.35 2.195 9.49 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.15 1.475 1.585 1.76 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.905 1.155 20.285 1.405 ;
 RECT 19.905 0.56 20.045 1.155 ;
 RECT 18.845 1.905 18.985 1.915 ;
 RECT 18.845 0.51 18.985 1.765 ;
 RECT 19.905 1.905 20.045 1.91 ;
 RECT 18.845 1.765 20.045 1.905 ;
 RECT 19.905 1.405 20.045 1.765 ;
 END
 ANTENNADIFFAREA 0.568 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.745 2.115 10.075 2.47 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.23 1.795 7.49 2.04 ;
 RECT 6.69 1.795 6.92 1.83 ;
 RECT 6.69 1.655 7.49 1.795 ;
 RECT 6.69 1.62 6.92 1.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 OBS
 LAYER PO ;
 RECT 14.255 1.6 14.355 2.39 ;
 RECT 11.23 0.195 11.33 1.29 ;
 RECT 12.125 1.39 12.32 1.405 ;
 RECT 2.785 0.285 2.885 0.505 ;
 RECT 4.495 0.285 4.595 1.24 ;
 RECT 2.785 0.185 11.33 0.195 ;
 RECT 2.785 0.195 4.595 0.285 ;
 RECT 4.495 0.095 11.33 0.185 ;
 RECT 11.23 1.29 12.32 1.39 ;
 RECT 2.67 0.505 2.9 0.715 ;
 RECT 12.125 1.405 12.355 1.615 ;
 RECT 22.51 1.245 22.61 2.02 ;
 RECT 22.38 1.035 22.61 1.245 ;
 RECT 12.62 0.105 15.445 0.205 ;
 RECT 12.62 0.205 12.72 1.91 ;
 RECT 15.345 0.205 15.445 1.265 ;
 RECT 11.8 1.71 11.9 1.91 ;
 RECT 10.715 1.61 11.9 1.71 ;
 RECT 10.715 0.475 10.815 1.61 ;
 RECT 11.265 1.71 11.365 2.425 ;
 RECT 7.38 0.475 7.48 0.895 ;
 RECT 11.8 1.91 12.72 2.01 ;
 RECT 7.38 0.375 10.815 0.475 ;
 RECT 7.255 0.895 7.485 1.105 ;
 RECT 12.93 0.455 14.86 0.535 ;
 RECT 14.63 0.535 14.86 0.6 ;
 RECT 14.63 0.39 14.86 0.435 ;
 RECT 13.01 0.435 14.86 0.455 ;
 RECT 12.93 0.535 13.16 0.665 ;
 RECT 13.785 0.535 14.015 0.835 ;
 RECT 13.785 0.835 13.885 2.39 ;
 RECT 22.815 0.215 22.915 0.995 ;
 RECT 22.815 0.995 23.055 1.205 ;
 RECT 22.815 1.205 22.915 2 ;
 RECT 25.21 0.375 25.31 0.99 ;
 RECT 25.21 0.99 25.46 1.2 ;
 RECT 25.21 1.2 25.31 2.27 ;
 RECT 25.21 2.27 25.495 2.48 ;
 RECT 10.195 0.655 10.295 2.305 ;
 RECT 10.5 2.3 10.73 2.305 ;
 RECT 10.5 2.405 10.73 2.51 ;
 RECT 10.195 2.305 10.73 2.405 ;
 RECT 22.035 0.21 22.135 0.755 ;
 RECT 22.035 0.855 22.135 2.2 ;
 RECT 24.9 1.125 25 2.2 ;
 RECT 21.07 0.755 22.605 0.84 ;
 RECT 21.07 0.84 22.6 0.855 ;
 RECT 22.505 0.215 22.605 0.755 ;
 RECT 21.07 0.595 21.3 0.755 ;
 RECT 22.035 2.2 25 2.3 ;
 RECT 23.725 1.06 23.825 1.14 ;
 RECT 23.725 0.38 23.825 0.96 ;
 RECT 23.725 1.14 23.995 1.24 ;
 RECT 23.895 1.24 23.995 1.84 ;
 RECT 23.305 0.935 23.535 0.96 ;
 RECT 23.305 0.96 23.825 1.06 ;
 RECT 23.305 1.06 23.535 1.145 ;
 RECT 24.09 0.22 24.32 0.28 ;
 RECT 24.09 0.38 24.32 0.43 ;
 RECT 23.725 0.28 24.32 0.38 ;
 RECT 7.98 1.575 8.08 2.485 ;
 RECT 8.49 1.575 8.72 1.685 ;
 RECT 7.98 1.475 8.72 1.575 ;
 RECT 25.91 0.195 26.01 2.665 ;
 RECT 24.9 0.095 26.01 0.195 ;
 RECT 21.275 1.245 21.375 2.665 ;
 RECT 24.9 0.195 25 0.945 ;
 RECT 21.275 1.2 21.56 1.245 ;
 RECT 21.33 1.035 21.56 1.1 ;
 RECT 21.275 2.665 26.01 2.765 ;
 RECT 21.275 1.1 21.605 1.2 ;
 RECT 12.205 0.795 12.37 0.925 ;
 RECT 11.525 0.885 11.755 0.925 ;
 RECT 11.525 1.025 11.755 1.095 ;
 RECT 11.525 0.925 12.37 1.025 ;
 RECT 12.205 0.585 12.435 0.795 ;
 RECT 3.755 1.435 3.855 2.4 ;
 RECT 3.795 0.65 3.895 1.19 ;
 RECT 3.755 1.19 3.985 1.435 ;
 RECT 3.26 1.665 3.36 2.385 ;
 RECT 2.72 1.445 2.965 1.565 ;
 RECT 2.72 1.665 2.965 1.69 ;
 RECT 2.72 1.565 3.36 1.665 ;
 RECT 2.375 1.62 2.475 2.675 ;
 RECT 3.305 0.47 3.59 0.705 ;
 RECT 3.305 0.705 3.405 1.155 ;
 RECT 2.39 0.715 2.49 1.155 ;
 RECT 2.39 1.155 3.405 1.255 ;
 RECT 2.39 1.255 2.49 1.52 ;
 RECT 1.815 1.44 2.06 1.52 ;
 RECT 1.815 1.52 2.49 1.62 ;
 RECT 1.815 1.62 2.06 1.69 ;
 RECT 5.175 1.79 5.275 2.675 ;
 RECT 2.375 2.675 5.275 2.775 ;
 RECT 9.8 0.655 9.9 1.16 ;
 RECT 9.185 1.155 9.415 1.16 ;
 RECT 9.185 1.26 9.415 1.39 ;
 RECT 9.185 1.16 9.9 1.26 ;
 RECT 1.535 0.49 1.635 1.495 ;
 RECT 1.34 1.495 1.635 1.745 ;
 RECT 1.535 1.745 1.635 2.37 ;
 RECT 1.06 0.445 1.16 1.17 ;
 RECT 1.06 1.27 1.16 2.465 ;
 RECT 0.2 1.27 0.43 1.385 ;
 RECT 0.2 1.17 1.16 1.27 ;
 RECT 8.905 0.655 9.005 1.18 ;
 RECT 8.905 1.28 9.005 1.655 ;
 RECT 7.99 0.66 8.09 1.18 ;
 RECT 8.905 1.655 9.865 1.755 ;
 RECT 9.765 1.755 9.865 2.255 ;
 RECT 8.905 1.755 9.005 2.51 ;
 RECT 7.99 1.18 9.005 1.28 ;
 RECT 9.765 2.255 9.995 2.465 ;
 RECT 4.195 0.715 4.295 1.595 ;
 RECT 4.23 1.72 4.33 2.28 ;
 RECT 4.075 0.485 4.315 0.715 ;
 RECT 4.195 1.595 4.33 1.72 ;
 RECT 4.215 2.28 4.445 2.49 ;
 RECT 19.105 1.25 19.355 1.33 ;
 RECT 19.105 1.43 19.355 1.46 ;
 RECT 19.105 1.33 19.785 1.43 ;
 RECT 19.685 0.385 19.785 1.33 ;
 RECT 19.685 1.43 19.785 2.575 ;
 RECT 19.105 0.385 19.205 1.25 ;
 RECT 19.105 1.46 19.205 2.575 ;
 RECT 16.225 0.77 16.325 2.155 ;
 RECT 16.225 0.55 16.325 0.56 ;
 RECT 16.225 0.56 16.48 0.77 ;
 RECT 16.86 0.43 16.96 1.245 ;
 RECT 17.59 0.39 17.69 1.4 ;
 RECT 17.59 1.5 17.69 2.37 ;
 RECT 18.08 0.51 18.18 1.4 ;
 RECT 18.08 1.5 18.18 2.37 ;
 RECT 16.795 0.22 17.025 0.29 ;
 RECT 16.795 0.39 17.025 0.43 ;
 RECT 16.795 0.29 17.69 0.39 ;
 RECT 17.59 1.4 18.18 1.5 ;
 RECT 16.78 1.245 17.01 1.455 ;
 RECT 15.285 1.445 15.385 2.035 ;
 RECT 15.27 2.035 15.5 2.245 ;
 RECT 15.755 0.55 15.855 2.69 ;
 RECT 6.685 1.58 6.785 1.62 ;
 RECT 6.425 1.01 6.525 1.48 ;
 RECT 6.685 1.83 6.785 2.69 ;
 RECT 6.685 1.62 6.92 1.83 ;
 RECT 6.425 1.48 6.785 1.58 ;
 RECT 6.685 2.69 15.855 2.79 ;
 RECT 6.125 0.98 6.225 1.615 ;
 RECT 5.985 1.615 6.225 1.825 ;
 RECT 6.125 1.825 6.225 2.51 ;
 RECT 20.29 0.205 20.455 0.22 ;
 RECT 18.465 0.205 18.63 0.22 ;
 RECT 18.4 0.22 18.63 0.43 ;
 RECT 18.465 0.105 20.455 0.205 ;
 RECT 20.29 0.22 20.52 0.43 ;
 RECT 14.255 0.73 14.355 1.39 ;
 RECT 14.12 1.39 14.355 1.6 ;
 LAYER CO ;
 RECT 6.905 2.11 7.035 2.24 ;
 RECT 19.41 0.62 19.54 0.75 ;
 RECT 5.395 2.135 5.525 2.265 ;
 RECT 3.01 1.99 3.14 2.12 ;
 RECT 3.975 1.995 4.105 2.125 ;
 RECT 1.95 0.145 2.08 0.275 ;
 RECT 10.98 1.9 11.11 2.03 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 2.085 2.345 2.215 2.475 ;
 RECT 23.035 0.435 23.165 0.565 ;
 RECT 17.33 1.705 17.46 1.835 ;
 RECT 6.685 1.23 6.815 1.36 ;
 RECT 15.505 1.705 15.635 1.835 ;
 RECT 5.875 2.075 6.005 2.205 ;
 RECT 3.525 0.88 3.655 1.01 ;
 RECT 0.25 1.215 0.38 1.345 ;
 RECT 9.815 2.295 9.945 2.425 ;
 RECT 18.45 0.26 18.58 0.39 ;
 RECT 4.265 2.32 4.395 2.45 ;
 RECT 2.72 0.545 2.85 0.675 ;
 RECT 19.175 1.29 19.305 1.42 ;
 RECT 16.83 1.285 16.96 1.415 ;
 RECT 14.68 0.43 14.81 0.56 ;
 RECT 16.3 0.6 16.43 0.73 ;
 RECT 16.845 0.26 16.975 0.39 ;
 RECT 15.32 2.075 15.45 2.205 ;
 RECT 6.74 1.66 6.87 1.79 ;
 RECT 6.035 1.655 6.165 1.785 ;
 RECT 20.34 0.26 20.47 0.39 ;
 RECT 25.28 1.03 25.41 1.16 ;
 RECT 12.98 0.495 13.11 0.625 ;
 RECT 14.17 1.43 14.3 1.56 ;
 RECT 12.255 0.625 12.385 0.755 ;
 RECT 12.175 1.445 12.305 1.575 ;
 RECT 22.43 1.075 22.56 1.205 ;
 RECT 7.305 0.935 7.435 1.065 ;
 RECT 23.355 0.975 23.485 1.105 ;
 RECT 13.835 0.665 13.965 0.795 ;
 RECT 22.875 1.035 23.005 1.165 ;
 RECT 25.315 2.31 25.445 2.44 ;
 RECT 10.55 2.34 10.68 2.47 ;
 RECT 21.12 0.635 21.25 0.765 ;
 RECT 24.14 0.26 24.27 0.39 ;
 RECT 8.54 1.515 8.67 1.645 ;
 RECT 21.38 1.075 21.51 1.205 ;
 RECT 11.575 0.925 11.705 1.055 ;
 RECT 24.485 1.49 24.615 1.62 ;
 RECT 3.055 0.88 3.185 1.01 ;
 RECT 11.485 1.87 11.615 2 ;
 RECT 4.925 2.11 5.055 2.24 ;
 RECT 4.74 0.32 4.87 0.45 ;
 RECT 22.255 0.135 22.385 0.265 ;
 RECT 1.875 1.495 2.005 1.625 ;
 RECT 1.88 0.975 2.01 1.105 ;
 RECT 1.755 1.995 1.885 2.125 ;
 RECT 8.655 1.995 8.785 2.125 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 8.21 2.07 8.34 2.2 ;
 RECT 10.98 0.595 11.11 0.725 ;
 RECT 2.775 1.49 2.905 1.62 ;
 RECT 9.235 1.195 9.365 1.325 ;
 RECT 18.85 1.725 18.98 1.855 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 6.415 2.045 6.545 2.175 ;
 RECT 1.4 1.55 1.53 1.68 ;
 RECT 13.535 1.835 13.665 1.965 ;
 RECT 13.405 0.765 13.535 0.895 ;
 RECT 1.28 0.74 1.41 0.87 ;
 RECT 24.65 0.12 24.78 0.25 ;
 RECT 4.13 0.53 4.26 0.66 ;
 RECT 18.85 0.62 18.98 0.75 ;
 RECT 12.38 2.38 12.51 2.51 ;
 RECT 8.655 0.905 8.785 1.035 ;
 RECT 21.785 1.425 21.915 1.555 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 16.57 0.92 16.7 1.05 ;
 RECT 22.255 1.475 22.385 1.605 ;
 RECT 10.455 0.875 10.585 1.005 ;
 RECT 2.66 0.935 2.79 1.065 ;
 RECT 14.475 1.835 14.605 1.965 ;
 RECT 3.505 1.965 3.635 2.095 ;
 RECT 26.21 1.475 26.34 1.605 ;
 RECT 18.335 1.705 18.465 1.835 ;
 RECT 19.91 1.71 20.04 1.84 ;
 RECT 17.33 0.975 17.46 1.105 ;
 RECT 0.81 0.74 0.94 0.87 ;
 RECT 2.595 1.825 2.725 1.955 ;
 RECT 10.455 1.945 10.585 2.075 ;
 RECT 1.28 2.05 1.41 2.18 ;
 RECT 21.535 0.505 21.665 0.635 ;
 RECT 7.73 2.015 7.86 2.145 ;
 RECT 23.47 0.12 23.6 0.25 ;
 RECT 23.035 1.485 23.165 1.615 ;
 RECT 25.43 1.465 25.56 1.595 ;
 RECT 15.975 1.705 16.105 1.835 ;
 RECT 25.43 0.595 25.56 0.725 ;
 RECT 3.805 1.235 3.935 1.365 ;
 RECT 9.355 2.225 9.485 2.355 ;
 RECT 18.335 0.975 18.465 1.105 ;
 RECT 19.325 2.64 19.455 2.77 ;
 RECT 0.81 2.115 0.94 2.245 ;
 RECT 17.82 0.36 17.95 0.49 ;
 RECT 19.91 0.63 20.04 0.76 ;
 RECT 23.975 0.595 24.105 0.725 ;
 RECT 3.41 0.525 3.54 0.655 ;
 RECT 4.525 1.675 4.655 1.805 ;
 RECT 16.45 1.705 16.58 1.835 ;
 RECT 17.735 2.64 17.865 2.77 ;
 RECT 24.115 1.405 24.245 1.535 ;
 RECT 7.735 0.905 7.865 1.035 ;
 RECT 5.875 0.315 6.005 0.445 ;
 RECT 8.21 0.905 8.34 1.035 ;
 RECT 11.485 0.595 11.615 0.725 ;
 RECT 9.545 0.62 9.675 0.75 ;
 RECT 23.64 1.445 23.77 1.575 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 14.51 1.035 14.64 1.165 ;
 RECT 15.095 0.91 15.225 1.04 ;
 LAYER M1 ;
 RECT 7.66 0.9 7.935 1.04 ;
 RECT 1.795 1.63 1.935 1.99 ;
 RECT 1.795 1.475 2.1 1.63 ;
 RECT 1.875 0.905 2.015 1.475 ;
 RECT 1.685 1.99 1.935 2.13 ;
 RECT 3.465 1.06 3.605 1.67 ;
 RECT 3.465 1.81 3.605 1.96 ;
 RECT 3.465 1.79 4.925 1.81 ;
 RECT 3.465 0.805 3.66 1.06 ;
 RECT 3.43 1.96 3.71 2.1 ;
 RECT 3.465 1.67 6.22 1.79 ;
 RECT 4.75 1.65 6.22 1.67 ;
 RECT 5.985 1.615 6.215 1.65 ;
 RECT 5.985 1.79 6.215 1.825 ;
 RECT 23.97 0.73 24.11 1.04 ;
 RECT 24.11 1.18 24.25 1.605 ;
 RECT 23.905 0.59 24.18 0.73 ;
 RECT 25.23 0.99 25.46 1.04 ;
 RECT 23.97 1.04 25.46 1.18 ;
 RECT 25.23 1.18 25.46 1.2 ;
 RECT 24.09 0.29 24.46 0.43 ;
 RECT 24.32 0.43 24.46 0.71 ;
 RECT 24.09 0.22 24.32 0.29 ;
 RECT 25.74 0.85 25.88 1.385 ;
 RECT 25.425 1.525 25.565 1.73 ;
 RECT 24.32 0.71 25.88 0.85 ;
 RECT 25.425 0.51 25.565 0.71 ;
 RECT 25.425 1.385 25.88 1.525 ;
 RECT 21.33 1.225 21.56 1.245 ;
 RECT 21.33 1.195 21.92 1.225 ;
 RECT 21.47 1.015 21.78 1.035 ;
 RECT 21.33 1.035 21.78 1.055 ;
 RECT 21.605 0.64 21.745 1.015 ;
 RECT 21.78 1.225 21.92 1.75 ;
 RECT 21.485 0.5 21.745 0.64 ;
 RECT 22.38 1.035 22.61 1.055 ;
 RECT 22.38 1.195 22.61 1.245 ;
 RECT 21.33 1.055 22.61 1.195 ;
 RECT 23.35 1.145 23.49 1.345 ;
 RECT 23.03 1.485 23.17 1.76 ;
 RECT 23.35 0.73 23.49 0.935 ;
 RECT 23.03 0.355 23.17 0.59 ;
 RECT 23.03 1.345 23.49 1.485 ;
 RECT 23.305 0.935 23.535 1.145 ;
 RECT 23.03 0.59 23.49 0.73 ;
 RECT 20.29 0.36 20.52 0.43 ;
 RECT 21.885 0.36 22.025 0.565 ;
 RECT 20.29 0.22 22.025 0.36 ;
 RECT 22.625 0.705 22.765 0.75 ;
 RECT 22.75 0.995 23.055 1.205 ;
 RECT 22.75 0.89 22.89 0.995 ;
 RECT 22.625 0.75 22.89 0.89 ;
 RECT 21.885 0.565 22.765 0.705 ;
 RECT 15.525 0.775 15.665 1.405 ;
 RECT 16.25 0.56 16.48 0.635 ;
 RECT 14.505 1.405 15.665 1.545 ;
 RECT 14.505 1.545 14.645 1.83 ;
 RECT 14.505 1.17 14.645 1.405 ;
 RECT 13.46 1.83 14.71 1.97 ;
 RECT 14.435 1.03 14.715 1.17 ;
 RECT 18.445 0.43 18.585 0.635 ;
 RECT 18.4 0.36 18.63 0.43 ;
 RECT 15.525 0.635 18.585 0.775 ;
 RECT 19.125 0.36 19.265 1.25 ;
 RECT 18.4 0.22 19.265 0.36 ;
 RECT 19.125 1.25 19.355 1.46 ;
 RECT 14.63 0.28 17.025 0.42 ;
 RECT 14.63 0.42 14.86 0.6 ;
 RECT 16.795 0.22 17.025 0.28 ;
 RECT 16.795 0.42 17.025 0.43 ;
 RECT 11.48 0.525 11.62 0.885 ;
 RECT 11.48 1.095 11.62 2.065 ;
 RECT 11.48 0.885 11.755 1.095 ;
 RECT 9.355 1.66 9.495 1.915 ;
 RECT 9 1.915 9.495 2.055 ;
 RECT 8.205 1.04 8.345 2.34 ;
 RECT 8.205 0.895 8.345 0.9 ;
 RECT 9 2.055 9.14 2.34 ;
 RECT 8.135 0.9 8.41 1.04 ;
 RECT 8.205 2.34 9.14 2.48 ;
 RECT 9.355 1.52 11.115 1.66 ;
 RECT 10.975 0.525 11.115 1.52 ;
 RECT 10.975 1.66 11.115 2.11 ;
 RECT 10.45 0.765 10.59 1.52 ;
 RECT 10.45 1.66 10.59 2.145 ;
 RECT 13.785 0.57 14.015 0.95 ;
 RECT 12.205 0.585 13.16 0.63 ;
 RECT 12.93 0.63 13.16 0.665 ;
 RECT 12.93 0.455 13.16 0.49 ;
 RECT 12.23 0.49 13.16 0.585 ;
 RECT 12.205 0.63 12.435 0.795 ;
 RECT 3.8 0.895 7.485 1.035 ;
 RECT 7.255 1.035 7.485 1.105 ;
 RECT 3.8 0.66 3.94 0.895 ;
 RECT 3.34 0.52 3.94 0.66 ;
 RECT 13.775 1.23 13.915 1.42 ;
 RECT 11.925 1.09 13.915 1.23 ;
 RECT 11.925 0.385 12.065 1.09 ;
 RECT 9.915 0.385 10.055 0.895 ;
 RECT 9.91 0.255 12.065 0.385 ;
 RECT 9.91 0.245 12.06 0.255 ;
 RECT 9.915 0.22 10.055 0.245 ;
 RECT 9 0.895 10.055 1.035 ;
 RECT 9 0.745 9.14 0.895 ;
 RECT 4.08 0.605 9.14 0.745 ;
 RECT 4.08 0.485 4.395 0.605 ;
 RECT 14.12 1.39 14.35 1.42 ;
 RECT 13.775 1.42 14.35 1.56 ;
 RECT 14.12 1.56 14.35 1.6 ;
 RECT 2.655 1.67 2.795 1.82 ;
 RECT 2.655 1.96 2.795 2.25 ;
 RECT 2.655 0.715 2.795 1.44 ;
 RECT 2.655 1.44 2.91 1.67 ;
 RECT 2.655 0.505 2.9 0.715 ;
 RECT 2.525 1.82 2.795 1.96 ;
 RECT 0.585 0.875 0.725 1.195 ;
 RECT 0.585 1.335 0.725 2.11 ;
 RECT 0.585 2.25 0.725 2.255 ;
 RECT 0.585 2.11 1.01 2.25 ;
 RECT 0.585 0.735 1.01 0.875 ;
 RECT 1.555 0.6 1.695 1.195 ;
 RECT 0.585 1.195 1.695 1.335 ;
 RECT 3.05 0.36 3.19 1.915 ;
 RECT 2.285 0.36 2.425 0.46 ;
 RECT 3.005 1.915 3.19 2.17 ;
 RECT 2.285 0.22 3.19 0.36 ;
 RECT 1.555 0.46 2.425 0.6 ;
 RECT 16.335 1.7 16.63 1.84 ;
 RECT 16.335 1.84 16.475 2.075 ;
 RECT 15.64 1.84 15.78 2.075 ;
 RECT 15.445 1.7 15.78 1.84 ;
 RECT 15.64 2.075 16.475 2.215 ;
 RECT 16.53 1.055 16.67 1.245 ;
 RECT 15.97 1.385 16.11 1.625 ;
 RECT 16.78 1.385 17.01 1.455 ;
 RECT 15.97 1.245 17.01 1.385 ;
 RECT 16.5 0.915 16.8 1.055 ;
 RECT 15.94 1.625 16.195 1.92 ;
 RECT 17.04 2.205 17.18 2.39 ;
 RECT 12.895 2.39 17.18 2.53 ;
 RECT 12.895 1.895 13.035 2.39 ;
 RECT 11.77 1.755 13.035 1.895 ;
 RECT 11.77 1.895 11.91 2.34 ;
 RECT 10.5 2.3 10.73 2.34 ;
 RECT 10.5 2.48 10.73 2.51 ;
 RECT 10.5 2.34 11.91 2.48 ;
 RECT 17.04 2.065 21.065 2.205 ;
 RECT 20.925 2.205 21.065 2.52 ;
 RECT 25.265 2.48 25.405 2.52 ;
 RECT 20.925 2.52 25.405 2.66 ;
 RECT 25.265 2.27 25.495 2.48 ;
 RECT 13.175 1.56 13.315 2.11 ;
 RECT 13.175 2.11 15.5 2.245 ;
 RECT 13.175 2.245 15.495 2.25 ;
 RECT 15.27 2.035 15.5 2.11 ;
 RECT 12.125 1.405 12.355 1.42 ;
 RECT 12.125 1.56 12.355 1.615 ;
 RECT 12.125 1.42 13.315 1.56 ;
 RECT 8.65 1.685 9.195 1.775 ;
 RECT 9.055 1.33 9.195 1.635 ;
 RECT 8.49 1.635 9.195 1.685 ;
 RECT 8.65 1.04 8.79 1.475 ;
 RECT 8.49 1.475 8.79 1.635 ;
 RECT 8.65 1.775 8.79 2.18 ;
 RECT 9.055 1.19 9.415 1.33 ;
 RECT 8.58 0.9 8.855 1.04 ;
 RECT 3.905 2.105 5.125 2.13 ;
 RECT 3.905 1.99 4.935 2.105 ;
 RECT 4.77 2.13 5.125 2.245 ;
 RECT 3.75 1.225 7.115 1.25 ;
 RECT 6.41 1.365 6.55 2.25 ;
 RECT 3.75 1.215 3.98 1.225 ;
 RECT 3.75 1.365 3.98 1.39 ;
 RECT 7.725 1.04 7.865 1.25 ;
 RECT 7.725 1.39 7.865 2.215 ;
 RECT 7.725 0.885 7.865 0.9 ;
 RECT 3.75 1.25 7.865 1.365 ;
 RECT 6.975 1.365 7.865 1.39 ;
 END
END RDFFSRASX1

MACRO RDFFSRASX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 29.76 BY 2.88 ;
 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.155 1.475 1.57 1.76 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.72 2.115 10.1 2.48 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 22.905 0.515 23.29 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.86 0.08 2.14 0.295 ;
 RECT 26.59 0.08 26.83 0.26 ;
 RECT 5.79 0.31 6.08 0.45 ;
 RECT 9.475 0.615 9.745 0.755 ;
 RECT 13.4 0.275 14.425 0.415 ;
 RECT 17.98 0.335 18.245 0.495 ;
 RECT 18.985 0.335 19.25 0.495 ;
 RECT 14.285 0.75 15.23 0.89 ;
 RECT 0 -0.08 29.76 0.08 ;
 RECT 1.275 0.08 1.415 0.97 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 4.685 0.08 4.92 0.46 ;
 RECT 20.5 0.08 20.64 0.82 ;
 RECT 21.565 0.08 21.705 0.82 ;
 RECT 24.24 0.08 24.38 0.36 ;
 RECT 25.455 0.08 25.595 0.35 ;
 RECT 5.87 0.08 6.01 0.31 ;
 RECT 9.54 0.08 9.68 0.615 ;
 RECT 13.4 0.415 13.54 0.945 ;
 RECT 13.4 0.08 13.54 0.275 ;
 RECT 18.035 0.08 18.175 0.335 ;
 RECT 19.04 0.08 19.18 0.335 ;
 RECT 15.09 0.89 15.23 1.11 ;
 RECT 14.285 0.415 14.425 0.75 ;
 END
 END VSS

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.23 1.795 7.485 2.045 ;
 RECT 6.69 1.655 7.485 1.795 ;
 RECT 6.69 1.795 6.92 1.83 ;
 RECT 6.69 1.62 6.92 1.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 28.11 1.435 28.47 1.8 ;
 RECT 26.47 1.99 28.335 2.13 ;
 RECT 24.24 2.22 26.61 2.36 ;
 RECT 26.47 1.435 26.61 1.99 ;
 RECT 28.195 1.8 28.335 1.99 ;
 RECT 24.24 1.39 24.38 2.22 ;
 RECT 25.625 1.37 25.765 2.22 ;
 RECT 26.47 2.13 26.61 2.22 ;
 END
 END VDDG

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 4.175 2.27 4.405 2.48 ;
 RECT 9.285 2.215 9.56 2.355 ;
 RECT 0 2.8 29.76 2.96 ;
 RECT 2.015 2.34 2.265 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.275 1.98 1.415 2.8 ;
 RECT 6.9 2 7.04 2.8 ;
 RECT 5.87 1.98 6.01 2.8 ;
 RECT 5.39 2.07 5.53 2.8 ;
 RECT 9.35 2.195 9.49 2.215 ;
 RECT 12.31 2.335 12.58 2.8 ;
 RECT 20.415 2.57 20.555 2.8 ;
 RECT 17.95 2.57 18.09 2.8 ;
 RECT 18.955 2.57 19.095 2.8 ;
 RECT 21.48 2.57 21.62 2.8 ;
 RECT 4.22 2.48 4.36 2.8 ;
 RECT 9.35 2.355 9.49 2.8 ;
 END
 END VDD

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.18 1.145 0.445 1.41 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.43 1.16 17.735 1.445 ;
 RECT 17.545 0.915 17.685 1.16 ;
 RECT 17.545 1.84 17.685 1.885 ;
 RECT 17.545 1.445 17.685 1.7 ;
 RECT 18.55 1.84 18.69 1.885 ;
 RECT 18.55 0.915 18.69 1.7 ;
 RECT 19.525 1.84 19.665 1.885 ;
 RECT 19.525 0.915 19.665 1.7 ;
 RECT 17.545 1.7 19.665 1.84 ;
 END
 ANTENNADIFFAREA 1.145 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 21 0.82 21.29 1.08 ;
 RECT 21 0.56 21.14 0.82 ;
 RECT 21 1.905 21.14 1.91 ;
 RECT 21 1.08 21.14 1.765 ;
 RECT 22.065 1.905 22.205 1.91 ;
 RECT 22.065 0.56 22.205 1.765 ;
 RECT 19.94 1.905 20.08 1.915 ;
 RECT 19.94 0.51 20.08 1.765 ;
 RECT 19.94 1.765 22.205 1.905 ;
 END
 ANTENNADIFFAREA 0.937 ;
 END Q

 OBS
 LAYER PO ;
 RECT 25.715 0.28 26.31 0.38 ;
 RECT 24.025 0.855 24.125 2.2 ;
 RECT 26.89 1.125 26.99 2.2 ;
 RECT 23.06 0.755 24.595 0.84 ;
 RECT 23.06 0.84 24.59 0.855 ;
 RECT 24.495 0.215 24.595 0.755 ;
 RECT 24.025 0.21 24.125 0.755 ;
 RECT 23.06 0.595 23.29 0.755 ;
 RECT 24.025 2.2 26.99 2.3 ;
 RECT 10.195 0.655 10.295 2.305 ;
 RECT 10.5 2.3 10.73 2.305 ;
 RECT 10.5 2.405 10.73 2.51 ;
 RECT 10.195 2.305 10.73 2.405 ;
 RECT 20.185 1.33 21.945 1.43 ;
 RECT 21.265 1.43 21.365 2.455 ;
 RECT 21.845 0.195 21.945 1.33 ;
 RECT 20.185 1.2 20.395 1.33 ;
 RECT 20.185 1.43 20.395 1.435 ;
 RECT 20.2 0.385 20.3 1.2 ;
 RECT 20.2 1.435 20.3 2.455 ;
 RECT 20.78 0.385 20.88 1.33 ;
 RECT 20.78 1.43 20.88 2.46 ;
 RECT 21.265 0.385 21.365 1.33 ;
 RECT 21.845 1.43 21.945 2.465 ;
 RECT 22.475 0.195 22.705 0.43 ;
 RECT 21.845 0.095 22.705 0.195 ;
 RECT 14.255 0.73 14.355 1.39 ;
 RECT 14.12 1.39 14.355 1.6 ;
 RECT 14.255 1.6 14.355 2.39 ;
 RECT 12.93 0.455 14.86 0.535 ;
 RECT 14.63 0.535 14.86 0.6 ;
 RECT 13.785 0.535 14.015 0.835 ;
 RECT 13.785 0.835 13.885 2.39 ;
 RECT 14.63 0.39 14.86 0.435 ;
 RECT 13.01 0.435 14.86 0.455 ;
 RECT 12.93 0.535 13.16 0.665 ;
 RECT 15.285 1.445 15.385 2.035 ;
 RECT 15.27 2.035 15.5 2.245 ;
 RECT 17.81 0.39 17.91 1.4 ;
 RECT 17.81 1.5 17.91 2.37 ;
 RECT 16.86 0.43 16.96 1.245 ;
 RECT 19.305 0.51 19.405 1.4 ;
 RECT 19.305 1.5 19.405 2.37 ;
 RECT 18.815 0.515 18.915 1.4 ;
 RECT 18.815 1.5 18.915 2.37 ;
 RECT 17.81 1.4 19.405 1.5 ;
 RECT 18.3 0.51 18.4 1.4 ;
 RECT 18.3 1.5 18.4 2.37 ;
 RECT 16.795 0.22 17.025 0.29 ;
 RECT 16.795 0.39 17.025 0.43 ;
 RECT 16.795 0.29 17.91 0.39 ;
 RECT 16.81 1.245 17.04 1.455 ;
 RECT 16.225 0.77 16.325 2.155 ;
 RECT 16.225 0.55 16.325 0.56 ;
 RECT 16.225 0.56 16.48 0.77 ;
 RECT 27.2 0.375 27.3 0.99 ;
 RECT 27.2 0.99 27.45 1.2 ;
 RECT 27.2 1.2 27.3 2.27 ;
 RECT 27.2 2.27 27.485 2.48 ;
 RECT 24.805 0.215 24.905 0.995 ;
 RECT 24.805 0.995 25.045 1.205 ;
 RECT 24.805 1.205 24.905 2 ;
 RECT 15.755 0.55 15.855 2.69 ;
 RECT 6.685 1.58 6.785 1.62 ;
 RECT 6.425 1.01 6.525 1.48 ;
 RECT 6.685 1.83 6.785 2.69 ;
 RECT 6.685 1.62 6.92 1.83 ;
 RECT 6.425 1.48 6.785 1.58 ;
 RECT 6.685 2.69 15.855 2.79 ;
 RECT 11.23 0.195 11.33 1.29 ;
 RECT 12.125 1.39 12.32 1.405 ;
 RECT 2.785 0.285 2.885 0.505 ;
 RECT 4.495 0.285 4.595 1.24 ;
 RECT 2.785 0.185 11.33 0.195 ;
 RECT 2.785 0.195 4.595 0.285 ;
 RECT 4.495 0.095 11.33 0.185 ;
 RECT 11.23 1.29 12.32 1.39 ;
 RECT 2.67 0.505 2.9 0.715 ;
 RECT 12.125 1.405 12.355 1.615 ;
 RECT 3.755 1.5 3.855 2.4 ;
 RECT 3.755 1.435 3.895 1.5 ;
 RECT 3.795 0.65 3.895 1.2 ;
 RECT 3.755 1.2 3.985 1.435 ;
 RECT 2.375 1.62 2.475 2.675 ;
 RECT 3.305 0.47 3.59 0.705 ;
 RECT 3.305 0.705 3.405 1.155 ;
 RECT 2.39 0.715 2.49 1.155 ;
 RECT 2.39 1.155 3.405 1.255 ;
 RECT 2.39 1.255 2.49 1.52 ;
 RECT 2.375 2.675 5.275 2.775 ;
 RECT 5.175 1.79 5.275 2.675 ;
 RECT 1.815 1.44 2.06 1.52 ;
 RECT 1.815 1.52 2.49 1.62 ;
 RECT 1.815 1.62 2.06 1.69 ;
 RECT 9.8 0.655 9.9 1.16 ;
 RECT 9.185 1.26 9.415 1.395 ;
 RECT 9.185 1.16 9.9 1.26 ;
 RECT 1.535 0.49 1.635 1.495 ;
 RECT 1.34 1.495 1.635 1.745 ;
 RECT 1.535 1.745 1.635 2.37 ;
 RECT 3.26 1.665 3.36 2.345 ;
 RECT 2.72 1.445 2.965 1.565 ;
 RECT 2.72 1.565 3.36 1.665 ;
 RECT 2.72 1.665 2.965 1.69 ;
 RECT 1.06 0.405 1.16 1.175 ;
 RECT 1.06 1.275 1.16 2.465 ;
 RECT 0.205 1.275 0.435 1.39 ;
 RECT 0.205 1.175 1.16 1.275 ;
 RECT 8.905 0.655 9.005 1.18 ;
 RECT 8.905 1.28 9.005 1.655 ;
 RECT 7.99 0.66 8.09 1.18 ;
 RECT 8.905 1.655 9.865 1.755 ;
 RECT 9.765 1.755 9.865 2.265 ;
 RECT 8.905 1.755 9.005 2.51 ;
 RECT 7.99 1.18 9.005 1.28 ;
 RECT 9.765 2.265 9.995 2.475 ;
 RECT 4.195 0.715 4.295 1.61 ;
 RECT 4.23 1.71 4.33 2.27 ;
 RECT 4.075 0.485 4.315 0.715 ;
 RECT 4.195 1.61 4.33 1.71 ;
 RECT 4.175 2.27 4.405 2.48 ;
 RECT 27.9 0.195 28 2.665 ;
 RECT 26.89 0.095 28 0.195 ;
 RECT 23.265 1.245 23.365 2.665 ;
 RECT 26.89 0.195 26.99 0.945 ;
 RECT 23.265 1.2 23.55 1.245 ;
 RECT 23.32 1.035 23.55 1.1 ;
 RECT 23.265 2.665 28 2.765 ;
 RECT 23.265 1.1 23.595 1.2 ;
 RECT 6.125 0.98 6.225 1.615 ;
 RECT 5.985 1.615 6.225 1.825 ;
 RECT 6.125 1.825 6.225 2.51 ;
 RECT 12.62 0.105 15.445 0.205 ;
 RECT 12.62 0.205 12.72 1.91 ;
 RECT 15.345 0.205 15.445 1.265 ;
 RECT 11.8 1.71 11.9 1.91 ;
 RECT 10.715 1.61 11.9 1.71 ;
 RECT 10.715 0.475 10.815 1.61 ;
 RECT 11.265 1.71 11.365 2.425 ;
 RECT 7.38 0.475 7.48 0.895 ;
 RECT 11.8 1.91 12.72 2.01 ;
 RECT 7.38 0.375 10.815 0.475 ;
 RECT 7.255 0.895 7.485 1.105 ;
 RECT 7.98 1.575 8.08 2.485 ;
 RECT 8.49 1.575 8.72 1.685 ;
 RECT 7.98 1.475 8.72 1.575 ;
 RECT 24.5 1.245 24.6 2.02 ;
 RECT 24.37 1.035 24.6 1.245 ;
 RECT 11.525 0.885 11.755 0.925 ;
 RECT 11.525 0.925 12.37 1.025 ;
 RECT 11.525 1.025 11.755 1.095 ;
 RECT 12.205 0.795 12.37 0.925 ;
 RECT 12.205 0.585 12.435 0.795 ;
 RECT 25.715 0.38 25.815 0.96 ;
 RECT 25.715 1.06 25.815 1.14 ;
 RECT 25.295 0.935 25.525 0.96 ;
 RECT 25.295 0.96 25.815 1.06 ;
 RECT 25.295 1.06 25.525 1.145 ;
 RECT 25.715 1.14 25.985 1.24 ;
 RECT 25.885 1.24 25.985 1.84 ;
 RECT 26.08 0.22 26.31 0.28 ;
 RECT 26.08 0.38 26.31 0.43 ;
 LAYER CO ;
 RECT 26.64 0.12 26.77 0.25 ;
 RECT 3.41 0.525 3.54 0.655 ;
 RECT 17.55 1.705 17.68 1.835 ;
 RECT 8.655 1.995 8.785 2.125 ;
 RECT 20.225 1.25 20.355 1.38 ;
 RECT 5.875 2.075 6.005 2.205 ;
 RECT 10.98 0.595 11.11 0.725 ;
 RECT 2.595 1.825 2.725 1.955 ;
 RECT 21.485 2.64 21.615 2.77 ;
 RECT 19.945 1.725 20.075 1.855 ;
 RECT 13.405 0.765 13.535 0.895 ;
 RECT 18.04 0.36 18.17 0.49 ;
 RECT 19.945 0.62 20.075 0.75 ;
 RECT 19.53 0.975 19.66 1.105 ;
 RECT 24.245 1.475 24.375 1.605 ;
 RECT 0.255 1.22 0.385 1.35 ;
 RECT 9.815 2.305 9.945 2.435 ;
 RECT 4.225 2.31 4.355 2.44 ;
 RECT 25.345 0.975 25.475 1.105 ;
 RECT 13.835 0.665 13.965 0.795 ;
 RECT 16.86 1.285 16.99 1.415 ;
 RECT 14.68 0.43 14.81 0.56 ;
 RECT 23.37 1.075 23.5 1.205 ;
 RECT 6.035 1.655 6.165 1.785 ;
 RECT 7.305 0.935 7.435 1.065 ;
 RECT 11.575 0.925 11.705 1.055 ;
 RECT 2.72 0.545 2.85 0.675 ;
 RECT 8.54 1.515 8.67 1.645 ;
 RECT 24.42 1.075 24.55 1.205 ;
 RECT 12.255 0.625 12.385 0.755 ;
 RECT 26.13 0.26 26.26 0.39 ;
 RECT 23.11 0.635 23.24 0.765 ;
 RECT 10.55 2.34 10.68 2.47 ;
 RECT 22.525 0.26 22.655 0.39 ;
 RECT 14.17 1.43 14.3 1.56 ;
 RECT 27.27 1.03 27.4 1.16 ;
 RECT 12.98 0.495 13.11 0.625 ;
 RECT 15.32 2.075 15.45 2.205 ;
 RECT 16.845 0.26 16.975 0.39 ;
 RECT 16.3 0.6 16.43 0.73 ;
 RECT 27.305 2.31 27.435 2.44 ;
 RECT 24.865 1.035 24.995 1.165 ;
 RECT 6.74 1.66 6.87 1.79 ;
 RECT 12.175 1.445 12.305 1.575 ;
 RECT 5.395 2.135 5.525 2.265 ;
 RECT 1.28 2.05 1.41 2.18 ;
 RECT 1.755 1.995 1.885 2.125 ;
 RECT 14.475 1.835 14.605 1.965 ;
 RECT 9.545 0.62 9.675 0.75 ;
 RECT 13.535 1.835 13.665 1.965 ;
 RECT 16.45 1.705 16.58 1.835 ;
 RECT 11.485 0.595 11.615 0.725 ;
 RECT 18.96 2.64 19.09 2.77 ;
 RECT 3.805 1.25 3.935 1.38 ;
 RECT 11.485 1.87 11.615 2 ;
 RECT 5.875 0.315 6.005 0.445 ;
 RECT 25.965 0.595 26.095 0.725 ;
 RECT 4.925 2.11 5.055 2.24 ;
 RECT 6.415 2.045 6.545 2.175 ;
 RECT 0.81 2.115 0.94 2.245 ;
 RECT 7.73 2.015 7.86 2.145 ;
 RECT 25.025 0.435 25.155 0.565 ;
 RECT 1.28 0.74 1.41 0.87 ;
 RECT 9.355 2.225 9.485 2.355 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 25.025 1.485 25.155 1.615 ;
 RECT 26.475 1.49 26.605 1.62 ;
 RECT 22.07 0.63 22.2 0.76 ;
 RECT 3.525 0.88 3.655 1.01 ;
 RECT 15.975 1.705 16.105 1.835 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 9.235 1.2 9.365 1.33 ;
 RECT 1.88 0.975 2.01 1.105 ;
 RECT 25.46 0.12 25.59 0.25 ;
 RECT 4.13 0.53 4.26 0.66 ;
 RECT 23.525 0.505 23.655 0.635 ;
 RECT 18.555 1.705 18.685 1.835 ;
 RECT 8.21 0.905 8.34 1.035 ;
 RECT 17.955 2.64 18.085 2.77 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 3.055 0.88 3.185 1.01 ;
 RECT 3.01 1.965 3.14 2.095 ;
 RECT 2.775 1.49 2.905 1.62 ;
 RECT 1.875 1.495 2.005 1.625 ;
 RECT 3.975 1.965 4.105 2.095 ;
 RECT 12.38 2.38 12.51 2.51 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 15.505 1.705 15.635 1.835 ;
 RECT 24.245 0.135 24.375 0.265 ;
 RECT 10.98 1.9 11.11 2.03 ;
 RECT 27.42 0.595 27.55 0.725 ;
 RECT 25.63 1.445 25.76 1.575 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 26.105 1.405 26.235 1.535 ;
 RECT 4.455 1.68 4.585 1.81 ;
 RECT 6.905 2.11 7.035 2.24 ;
 RECT 21.005 0.63 21.135 0.76 ;
 RECT 7.735 0.905 7.865 1.035 ;
 RECT 8.21 2.07 8.34 2.2 ;
 RECT 27.42 1.465 27.55 1.595 ;
 RECT 21.005 1.71 21.135 1.84 ;
 RECT 14.51 1.035 14.64 1.165 ;
 RECT 1.4 1.55 1.53 1.68 ;
 RECT 2.66 0.935 2.79 1.065 ;
 RECT 17.55 0.975 17.68 1.105 ;
 RECT 16.57 0.92 16.7 1.05 ;
 RECT 15.095 0.91 15.225 1.04 ;
 RECT 22.07 1.71 22.2 1.84 ;
 RECT 19.53 1.705 19.66 1.835 ;
 RECT 23.775 1.425 23.905 1.555 ;
 RECT 20.505 0.62 20.635 0.75 ;
 RECT 4.74 0.32 4.87 0.45 ;
 RECT 3.505 1.935 3.635 2.065 ;
 RECT 18.555 0.975 18.685 1.105 ;
 RECT 2.085 2.345 2.215 2.475 ;
 RECT 10.455 1.945 10.585 2.075 ;
 RECT 28.2 1.475 28.33 1.605 ;
 RECT 0.81 0.74 0.94 0.87 ;
 RECT 20.42 2.64 20.55 2.77 ;
 RECT 6.685 1.23 6.815 1.36 ;
 RECT 1.95 0.145 2.08 0.275 ;
 RECT 21.57 0.62 21.7 0.75 ;
 RECT 19.045 0.36 19.175 0.49 ;
 RECT 8.655 0.905 8.785 1.035 ;
 RECT 10.455 0.875 10.585 1.005 ;
 LAYER M1 ;
 RECT 1.795 1.475 2.1 1.63 ;
 RECT 1.875 0.905 2.015 1.475 ;
 RECT 1.685 1.99 1.935 2.13 ;
 RECT 25.96 0.73 26.1 1.04 ;
 RECT 26.1 1.18 26.24 1.605 ;
 RECT 25.895 0.59 26.17 0.73 ;
 RECT 27.22 0.99 27.45 1.04 ;
 RECT 25.96 1.04 27.45 1.18 ;
 RECT 27.22 1.18 27.45 1.2 ;
 RECT 26.08 0.29 26.45 0.43 ;
 RECT 26.31 0.43 26.45 0.71 ;
 RECT 26.08 0.22 26.31 0.29 ;
 RECT 27.73 0.85 27.87 1.385 ;
 RECT 27.415 1.525 27.555 1.73 ;
 RECT 26.31 0.71 27.87 0.85 ;
 RECT 27.415 0.51 27.555 0.71 ;
 RECT 27.415 1.385 27.87 1.525 ;
 RECT 25.34 1.145 25.48 1.345 ;
 RECT 25.02 1.485 25.16 1.76 ;
 RECT 25.34 0.73 25.48 0.935 ;
 RECT 25.02 0.355 25.16 0.59 ;
 RECT 25.02 1.345 25.48 1.485 ;
 RECT 25.295 0.935 25.525 1.145 ;
 RECT 25.02 0.59 25.48 0.73 ;
 RECT 23.32 1.225 23.55 1.245 ;
 RECT 23.32 1.195 23.91 1.225 ;
 RECT 23.46 1.015 23.77 1.035 ;
 RECT 23.32 1.035 23.77 1.055 ;
 RECT 23.595 0.64 23.735 1.015 ;
 RECT 23.77 1.225 23.91 1.75 ;
 RECT 23.475 0.5 23.735 0.64 ;
 RECT 24.37 1.035 24.6 1.055 ;
 RECT 24.37 1.195 24.6 1.245 ;
 RECT 23.32 1.055 24.6 1.195 ;
 RECT 22.475 0.36 22.705 0.43 ;
 RECT 22.475 0.22 24.015 0.36 ;
 RECT 23.875 0.36 24.015 0.565 ;
 RECT 24.615 0.705 24.755 0.75 ;
 RECT 24.74 0.995 25.045 1.205 ;
 RECT 24.74 0.89 24.88 0.995 ;
 RECT 24.615 0.75 24.88 0.89 ;
 RECT 23.875 0.565 24.755 0.705 ;
 RECT 15.525 0.775 15.665 1.405 ;
 RECT 16.25 0.56 16.48 0.635 ;
 RECT 14.505 1.405 15.665 1.545 ;
 RECT 14.505 1.545 14.645 1.83 ;
 RECT 14.505 1.17 14.645 1.405 ;
 RECT 13.46 1.83 14.71 1.97 ;
 RECT 14.435 1.03 14.715 1.17 ;
 RECT 19.54 0.36 19.68 0.635 ;
 RECT 15.525 0.635 19.68 0.775 ;
 RECT 20.22 0.36 20.36 1.46 ;
 RECT 19.54 0.22 20.36 0.36 ;
 RECT 12.205 0.585 13.16 0.63 ;
 RECT 12.205 0.63 12.435 0.795 ;
 RECT 12.23 0.49 13.16 0.585 ;
 RECT 12.93 0.455 13.16 0.49 ;
 RECT 12.93 0.63 13.16 0.665 ;
 RECT 13.785 0.57 14.015 0.95 ;
 RECT 16.795 0.22 17.025 0.28 ;
 RECT 16.795 0.42 17.025 0.43 ;
 RECT 14.63 0.28 17.025 0.42 ;
 RECT 14.63 0.42 14.86 0.6 ;
 RECT 11.48 0.525 11.62 0.885 ;
 RECT 11.48 1.095 11.62 2.065 ;
 RECT 11.48 0.885 11.755 1.095 ;
 RECT 9.365 1.66 9.505 1.915 ;
 RECT 9 1.915 9.505 2.055 ;
 RECT 8.205 1.04 8.345 2.34 ;
 RECT 8.205 0.895 8.345 0.9 ;
 RECT 9 2.055 9.14 2.34 ;
 RECT 8.135 0.9 8.41 1.04 ;
 RECT 8.205 2.34 9.14 2.48 ;
 RECT 9.365 1.52 11.115 1.66 ;
 RECT 10.45 0.765 10.59 1.52 ;
 RECT 10.45 1.66 10.59 2.145 ;
 RECT 10.975 0.525 11.115 1.52 ;
 RECT 10.975 1.66 11.115 2.11 ;
 RECT 3.8 0.895 7.485 1.035 ;
 RECT 7.255 1.035 7.485 1.105 ;
 RECT 3.8 0.66 3.94 0.895 ;
 RECT 3.34 0.52 3.94 0.66 ;
 RECT 13.775 1.23 13.915 1.42 ;
 RECT 11.925 1.09 13.915 1.23 ;
 RECT 11.925 0.385 12.065 1.09 ;
 RECT 9.915 0.385 10.055 0.895 ;
 RECT 9.91 0.255 12.065 0.385 ;
 RECT 9.91 0.245 12.06 0.255 ;
 RECT 9.915 0.22 10.055 0.245 ;
 RECT 9 0.895 10.055 1.035 ;
 RECT 9 0.745 9.14 0.895 ;
 RECT 4.08 0.605 9.14 0.745 ;
 RECT 4.08 0.485 4.395 0.605 ;
 RECT 14.12 1.39 14.35 1.42 ;
 RECT 13.775 1.42 14.35 1.56 ;
 RECT 14.12 1.56 14.35 1.6 ;
 RECT 2.655 1.67 2.795 1.82 ;
 RECT 2.655 1.96 2.795 2.25 ;
 RECT 2.655 0.715 2.795 1.44 ;
 RECT 2.655 1.44 2.91 1.67 ;
 RECT 2.655 0.505 2.9 0.715 ;
 RECT 2.525 1.82 2.795 1.96 ;
 RECT 0.585 1.335 0.725 2.11 ;
 RECT 0.585 2.25 0.725 2.255 ;
 RECT 0.585 0.875 0.725 1.195 ;
 RECT 0.585 2.11 1.01 2.25 ;
 RECT 0.585 0.735 1.01 0.875 ;
 RECT 0.585 1.195 1.695 1.335 ;
 RECT 1.555 0.6 1.695 1.195 ;
 RECT 3.05 0.36 3.19 1.96 ;
 RECT 2.285 0.36 2.425 0.46 ;
 RECT 2.94 1.96 3.21 2.1 ;
 RECT 1.555 0.46 2.425 0.6 ;
 RECT 2.285 0.22 3.19 0.36 ;
 RECT 12.895 1.895 13.035 2.39 ;
 RECT 16.835 2.205 16.975 2.39 ;
 RECT 12.895 2.39 16.975 2.53 ;
 RECT 11.77 1.755 13.035 1.895 ;
 RECT 11.77 1.895 11.91 2.34 ;
 RECT 10.5 2.3 10.73 2.34 ;
 RECT 10.5 2.48 10.73 2.51 ;
 RECT 10.5 2.34 11.91 2.48 ;
 RECT 16.835 2.065 23.055 2.205 ;
 RECT 22.915 2.205 23.055 2.52 ;
 RECT 27.255 2.48 27.395 2.52 ;
 RECT 22.915 2.52 27.395 2.66 ;
 RECT 27.255 2.27 27.485 2.48 ;
 RECT 16.335 1.7 16.63 1.84 ;
 RECT 16.335 1.84 16.475 2.075 ;
 RECT 15.64 1.84 15.78 2.075 ;
 RECT 15.445 1.7 15.78 1.84 ;
 RECT 15.64 2.075 16.475 2.215 ;
 RECT 16.53 1.055 16.67 1.245 ;
 RECT 15.97 1.385 16.11 1.625 ;
 RECT 15.97 1.245 17.04 1.385 ;
 RECT 16.81 1.385 17.04 1.455 ;
 RECT 16.5 0.915 16.8 1.055 ;
 RECT 15.94 1.625 16.195 1.92 ;
 RECT 13.175 1.56 13.315 2.11 ;
 RECT 13.175 2.11 15.5 2.245 ;
 RECT 13.175 2.245 15.495 2.25 ;
 RECT 15.27 2.035 15.5 2.11 ;
 RECT 12.125 1.405 12.355 1.42 ;
 RECT 12.125 1.56 12.355 1.615 ;
 RECT 12.125 1.42 13.315 1.56 ;
 RECT 8.65 1.685 9.225 1.775 ;
 RECT 9.085 1.335 9.225 1.635 ;
 RECT 8.49 1.635 9.225 1.685 ;
 RECT 8.65 1.04 8.79 1.475 ;
 RECT 8.49 1.475 8.79 1.635 ;
 RECT 8.65 1.775 8.79 2.18 ;
 RECT 9.085 1.195 9.435 1.335 ;
 RECT 8.58 0.9 8.855 1.04 ;
 RECT 3.8 1.225 7.115 1.25 ;
 RECT 6.41 1.365 6.55 2.25 ;
 RECT 3.8 1.365 4.14 1.4 ;
 RECT 3.8 1.18 3.94 1.225 ;
 RECT 3.8 1.4 3.94 1.45 ;
 RECT 3.8 1.25 7.865 1.365 ;
 RECT 7.725 0.885 7.865 0.9 ;
 RECT 7.725 1.04 7.865 1.25 ;
 RECT 6.975 1.365 7.865 1.39 ;
 RECT 7.725 1.39 7.865 2.215 ;
 RECT 7.66 0.9 7.935 1.04 ;
 RECT 4.85 2.1 5.125 2.245 ;
 RECT 3.905 1.96 5.125 2.1 ;
 RECT 3.52 1.79 5.175 1.815 ;
 RECT 3.52 1.815 3.71 1.93 ;
 RECT 3.52 0.805 3.66 1.675 ;
 RECT 3.43 1.93 3.71 2.07 ;
 RECT 3.52 1.675 6.22 1.79 ;
 RECT 4.995 1.65 6.22 1.675 ;
 RECT 5.985 1.615 6.215 1.65 ;
 RECT 5.985 1.79 6.215 1.825 ;
 RECT 1.795 1.63 1.935 1.99 ;
 END
END RDFFSRASX2

MACRO RDFFNSRASRQX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.84 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.895 0.52 21.265 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.125 1.435 26.465 1.8 ;
 RECT 24.445 1.99 26.31 2.13 ;
 RECT 22.215 2.22 24.585 2.36 ;
 RECT 26.17 1.8 26.31 1.99 ;
 RECT 24.445 1.435 24.585 1.99 ;
 RECT 22.215 1.39 22.355 2.22 ;
 RECT 23.6 1.37 23.74 2.22 ;
 RECT 24.445 2.13 24.585 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.17 1.135 0.465 1.405 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.825 0.08 2.105 0.295 ;
 RECT 24.565 0.08 24.805 0.26 ;
 RECT 5.755 0.31 6.045 0.45 ;
 RECT 13.365 0.275 14.39 0.415 ;
 RECT 9.44 0.615 9.71 0.755 ;
 RECT 14.25 0.75 15.195 0.89 ;
 RECT 0 -0.08 27.84 0.08 ;
 RECT 1.305 0.08 1.445 0.97 ;
 RECT 4.65 0.08 4.885 0.46 ;
 RECT 0.335 0.08 0.475 0.775 ;
 RECT 19.37 0.08 19.51 0.82 ;
 RECT 22.215 0.08 22.355 0.36 ;
 RECT 23.43 0.08 23.57 0.35 ;
 RECT 5.835 0.08 5.975 0.31 ;
 RECT 13.365 0.415 13.505 0.945 ;
 RECT 13.365 0.08 13.505 0.275 ;
 RECT 9.505 0.08 9.645 0.615 ;
 RECT 15.055 0.89 15.195 1.11 ;
 RECT 14.25 0.415 14.39 0.75 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 19.225 2.6 19.49 2.8 ;
 RECT 9.25 2.215 9.525 2.355 ;
 RECT 0 2.8 27.84 2.96 ;
 RECT 1.98 2.34 2.23 2.8 ;
 RECT 0.335 1.74 0.475 2.8 ;
 RECT 1.305 1.98 1.445 2.8 ;
 RECT 5.835 1.98 5.975 2.8 ;
 RECT 6.865 2 7.005 2.8 ;
 RECT 5.355 2.07 5.495 2.8 ;
 RECT 12.275 2.335 12.545 2.8 ;
 RECT 9.315 2.355 9.455 2.8 ;
 RECT 9.315 2.195 9.455 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.15 1.475 1.59 1.76 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.44 1.145 18.95 1.405 ;
 RECT 18.81 0.51 18.95 1.145 ;
 RECT 19.87 1.905 20.01 1.91 ;
 RECT 18.81 1.765 20.01 1.905 ;
 RECT 19.87 0.56 20.01 1.765 ;
 RECT 18.81 1.905 18.95 1.915 ;
 RECT 18.81 1.405 18.95 1.765 ;
 END
 ANTENNADIFFAREA 0.787 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.73 2.255 10.04 2.465 ;
 RECT 9.765 2.12 10.04 2.255 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.035 0.745 4.36 0.765 ;
 RECT 4.035 0.485 4.36 0.605 ;
 RECT 8.965 0.91 10.02 1.05 ;
 RECT 9.875 0.245 12.025 0.255 ;
 RECT 9.875 0.255 12.03 0.385 ;
 RECT 11.89 1.09 13.88 1.23 ;
 RECT 14.085 1.56 14.315 1.6 ;
 RECT 13.74 1.42 14.315 1.56 ;
 RECT 14.085 1.39 14.315 1.42 ;
 RECT 4.035 0.605 9.105 0.745 ;
 RECT 8.965 0.745 9.105 0.91 ;
 RECT 11.89 0.385 12.03 1.09 ;
 RECT 9.88 0.385 10.02 0.91 ;
 RECT 13.74 1.23 13.88 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.23 1.795 7.49 2.05 ;
 RECT 6.655 1.655 7.49 1.795 ;
 RECT 6.655 1.795 6.885 1.83 ;
 RECT 6.655 1.62 6.885 1.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 OBS
 LAYER PO ;
 RECT 20.255 0.22 20.485 0.275 ;
 RECT 20.255 0.375 20.485 0.43 ;
 RECT 19.65 0.275 20.485 0.375 ;
 RECT 14.22 0.73 14.32 1.39 ;
 RECT 14.085 1.39 14.32 1.6 ;
 RECT 14.22 1.6 14.32 2.39 ;
 RECT 2.405 0.285 2.505 1.52 ;
 RECT 1.905 1.52 2.505 1.62 ;
 RECT 2.405 0.185 11.295 0.195 ;
 RECT 4.46 0.095 11.295 0.185 ;
 RECT 2.405 0.195 4.56 0.285 ;
 RECT 11.195 0.195 11.295 1.29 ;
 RECT 12.09 1.39 12.285 1.405 ;
 RECT 3.225 1.565 3.325 2.675 ;
 RECT 2.34 1.62 2.44 2.675 ;
 RECT 1.905 1.44 2.15 1.52 ;
 RECT 1.905 1.62 2.15 1.69 ;
 RECT 4.46 0.285 4.56 1.24 ;
 RECT 11.195 1.29 12.285 1.39 ;
 RECT 2.34 2.675 3.325 2.775 ;
 RECT 12.09 1.405 12.32 1.615 ;
 RECT 22.475 1.245 22.575 2.02 ;
 RECT 22.345 1.035 22.575 1.245 ;
 RECT 12.585 0.105 15.41 0.205 ;
 RECT 12.585 0.205 12.685 1.91 ;
 RECT 15.31 0.205 15.41 1.265 ;
 RECT 11.765 1.71 11.865 1.91 ;
 RECT 10.68 1.61 11.865 1.71 ;
 RECT 10.68 0.475 10.78 1.61 ;
 RECT 11.23 1.71 11.33 2.425 ;
 RECT 7.345 0.475 7.445 0.895 ;
 RECT 11.765 1.91 12.685 2.01 ;
 RECT 7.345 0.375 10.78 0.475 ;
 RECT 7.22 0.895 7.45 1.105 ;
 RECT 12.895 0.455 14.825 0.535 ;
 RECT 14.595 0.535 14.825 0.6 ;
 RECT 14.595 0.39 14.825 0.435 ;
 RECT 12.975 0.435 14.825 0.455 ;
 RECT 12.895 0.535 13.125 0.665 ;
 RECT 13.75 0.535 13.98 0.835 ;
 RECT 13.75 0.835 13.85 2.39 ;
 RECT 22.78 0.215 22.88 0.995 ;
 RECT 22.78 0.995 23.02 1.205 ;
 RECT 22.78 1.205 22.88 2 ;
 RECT 25.175 0.375 25.275 0.99 ;
 RECT 25.175 0.99 25.425 1.2 ;
 RECT 25.175 1.2 25.275 2.27 ;
 RECT 25.175 2.27 25.46 2.48 ;
 RECT 10.16 0.655 10.26 2.305 ;
 RECT 10.465 2.3 10.695 2.305 ;
 RECT 10.465 2.405 10.695 2.51 ;
 RECT 10.16 2.305 10.695 2.405 ;
 RECT 22 0.21 22.1 0.755 ;
 RECT 22 0.855 22.1 2.2 ;
 RECT 24.865 1.125 24.965 2.2 ;
 RECT 21.035 0.755 22.57 0.84 ;
 RECT 21.035 0.84 22.565 0.855 ;
 RECT 22.47 0.215 22.57 0.755 ;
 RECT 21.035 0.595 21.265 0.755 ;
 RECT 22 2.2 24.965 2.3 ;
 RECT 23.69 1.06 23.79 1.14 ;
 RECT 23.69 0.38 23.79 0.96 ;
 RECT 23.69 1.14 23.96 1.24 ;
 RECT 23.86 1.24 23.96 1.84 ;
 RECT 23.27 0.935 23.5 0.96 ;
 RECT 23.27 0.96 23.79 1.06 ;
 RECT 23.27 1.06 23.5 1.145 ;
 RECT 24.055 0.22 24.285 0.28 ;
 RECT 24.055 0.38 24.285 0.43 ;
 RECT 23.69 0.28 24.285 0.38 ;
 RECT 7.945 1.575 8.045 2.485 ;
 RECT 8.455 1.575 8.685 1.685 ;
 RECT 7.945 1.475 8.685 1.575 ;
 RECT 25.875 0.195 25.975 2.665 ;
 RECT 24.865 0.095 25.975 0.195 ;
 RECT 21.24 1.245 21.34 2.665 ;
 RECT 24.865 0.195 24.965 0.945 ;
 RECT 21.24 1.2 21.525 1.245 ;
 RECT 21.295 1.035 21.525 1.1 ;
 RECT 21.24 2.665 25.975 2.765 ;
 RECT 21.24 1.1 21.57 1.2 ;
 RECT 12.17 0.795 12.335 0.925 ;
 RECT 11.49 0.885 11.72 0.925 ;
 RECT 11.49 1.025 11.72 1.095 ;
 RECT 11.49 0.925 12.335 1.025 ;
 RECT 12.17 0.585 12.4 0.795 ;
 RECT 3.26 0.705 3.36 1.165 ;
 RECT 2.83 1.27 2.93 1.445 ;
 RECT 3.26 0.47 3.555 0.705 ;
 RECT 2.83 1.17 3.37 1.265 ;
 RECT 2.83 1.265 3.205 1.27 ;
 RECT 3.06 1.165 3.37 1.17 ;
 RECT 2.685 1.445 2.93 1.69 ;
 RECT 4.16 0.715 4.26 1.61 ;
 RECT 4.195 1.71 4.295 2.48 ;
 RECT 4.16 1.61 4.295 1.71 ;
 RECT 4.04 0.485 4.28 0.715 ;
 RECT 9.765 0.655 9.865 1.235 ;
 RECT 9.15 1.335 9.38 1.475 ;
 RECT 9.15 1.235 9.865 1.335 ;
 RECT 1.565 0.49 1.665 1.495 ;
 RECT 1.37 1.495 1.665 1.745 ;
 RECT 1.565 1.745 1.665 2.37 ;
 RECT 3.72 1.33 3.86 1.475 ;
 RECT 3.72 1.71 3.82 2.475 ;
 RECT 3.76 0.65 3.86 1.33 ;
 RECT 3.72 1.475 3.95 1.71 ;
 RECT 1.09 0.425 1.19 1.16 ;
 RECT 1.09 1.26 1.19 2.465 ;
 RECT 0.205 1.26 0.435 1.38 ;
 RECT 0.2 1.16 1.19 1.26 ;
 RECT 8.87 0.655 8.97 1.18 ;
 RECT 8.87 1.28 8.97 1.655 ;
 RECT 7.955 0.66 8.055 1.18 ;
 RECT 8.87 1.655 9.83 1.755 ;
 RECT 9.73 1.755 9.83 2.255 ;
 RECT 8.87 1.755 8.97 2.51 ;
 RECT 7.955 1.18 8.97 1.28 ;
 RECT 9.73 2.255 9.96 2.465 ;
 RECT 16.19 0.77 16.29 2.155 ;
 RECT 16.19 0.55 16.29 0.56 ;
 RECT 16.19 0.56 16.445 0.77 ;
 RECT 16.76 0.095 16.99 0.43 ;
 RECT 16.825 0.43 16.925 1.245 ;
 RECT 16.775 1.245 17.005 1.455 ;
 RECT 4.98 2.445 5.24 2.655 ;
 RECT 5.14 1.79 5.24 2.445 ;
 RECT 15.25 1.445 15.35 2.035 ;
 RECT 15.235 2.035 15.465 2.245 ;
 RECT 15.72 0.55 15.82 2.69 ;
 RECT 6.65 1.58 6.75 1.62 ;
 RECT 6.39 1.01 6.49 1.48 ;
 RECT 6.65 1.83 6.75 2.69 ;
 RECT 6.65 1.62 6.885 1.83 ;
 RECT 6.39 1.48 6.75 1.58 ;
 RECT 6.65 2.69 15.82 2.79 ;
 RECT 6.09 0.98 6.19 1.615 ;
 RECT 5.95 1.615 6.19 1.825 ;
 RECT 6.09 1.825 6.19 2.51 ;
 RECT 19.07 1.25 19.32 1.33 ;
 RECT 19.07 1.33 19.75 1.43 ;
 RECT 19.07 1.43 19.32 1.46 ;
 RECT 19.65 0.375 19.75 1.33 ;
 RECT 19.07 0.385 19.17 1.25 ;
 RECT 19.07 1.46 19.17 2.74 ;
 RECT 19.65 1.43 19.75 2.73 ;
 LAYER CO ;
 RECT 7.695 2.015 7.825 2.145 ;
 RECT 23.435 0.12 23.565 0.25 ;
 RECT 23 1.485 23.13 1.615 ;
 RECT 25.395 1.465 25.525 1.595 ;
 RECT 15.94 1.705 16.07 1.835 ;
 RECT 25.395 0.595 25.525 0.725 ;
 RECT 3.77 1.525 3.9 1.655 ;
 RECT 9.32 2.225 9.45 2.355 ;
 RECT 19.29 2.64 19.42 2.77 ;
 RECT 0.84 2.115 0.97 2.245 ;
 RECT 19.875 0.63 20.005 0.76 ;
 RECT 23.94 0.595 24.07 0.725 ;
 RECT 3.375 0.525 3.505 0.655 ;
 RECT 4.42 1.825 4.55 1.955 ;
 RECT 16.415 1.705 16.545 1.835 ;
 RECT 24.08 1.405 24.21 1.535 ;
 RECT 7.7 0.905 7.83 1.035 ;
 RECT 5.84 0.315 5.97 0.445 ;
 RECT 8.175 0.905 8.305 1.035 ;
 RECT 11.45 0.595 11.58 0.725 ;
 RECT 9.51 0.62 9.64 0.75 ;
 RECT 23.605 1.445 23.735 1.575 ;
 RECT 0.34 1.825 0.47 1.955 ;
 RECT 14.475 1.035 14.605 1.165 ;
 RECT 15.06 0.91 15.19 1.04 ;
 RECT 6.87 2.11 7 2.24 ;
 RECT 19.375 0.62 19.505 0.75 ;
 RECT 5.36 2.135 5.49 2.265 ;
 RECT 2.975 2.105 3.105 2.235 ;
 RECT 3.94 2.11 4.07 2.24 ;
 RECT 1.895 0.145 2.025 0.275 ;
 RECT 10.945 1.9 11.075 2.03 ;
 RECT 0.34 2.345 0.47 2.475 ;
 RECT 2.05 2.345 2.18 2.475 ;
 RECT 23 0.435 23.13 0.565 ;
 RECT 6.65 1.23 6.78 1.36 ;
 RECT 15.47 1.705 15.6 1.835 ;
 RECT 5.84 2.075 5.97 2.205 ;
 RECT 0.255 1.21 0.385 1.34 ;
 RECT 9.78 2.295 9.91 2.425 ;
 RECT 19.14 1.29 19.27 1.42 ;
 RECT 16.825 1.285 16.955 1.415 ;
 RECT 14.645 0.43 14.775 0.56 ;
 RECT 16.265 0.6 16.395 0.73 ;
 RECT 16.81 0.26 16.94 0.39 ;
 RECT 5.03 2.485 5.16 2.615 ;
 RECT 15.285 2.075 15.415 2.205 ;
 RECT 6.705 1.66 6.835 1.79 ;
 RECT 6 1.655 6.13 1.785 ;
 RECT 20.305 0.26 20.435 0.39 ;
 RECT 25.245 1.03 25.375 1.16 ;
 RECT 12.945 0.495 13.075 0.625 ;
 RECT 14.135 1.43 14.265 1.56 ;
 RECT 12.22 0.625 12.35 0.755 ;
 RECT 12.14 1.445 12.27 1.575 ;
 RECT 22.395 1.075 22.525 1.205 ;
 RECT 7.27 0.935 7.4 1.065 ;
 RECT 23.32 0.975 23.45 1.105 ;
 RECT 13.8 0.665 13.93 0.795 ;
 RECT 22.84 1.035 22.97 1.165 ;
 RECT 25.28 2.31 25.41 2.44 ;
 RECT 10.515 2.34 10.645 2.47 ;
 RECT 21.085 0.635 21.215 0.765 ;
 RECT 24.105 0.26 24.235 0.39 ;
 RECT 8.505 1.515 8.635 1.645 ;
 RECT 21.345 1.075 21.475 1.205 ;
 RECT 11.54 0.925 11.67 1.055 ;
 RECT 24.45 1.49 24.58 1.62 ;
 RECT 3.01 0.88 3.14 1.01 ;
 RECT 11.45 1.87 11.58 2 ;
 RECT 4.89 2.11 5.02 2.24 ;
 RECT 4.705 0.32 4.835 0.45 ;
 RECT 22.22 0.135 22.35 0.265 ;
 RECT 1.965 1.495 2.095 1.625 ;
 RECT 1.915 0.745 2.045 0.875 ;
 RECT 1.785 1.995 1.915 2.125 ;
 RECT 8.62 1.995 8.75 2.125 ;
 RECT 0.34 0.59 0.47 0.72 ;
 RECT 8.175 2.07 8.305 2.2 ;
 RECT 10.945 0.595 11.075 0.725 ;
 RECT 2.74 1.49 2.87 1.62 ;
 RECT 9.2 1.28 9.33 1.41 ;
 RECT 18.815 1.725 18.945 1.855 ;
 RECT 0.34 2.085 0.47 2.215 ;
 RECT 6.38 2.045 6.51 2.175 ;
 RECT 1.43 1.55 1.56 1.68 ;
 RECT 3.48 0.88 3.61 1.01 ;
 RECT 13.5 1.835 13.63 1.965 ;
 RECT 13.37 0.765 13.5 0.895 ;
 RECT 1.31 0.74 1.44 0.87 ;
 RECT 24.615 0.12 24.745 0.25 ;
 RECT 4.095 0.53 4.225 0.66 ;
 RECT 18.815 0.62 18.945 0.75 ;
 RECT 12.345 2.38 12.475 2.51 ;
 RECT 8.62 0.905 8.75 1.035 ;
 RECT 21.75 1.425 21.88 1.555 ;
 RECT 0.34 0.33 0.47 0.46 ;
 RECT 16.535 0.92 16.665 1.05 ;
 RECT 22.22 1.475 22.35 1.605 ;
 RECT 10.42 0.875 10.55 1.005 ;
 RECT 2.625 0.79 2.755 0.92 ;
 RECT 14.44 1.835 14.57 1.965 ;
 RECT 3.47 2.07 3.6 2.2 ;
 RECT 26.175 1.475 26.305 1.605 ;
 RECT 19.875 1.71 20.005 1.84 ;
 RECT 0.84 0.74 0.97 0.87 ;
 RECT 2.56 1.825 2.69 1.955 ;
 RECT 10.42 1.945 10.55 2.075 ;
 RECT 1.31 2.05 1.44 2.18 ;
 RECT 21.5 0.505 21.63 0.635 ;
 LAYER M1 ;
 RECT 4.43 1.365 4.57 1.5 ;
 RECT 3.6 1.64 4.105 1.675 ;
 RECT 3.6 1.5 4.57 1.64 ;
 RECT 7.69 1.04 7.83 1.25 ;
 RECT 7.69 1.39 7.83 2.215 ;
 RECT 7.69 0.885 7.83 0.9 ;
 RECT 4.43 1.25 7.83 1.365 ;
 RECT 6.94 1.365 7.83 1.39 ;
 RECT 7.625 0.9 7.9 1.04 ;
 RECT 23.935 0.73 24.075 1.04 ;
 RECT 24.075 1.18 24.215 1.605 ;
 RECT 23.87 0.59 24.145 0.73 ;
 RECT 25.195 0.99 25.425 1.04 ;
 RECT 23.935 1.04 25.425 1.18 ;
 RECT 25.195 1.18 25.425 1.2 ;
 RECT 24.055 0.29 24.425 0.43 ;
 RECT 24.285 0.43 24.425 0.71 ;
 RECT 24.055 0.22 24.285 0.29 ;
 RECT 25.705 0.85 25.845 1.385 ;
 RECT 25.39 1.525 25.53 1.73 ;
 RECT 24.285 0.71 25.845 0.85 ;
 RECT 25.39 0.51 25.53 0.71 ;
 RECT 25.39 1.385 25.845 1.525 ;
 RECT 21.295 1.225 21.525 1.245 ;
 RECT 21.295 1.195 21.885 1.225 ;
 RECT 21.435 1.015 21.745 1.035 ;
 RECT 21.295 1.035 21.745 1.055 ;
 RECT 21.57 0.64 21.71 1.015 ;
 RECT 21.745 1.225 21.885 1.75 ;
 RECT 21.45 0.5 21.71 0.64 ;
 RECT 22.345 1.035 22.575 1.055 ;
 RECT 22.345 1.195 22.575 1.245 ;
 RECT 21.295 1.055 22.575 1.195 ;
 RECT 23.315 1.145 23.455 1.345 ;
 RECT 22.995 1.485 23.135 1.76 ;
 RECT 23.315 0.73 23.455 0.935 ;
 RECT 22.995 0.355 23.135 0.59 ;
 RECT 22.995 1.345 23.455 1.485 ;
 RECT 23.27 0.935 23.5 1.145 ;
 RECT 22.995 0.59 23.455 0.73 ;
 RECT 20.255 0.36 20.485 0.43 ;
 RECT 21.85 0.36 21.99 0.565 ;
 RECT 20.255 0.22 21.99 0.36 ;
 RECT 22.59 0.705 22.73 0.75 ;
 RECT 22.715 0.995 23.02 1.205 ;
 RECT 22.715 0.89 22.855 0.995 ;
 RECT 22.59 0.75 22.855 0.89 ;
 RECT 21.85 0.565 22.73 0.705 ;
 RECT 18.41 0.36 18.55 0.635 ;
 RECT 15.49 0.635 18.55 0.775 ;
 RECT 14.47 1.545 14.61 1.83 ;
 RECT 14.47 1.17 14.61 1.405 ;
 RECT 13.425 1.83 14.675 1.97 ;
 RECT 14.4 1.03 14.68 1.17 ;
 RECT 15.49 0.775 15.63 1.405 ;
 RECT 16.215 0.56 16.445 0.635 ;
 RECT 14.47 1.405 15.63 1.545 ;
 RECT 19.09 0.36 19.23 1.25 ;
 RECT 19.09 1.25 19.32 1.46 ;
 RECT 18.41 0.22 19.23 0.36 ;
 RECT 14.595 0.28 16.99 0.42 ;
 RECT 14.595 0.42 14.825 0.6 ;
 RECT 16.76 0.22 16.99 0.28 ;
 RECT 16.76 0.42 16.99 0.43 ;
 RECT 11.445 0.525 11.585 0.885 ;
 RECT 11.445 1.095 11.585 2.065 ;
 RECT 11.445 0.885 11.72 1.095 ;
 RECT 8.965 2.055 9.105 2.34 ;
 RECT 8.17 2.34 9.105 2.48 ;
 RECT 9.485 1.66 9.625 1.915 ;
 RECT 8.965 1.915 9.625 2.055 ;
 RECT 8.17 1.04 8.31 2.34 ;
 RECT 8.17 0.895 8.31 0.9 ;
 RECT 8.1 0.9 8.375 1.04 ;
 RECT 10.94 0.525 11.08 1.52 ;
 RECT 10.94 1.66 11.08 2.11 ;
 RECT 10.415 0.765 10.555 1.52 ;
 RECT 10.415 1.66 10.555 2.145 ;
 RECT 9.485 1.52 11.08 1.66 ;
 RECT 13.75 0.57 13.98 0.95 ;
 RECT 12.17 0.585 13.125 0.63 ;
 RECT 12.17 0.63 12.4 0.795 ;
 RECT 12.195 0.49 13.125 0.585 ;
 RECT 12.895 0.455 13.125 0.49 ;
 RECT 12.895 0.63 13.125 0.665 ;
 RECT 0.615 1.335 0.755 2.11 ;
 RECT 0.615 2.25 0.755 2.255 ;
 RECT 0.615 0.875 0.755 1.195 ;
 RECT 0.615 2.11 1.04 2.25 ;
 RECT 0.615 0.735 1.04 0.875 ;
 RECT 0.615 1.195 1.725 1.335 ;
 RECT 1.585 0.6 1.725 1.195 ;
 RECT 2.33 0.36 2.47 0.46 ;
 RECT 3.005 0.97 3.155 1.095 ;
 RECT 3.015 1.095 3.155 2.035 ;
 RECT 3.005 0.36 3.145 0.97 ;
 RECT 2.33 0.22 3.145 0.36 ;
 RECT 2.97 2.17 3.11 2.305 ;
 RECT 1.585 0.46 2.47 0.6 ;
 RECT 2.97 2.035 3.155 2.17 ;
 RECT 3.755 0.66 3.895 0.92 ;
 RECT 3.3 0.52 3.895 0.66 ;
 RECT 7.22 0.895 7.45 0.92 ;
 RECT 7.22 1.06 7.45 1.105 ;
 RECT 3.755 0.92 7.45 1.06 ;
 RECT 1.865 0.88 2.005 1.475 ;
 RECT 1.825 1.63 1.965 1.99 ;
 RECT 1.825 1.475 2.17 1.63 ;
 RECT 1.715 1.99 1.965 2.13 ;
 RECT 1.865 0.74 2.185 0.88 ;
 RECT 3.31 1.82 4.89 1.96 ;
 RECT 4.75 1.79 4.89 1.82 ;
 RECT 3.395 1.96 3.675 2.215 ;
 RECT 3.475 0.805 3.615 1.22 ;
 RECT 3.31 1.22 3.615 1.36 ;
 RECT 3.31 1.36 3.45 1.82 ;
 RECT 5.95 1.615 6.18 1.65 ;
 RECT 5.95 1.79 6.18 1.825 ;
 RECT 4.75 1.65 6.185 1.79 ;
 RECT 2.62 1.67 2.76 1.82 ;
 RECT 2.62 1.96 2.76 2.51 ;
 RECT 2.62 0.5 2.76 1.44 ;
 RECT 2.62 1.44 2.875 1.67 ;
 RECT 2.49 1.82 2.76 1.96 ;
 RECT 4.98 2.445 5.21 2.51 ;
 RECT 4.98 2.65 5.21 2.655 ;
 RECT 2.62 2.51 5.21 2.65 ;
 RECT 16.3 1.7 16.595 1.84 ;
 RECT 16.3 1.84 16.44 2.075 ;
 RECT 15.605 1.84 15.745 2.075 ;
 RECT 15.41 1.7 15.745 1.84 ;
 RECT 15.605 2.075 16.44 2.215 ;
 RECT 16.495 1.055 16.635 1.245 ;
 RECT 15.935 1.385 16.075 1.625 ;
 RECT 16.775 1.385 17.005 1.455 ;
 RECT 15.935 1.245 17.005 1.385 ;
 RECT 16.465 0.915 16.765 1.055 ;
 RECT 15.905 1.625 16.16 1.92 ;
 RECT 13.14 1.56 13.28 2.11 ;
 RECT 12.09 1.405 12.32 1.42 ;
 RECT 12.09 1.56 12.32 1.615 ;
 RECT 12.09 1.42 13.28 1.56 ;
 RECT 13.14 2.11 15.465 2.245 ;
 RECT 13.14 2.245 15.46 2.25 ;
 RECT 15.235 2.035 15.465 2.11 ;
 RECT 17.005 2.205 17.145 2.39 ;
 RECT 12.86 1.895 13 2.39 ;
 RECT 12.86 2.39 17.145 2.53 ;
 RECT 11.735 1.755 13 1.895 ;
 RECT 11.735 1.895 11.875 2.34 ;
 RECT 10.465 2.3 10.695 2.34 ;
 RECT 10.465 2.48 10.695 2.51 ;
 RECT 10.465 2.34 11.875 2.48 ;
 RECT 17.005 2.065 21.03 2.205 ;
 RECT 20.89 2.205 21.03 2.52 ;
 RECT 25.23 2.48 25.37 2.52 ;
 RECT 20.89 2.52 25.37 2.66 ;
 RECT 25.23 2.27 25.46 2.48 ;
 RECT 8.615 1.04 8.755 1.475 ;
 RECT 8.455 1.475 8.755 1.635 ;
 RECT 8.615 1.775 8.755 2.18 ;
 RECT 8.545 0.9 8.82 1.04 ;
 RECT 9.195 1.21 9.335 1.635 ;
 RECT 8.615 1.685 9.335 1.775 ;
 RECT 8.455 1.635 9.335 1.685 ;
 RECT 3.87 2.105 5.09 2.245 ;
 RECT 4.43 1.225 7.08 1.25 ;
 RECT 6.375 1.365 6.515 2.25 ;
 END
END RDFFNSRASRQX1

MACRO RDFFNSRASRQX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.84 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.895 0.51 21.265 0.89 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.125 1.435 26.465 1.8 ;
 RECT 24.445 1.99 26.31 2.13 ;
 RECT 22.215 2.22 24.585 2.36 ;
 RECT 26.17 1.8 26.31 1.99 ;
 RECT 24.445 1.435 24.585 1.99 ;
 RECT 22.215 1.39 22.355 2.22 ;
 RECT 23.6 1.37 23.74 2.22 ;
 RECT 24.445 2.13 24.585 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.18 1.15 0.465 1.4 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.825 0.08 2.105 0.295 ;
 RECT 24.565 0.08 24.805 0.26 ;
 RECT 5.755 0.31 6.045 0.45 ;
 RECT 13.365 0.275 14.39 0.415 ;
 RECT 9.44 0.615 9.71 0.755 ;
 RECT 14.25 0.75 15.195 0.89 ;
 RECT 0 -0.08 27.84 0.08 ;
 RECT 0.335 0.08 0.475 0.775 ;
 RECT 1.305 0.08 1.445 0.97 ;
 RECT 4.65 0.08 4.885 0.46 ;
 RECT 18.325 0.08 18.465 0.82 ;
 RECT 19.37 0.08 19.51 0.82 ;
 RECT 22.215 0.08 22.355 0.36 ;
 RECT 23.43 0.08 23.57 0.35 ;
 RECT 5.835 0.08 5.975 0.31 ;
 RECT 13.365 0.415 13.505 0.945 ;
 RECT 13.365 0.08 13.505 0.275 ;
 RECT 9.505 0.08 9.645 0.615 ;
 RECT 15.055 0.89 15.195 1.11 ;
 RECT 14.25 0.415 14.39 0.75 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 18.225 2.6 18.49 2.8 ;
 RECT 19.225 2.6 19.49 2.8 ;
 RECT 9.25 2.215 9.525 2.355 ;
 RECT 0 2.8 27.84 2.96 ;
 RECT 0.335 1.74 0.475 2.8 ;
 RECT 1.98 2.34 2.23 2.8 ;
 RECT 1.305 1.98 1.445 2.8 ;
 RECT 5.355 2.07 5.495 2.8 ;
 RECT 5.835 1.98 5.975 2.8 ;
 RECT 6.865 2 7.005 2.8 ;
 RECT 12.275 2.335 12.545 2.8 ;
 RECT 9.315 2.355 9.455 2.8 ;
 RECT 9.315 2.195 9.455 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 1.475 1.59 1.755 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.87 1.15 20.295 1.405 ;
 RECT 19.87 0.56 20.01 1.15 ;
 RECT 17.76 1.905 17.9 1.915 ;
 RECT 17.76 0.51 17.9 1.765 ;
 RECT 18.81 1.905 18.95 1.915 ;
 RECT 18.81 0.51 18.95 1.765 ;
 RECT 19.87 1.905 20.01 1.91 ;
 RECT 17.725 1.765 20.01 1.905 ;
 RECT 19.87 1.405 20.01 1.765 ;
 END
 ANTENNADIFFAREA 0.975 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.73 2.255 10.04 2.465 ;
 RECT 9.78 2.12 10.04 2.255 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.035 0.745 4.36 0.755 ;
 RECT 4.035 0.485 4.36 0.605 ;
 RECT 8.965 0.9 10.02 1.04 ;
 RECT 9.88 0.22 10.02 0.245 ;
 RECT 9.875 0.245 12.025 0.255 ;
 RECT 9.875 0.255 12.03 0.385 ;
 RECT 11.89 1.09 13.88 1.23 ;
 RECT 14.085 1.56 14.315 1.6 ;
 RECT 13.74 1.42 14.315 1.56 ;
 RECT 14.085 1.39 14.315 1.42 ;
 RECT 4.035 0.605 9.105 0.745 ;
 RECT 8.965 0.745 9.105 0.9 ;
 RECT 9.88 0.385 10.02 0.9 ;
 RECT 11.89 0.385 12.03 1.09 ;
 RECT 13.74 1.23 13.88 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.22 1.795 7.495 2.045 ;
 RECT 6.655 1.795 6.885 1.83 ;
 RECT 6.655 1.655 7.495 1.795 ;
 RECT 6.655 1.62 6.885 1.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 OBS
 LAYER PO ;
 RECT 20.255 0.22 20.485 0.275 ;
 RECT 20.255 0.375 20.485 0.43 ;
 RECT 19.65 0.275 20.485 0.375 ;
 RECT 14.22 0.73 14.32 1.39 ;
 RECT 14.085 1.39 14.32 1.6 ;
 RECT 14.22 1.6 14.32 2.39 ;
 RECT 2.405 0.285 2.505 1.52 ;
 RECT 1.905 1.52 2.505 1.62 ;
 RECT 2.405 0.185 11.295 0.195 ;
 RECT 4.46 0.095 11.295 0.185 ;
 RECT 2.405 0.195 4.56 0.285 ;
 RECT 11.195 0.195 11.295 1.29 ;
 RECT 12.09 1.39 12.285 1.405 ;
 RECT 3.225 1.565 3.325 2.675 ;
 RECT 2.34 1.62 2.44 2.675 ;
 RECT 1.905 1.44 2.15 1.52 ;
 RECT 1.905 1.62 2.15 1.69 ;
 RECT 4.46 0.285 4.56 1.24 ;
 RECT 11.195 1.29 12.285 1.39 ;
 RECT 2.34 2.675 3.325 2.775 ;
 RECT 12.09 1.405 12.32 1.615 ;
 RECT 22.475 1.245 22.575 2.02 ;
 RECT 22.345 1.035 22.575 1.245 ;
 RECT 12.585 0.105 15.41 0.205 ;
 RECT 12.585 0.205 12.685 1.91 ;
 RECT 15.31 0.205 15.41 1.265 ;
 RECT 11.765 1.71 11.865 1.91 ;
 RECT 10.68 1.61 11.865 1.71 ;
 RECT 10.68 0.475 10.78 1.61 ;
 RECT 11.23 1.71 11.33 2.425 ;
 RECT 7.345 0.475 7.445 0.895 ;
 RECT 11.765 1.91 12.685 2.01 ;
 RECT 7.345 0.375 10.78 0.475 ;
 RECT 7.22 0.895 7.45 1.105 ;
 RECT 12.895 0.455 14.825 0.535 ;
 RECT 14.595 0.535 14.825 0.6 ;
 RECT 14.595 0.39 14.825 0.435 ;
 RECT 12.975 0.435 14.825 0.455 ;
 RECT 12.895 0.535 13.125 0.665 ;
 RECT 13.75 0.535 13.98 0.835 ;
 RECT 13.75 0.835 13.85 2.39 ;
 RECT 22.78 0.215 22.88 0.995 ;
 RECT 22.78 0.995 23.02 1.205 ;
 RECT 22.78 1.205 22.88 2 ;
 RECT 25.175 0.375 25.275 0.99 ;
 RECT 25.175 0.99 25.425 1.2 ;
 RECT 25.175 1.2 25.275 2.27 ;
 RECT 25.175 2.27 25.46 2.48 ;
 RECT 10.16 0.655 10.26 2.305 ;
 RECT 10.465 2.3 10.695 2.305 ;
 RECT 10.465 2.405 10.695 2.51 ;
 RECT 10.16 2.305 10.695 2.405 ;
 RECT 22 0.21 22.1 0.755 ;
 RECT 22 0.855 22.1 2.2 ;
 RECT 24.865 1.125 24.965 2.2 ;
 RECT 21.035 0.755 22.57 0.84 ;
 RECT 21.035 0.84 22.565 0.855 ;
 RECT 22.47 0.215 22.57 0.755 ;
 RECT 21.035 0.595 21.265 0.755 ;
 RECT 22 2.2 24.965 2.3 ;
 RECT 23.69 1.06 23.79 1.14 ;
 RECT 23.69 0.38 23.79 0.96 ;
 RECT 23.69 1.14 23.96 1.24 ;
 RECT 23.86 1.24 23.96 1.84 ;
 RECT 23.27 0.935 23.5 0.96 ;
 RECT 23.27 0.96 23.79 1.06 ;
 RECT 23.27 1.06 23.5 1.145 ;
 RECT 24.055 0.22 24.285 0.28 ;
 RECT 24.055 0.38 24.285 0.43 ;
 RECT 23.69 0.28 24.285 0.38 ;
 RECT 7.945 1.575 8.045 2.485 ;
 RECT 8.455 1.575 8.685 1.685 ;
 RECT 7.945 1.475 8.685 1.575 ;
 RECT 25.875 0.195 25.975 2.665 ;
 RECT 24.865 0.095 25.975 0.195 ;
 RECT 21.24 1.245 21.34 2.665 ;
 RECT 24.865 0.195 24.965 0.945 ;
 RECT 21.24 1.2 21.525 1.245 ;
 RECT 21.295 1.035 21.525 1.1 ;
 RECT 21.24 2.665 25.975 2.765 ;
 RECT 21.24 1.1 21.57 1.2 ;
 RECT 12.17 0.795 12.335 0.925 ;
 RECT 11.49 0.885 11.72 0.925 ;
 RECT 11.49 1.025 11.72 1.095 ;
 RECT 11.49 0.925 12.335 1.025 ;
 RECT 12.17 0.585 12.4 0.795 ;
 RECT 3.26 0.705 3.36 1.165 ;
 RECT 2.83 1.27 2.93 1.445 ;
 RECT 3.26 0.47 3.555 0.705 ;
 RECT 2.83 1.17 3.37 1.265 ;
 RECT 2.83 1.265 3.205 1.27 ;
 RECT 3.06 1.165 3.37 1.17 ;
 RECT 2.685 1.445 2.93 1.69 ;
 RECT 4.16 0.715 4.26 1.61 ;
 RECT 4.195 1.71 4.295 2.48 ;
 RECT 4.16 1.61 4.295 1.71 ;
 RECT 4.04 0.485 4.28 0.715 ;
 RECT 9.765 0.655 9.865 1.205 ;
 RECT 9.15 1.305 9.38 1.475 ;
 RECT 9.15 1.205 9.865 1.305 ;
 RECT 1.565 0.49 1.665 1.495 ;
 RECT 1.37 1.495 1.665 1.745 ;
 RECT 1.565 1.745 1.665 2.37 ;
 RECT 3.72 1.37 3.86 1.475 ;
 RECT 3.72 1.33 3.85 1.37 ;
 RECT 3.72 1.71 3.82 2.475 ;
 RECT 3.75 0.65 3.85 1.33 ;
 RECT 3.72 1.475 3.95 1.71 ;
 RECT 0.85 0.27 1.19 0.52 ;
 RECT 1.09 0.52 1.19 1.16 ;
 RECT 1.09 1.26 1.19 2.465 ;
 RECT 0.21 1.26 0.44 1.38 ;
 RECT 0.21 1.16 1.19 1.26 ;
 RECT 8.87 0.655 8.97 1.18 ;
 RECT 8.87 1.28 8.97 1.655 ;
 RECT 7.955 0.66 8.055 1.18 ;
 RECT 8.87 1.655 9.83 1.755 ;
 RECT 9.73 1.755 9.83 2.255 ;
 RECT 8.87 1.755 8.97 2.51 ;
 RECT 7.955 1.18 8.97 1.28 ;
 RECT 9.73 2.255 9.96 2.465 ;
 RECT 16.19 0.77 16.29 2.155 ;
 RECT 16.19 0.55 16.29 0.56 ;
 RECT 16.19 0.56 16.445 0.77 ;
 RECT 16.825 0.43 16.925 1.245 ;
 RECT 16.775 1.245 17.005 1.455 ;
 RECT 16.76 0.22 16.99 0.43 ;
 RECT 4.98 2.445 5.24 2.655 ;
 RECT 5.14 1.79 5.24 2.445 ;
 RECT 15.25 1.445 15.35 2.035 ;
 RECT 15.235 2.035 15.465 2.245 ;
 RECT 15.72 0.55 15.82 2.69 ;
 RECT 6.65 1.58 6.75 1.62 ;
 RECT 6.39 1.01 6.49 1.48 ;
 RECT 6.65 1.83 6.75 2.69 ;
 RECT 6.65 1.62 6.885 1.83 ;
 RECT 6.39 1.48 6.75 1.58 ;
 RECT 6.65 2.69 15.82 2.79 ;
 RECT 6.09 0.98 6.19 1.615 ;
 RECT 5.95 1.615 6.19 1.825 ;
 RECT 6.09 1.825 6.19 2.51 ;
 RECT 17.265 1.33 19.75 1.43 ;
 RECT 17.265 1.265 17.495 1.33 ;
 RECT 18.015 1.43 18.115 2.74 ;
 RECT 19.65 0.375 19.75 1.33 ;
 RECT 18.015 0.385 18.115 1.33 ;
 RECT 17.265 1.43 17.495 1.475 ;
 RECT 18.595 1.43 18.695 2.73 ;
 RECT 18.595 0.385 18.695 1.33 ;
 RECT 19.07 0.385 19.17 1.33 ;
 RECT 19.07 1.43 19.17 2.74 ;
 RECT 19.65 1.43 19.75 2.73 ;
 LAYER CO ;
 RECT 24.45 1.49 24.58 1.62 ;
 RECT 3.01 0.88 3.14 1.01 ;
 RECT 11.45 1.87 11.58 2 ;
 RECT 4.89 2.11 5.02 2.24 ;
 RECT 4.705 0.32 4.835 0.45 ;
 RECT 16.415 1.705 16.545 1.835 ;
 RECT 24.08 1.405 24.21 1.535 ;
 RECT 7.7 0.905 7.83 1.035 ;
 RECT 0.91 0.325 1.04 0.455 ;
 RECT 5.84 0.315 5.97 0.445 ;
 RECT 8.175 0.905 8.305 1.035 ;
 RECT 11.45 0.595 11.58 0.725 ;
 RECT 9.51 0.62 9.64 0.75 ;
 RECT 23.605 1.445 23.735 1.575 ;
 RECT 0.34 1.825 0.47 1.955 ;
 RECT 14.475 1.035 14.605 1.165 ;
 RECT 15.06 0.91 15.19 1.04 ;
 RECT 6.87 2.11 7 2.24 ;
 RECT 19.375 0.62 19.505 0.75 ;
 RECT 5.36 2.135 5.49 2.265 ;
 RECT 2.975 2.105 3.105 2.235 ;
 RECT 3.94 2.11 4.07 2.24 ;
 RECT 1.895 0.145 2.025 0.275 ;
 RECT 10.945 1.9 11.075 2.03 ;
 RECT 0.34 2.345 0.47 2.475 ;
 RECT 2.05 2.345 2.18 2.475 ;
 RECT 23 0.435 23.13 0.565 ;
 RECT 6.65 1.23 6.78 1.36 ;
 RECT 15.47 1.705 15.6 1.835 ;
 RECT 5.84 2.075 5.97 2.205 ;
 RECT 3.48 0.88 3.61 1.01 ;
 RECT 13.5 1.835 13.63 1.965 ;
 RECT 0.26 1.21 0.39 1.34 ;
 RECT 9.78 2.295 9.91 2.425 ;
 RECT 17.315 1.305 17.445 1.435 ;
 RECT 16.825 1.285 16.955 1.415 ;
 RECT 14.645 0.43 14.775 0.56 ;
 RECT 16.265 0.6 16.395 0.73 ;
 RECT 16.81 0.26 16.94 0.39 ;
 RECT 5.03 2.485 5.16 2.615 ;
 RECT 15.285 2.075 15.415 2.205 ;
 RECT 6.705 1.66 6.835 1.79 ;
 RECT 6 1.655 6.13 1.785 ;
 RECT 20.305 0.26 20.435 0.39 ;
 RECT 25.245 1.03 25.375 1.16 ;
 RECT 12.945 0.495 13.075 0.625 ;
 RECT 14.135 1.43 14.265 1.56 ;
 RECT 12.22 0.625 12.35 0.755 ;
 RECT 12.14 1.445 12.27 1.575 ;
 RECT 22.395 1.075 22.525 1.205 ;
 RECT 7.27 0.935 7.4 1.065 ;
 RECT 23.32 0.975 23.45 1.105 ;
 RECT 13.8 0.665 13.93 0.795 ;
 RECT 22.84 1.035 22.97 1.165 ;
 RECT 25.28 2.31 25.41 2.44 ;
 RECT 10.515 2.34 10.645 2.47 ;
 RECT 21.085 0.635 21.215 0.765 ;
 RECT 24.105 0.26 24.235 0.39 ;
 RECT 8.505 1.515 8.635 1.645 ;
 RECT 21.345 1.075 21.475 1.205 ;
 RECT 11.54 0.925 11.67 1.055 ;
 RECT 22.22 0.135 22.35 0.265 ;
 RECT 1.965 1.495 2.095 1.625 ;
 RECT 1.915 0.745 2.045 0.875 ;
 RECT 1.785 1.995 1.915 2.125 ;
 RECT 8.62 1.995 8.75 2.125 ;
 RECT 0.34 0.59 0.47 0.72 ;
 RECT 8.175 2.07 8.305 2.2 ;
 RECT 10.945 0.595 11.075 0.725 ;
 RECT 2.74 1.49 2.87 1.62 ;
 RECT 9.2 1.28 9.33 1.41 ;
 RECT 18.815 1.725 18.945 1.855 ;
 RECT 0.34 2.085 0.47 2.215 ;
 RECT 6.38 2.045 6.51 2.175 ;
 RECT 1.43 1.55 1.56 1.68 ;
 RECT 18.29 2.64 18.42 2.77 ;
 RECT 18.33 0.62 18.46 0.75 ;
 RECT 17.765 1.725 17.895 1.855 ;
 RECT 17.765 0.62 17.895 0.75 ;
 RECT 13.37 0.765 13.5 0.895 ;
 RECT 1.31 0.74 1.44 0.87 ;
 RECT 24.615 0.12 24.745 0.25 ;
 RECT 4.095 0.53 4.225 0.66 ;
 RECT 18.815 0.62 18.945 0.75 ;
 RECT 12.345 2.38 12.475 2.51 ;
 RECT 8.62 0.905 8.75 1.035 ;
 RECT 21.75 1.425 21.88 1.555 ;
 RECT 0.34 0.33 0.47 0.46 ;
 RECT 16.535 0.92 16.665 1.05 ;
 RECT 22.22 1.475 22.35 1.605 ;
 RECT 10.42 0.875 10.55 1.005 ;
 RECT 2.625 0.79 2.755 0.92 ;
 RECT 14.44 1.835 14.57 1.965 ;
 RECT 3.47 2.07 3.6 2.2 ;
 RECT 26.175 1.475 26.305 1.605 ;
 RECT 19.875 1.71 20.005 1.84 ;
 RECT 0.84 0.74 0.97 0.87 ;
 RECT 2.56 1.825 2.69 1.955 ;
 RECT 10.42 1.945 10.55 2.075 ;
 RECT 1.31 2.05 1.44 2.18 ;
 RECT 21.5 0.505 21.63 0.635 ;
 RECT 7.695 2.015 7.825 2.145 ;
 RECT 23.435 0.12 23.565 0.25 ;
 RECT 23 1.485 23.13 1.615 ;
 RECT 25.395 1.465 25.525 1.595 ;
 RECT 15.94 1.705 16.07 1.835 ;
 RECT 25.395 0.595 25.525 0.725 ;
 RECT 3.77 1.525 3.9 1.655 ;
 RECT 9.32 2.225 9.45 2.355 ;
 RECT 19.29 2.64 19.42 2.77 ;
 RECT 0.84 2.115 0.97 2.245 ;
 RECT 19.875 0.63 20.005 0.76 ;
 RECT 23.94 0.595 24.07 0.725 ;
 RECT 3.375 0.525 3.505 0.655 ;
 RECT 4.42 1.825 4.55 1.955 ;
 LAYER M1 ;
 RECT 4.43 1.365 4.57 1.5 ;
 RECT 3.6 1.64 4.105 1.675 ;
 RECT 3.6 1.5 4.57 1.64 ;
 RECT 7.69 1.04 7.83 1.25 ;
 RECT 7.69 1.39 7.83 2.215 ;
 RECT 7.69 0.885 7.83 0.9 ;
 RECT 4.43 1.25 7.83 1.365 ;
 RECT 6.94 1.365 7.83 1.39 ;
 RECT 7.625 0.9 7.9 1.04 ;
 RECT 3.31 1.82 4.89 1.96 ;
 RECT 4.75 1.79 4.89 1.82 ;
 RECT 3.395 1.96 3.675 2.215 ;
 RECT 3.475 0.805 3.615 1.22 ;
 RECT 3.31 1.22 3.615 1.36 ;
 RECT 3.31 1.36 3.45 1.82 ;
 RECT 5.95 1.615 6.18 1.65 ;
 RECT 5.95 1.79 6.18 1.825 ;
 RECT 4.75 1.65 6.185 1.79 ;
 RECT 23.935 0.73 24.075 1.04 ;
 RECT 24.075 1.18 24.215 1.605 ;
 RECT 23.87 0.59 24.145 0.73 ;
 RECT 25.195 0.99 25.425 1.04 ;
 RECT 23.935 1.04 25.425 1.18 ;
 RECT 25.195 1.18 25.425 1.2 ;
 RECT 24.055 0.29 24.425 0.43 ;
 RECT 24.285 0.43 24.425 0.71 ;
 RECT 24.055 0.22 24.285 0.29 ;
 RECT 25.705 0.85 25.845 1.385 ;
 RECT 25.39 1.525 25.53 1.73 ;
 RECT 24.285 0.71 25.845 0.85 ;
 RECT 25.39 0.51 25.53 0.71 ;
 RECT 25.39 1.385 25.845 1.525 ;
 RECT 21.295 1.225 21.525 1.245 ;
 RECT 21.295 1.195 21.885 1.225 ;
 RECT 21.435 1.015 21.745 1.035 ;
 RECT 21.295 1.035 21.745 1.055 ;
 RECT 21.57 0.64 21.71 1.015 ;
 RECT 21.745 1.225 21.885 1.75 ;
 RECT 21.45 0.5 21.71 0.64 ;
 RECT 22.345 1.035 22.575 1.055 ;
 RECT 22.345 1.195 22.575 1.245 ;
 RECT 21.295 1.055 22.575 1.195 ;
 RECT 23.315 1.145 23.455 1.345 ;
 RECT 22.995 1.485 23.135 1.76 ;
 RECT 23.315 0.73 23.455 0.935 ;
 RECT 22.995 0.355 23.135 0.59 ;
 RECT 22.995 1.345 23.455 1.485 ;
 RECT 23.27 0.935 23.5 1.145 ;
 RECT 22.995 0.59 23.455 0.73 ;
 RECT 20.255 0.36 20.485 0.43 ;
 RECT 21.85 0.36 21.99 0.565 ;
 RECT 20.255 0.22 21.99 0.36 ;
 RECT 22.59 0.705 22.73 0.75 ;
 RECT 22.715 0.995 23.02 1.205 ;
 RECT 22.715 0.89 22.855 0.995 ;
 RECT 22.59 0.75 22.855 0.89 ;
 RECT 21.85 0.565 22.73 0.705 ;
 RECT 14.47 1.545 14.61 1.83 ;
 RECT 14.47 1.17 14.61 1.405 ;
 RECT 13.425 1.83 14.675 1.97 ;
 RECT 14.4 1.03 14.68 1.17 ;
 RECT 15.49 0.775 15.63 1.405 ;
 RECT 17.315 0.775 17.455 1.265 ;
 RECT 16.215 0.56 16.445 0.635 ;
 RECT 14.47 1.405 15.63 1.545 ;
 RECT 17.265 1.265 17.495 1.475 ;
 RECT 15.49 0.635 17.455 0.775 ;
 RECT 14.595 0.28 16.99 0.42 ;
 RECT 14.595 0.42 14.825 0.6 ;
 RECT 16.76 0.22 16.99 0.28 ;
 RECT 16.76 0.42 16.99 0.43 ;
 RECT 11.445 0.525 11.585 0.885 ;
 RECT 11.445 1.095 11.585 2.065 ;
 RECT 11.445 0.885 11.72 1.095 ;
 RECT 8.965 2.055 9.105 2.34 ;
 RECT 8.17 2.34 9.105 2.48 ;
 RECT 9.495 1.66 9.635 1.915 ;
 RECT 8.965 1.915 9.635 2.055 ;
 RECT 8.17 1.04 8.31 2.34 ;
 RECT 8.17 0.895 8.31 0.9 ;
 RECT 8.1 0.9 8.375 1.04 ;
 RECT 10.94 0.525 11.08 1.52 ;
 RECT 10.94 1.66 11.08 2.11 ;
 RECT 10.415 0.765 10.555 1.52 ;
 RECT 10.415 1.66 10.555 2.145 ;
 RECT 9.495 1.52 11.08 1.66 ;
 RECT 13.75 0.57 13.98 0.95 ;
 RECT 12.17 0.585 13.125 0.63 ;
 RECT 12.17 0.63 12.4 0.795 ;
 RECT 12.195 0.49 13.125 0.585 ;
 RECT 12.895 0.455 13.125 0.49 ;
 RECT 12.895 0.63 13.125 0.665 ;
 RECT 2.62 1.67 2.76 1.82 ;
 RECT 2.62 1.96 2.76 2.51 ;
 RECT 2.62 0.5 2.76 1.44 ;
 RECT 2.62 1.44 2.875 1.67 ;
 RECT 2.49 1.82 2.76 1.96 ;
 RECT 4.98 2.445 5.21 2.51 ;
 RECT 4.98 2.65 5.21 2.655 ;
 RECT 2.62 2.51 5.21 2.65 ;
 RECT 0.615 1.335 0.755 2.11 ;
 RECT 0.615 2.25 0.755 2.255 ;
 RECT 0.615 0.875 0.755 1.195 ;
 RECT 0.615 2.11 1.04 2.25 ;
 RECT 0.615 0.735 1.04 0.875 ;
 RECT 0.615 1.195 1.725 1.335 ;
 RECT 1.585 0.6 1.725 1.195 ;
 RECT 2.33 0.36 2.47 0.46 ;
 RECT 3.005 0.97 3.155 1.085 ;
 RECT 3.015 1.085 3.155 2.035 ;
 RECT 3.005 0.36 3.145 0.97 ;
 RECT 2.33 0.22 3.145 0.36 ;
 RECT 2.97 2.17 3.11 2.305 ;
 RECT 1.585 0.46 2.47 0.6 ;
 RECT 2.97 2.035 3.155 2.17 ;
 RECT 3.755 0.66 3.895 0.915 ;
 RECT 3.3 0.52 3.895 0.66 ;
 RECT 3.755 0.915 7.45 1.035 ;
 RECT 3.765 1.035 7.45 1.055 ;
 RECT 7.22 0.895 7.45 0.915 ;
 RECT 7.22 1.055 7.45 1.105 ;
 RECT 1.865 0.88 2.005 1.475 ;
 RECT 1.825 1.63 1.965 1.99 ;
 RECT 1.825 1.475 2.17 1.63 ;
 RECT 1.715 1.99 1.965 2.13 ;
 RECT 1.865 0.74 2.185 0.88 ;
 RECT 0.8 0.22 1.165 0.525 ;
 RECT 16.3 1.7 16.595 1.84 ;
 RECT 16.3 1.84 16.44 2.075 ;
 RECT 15.605 1.84 15.745 2.075 ;
 RECT 15.41 1.7 15.745 1.84 ;
 RECT 15.605 2.075 16.44 2.215 ;
 RECT 16.495 1.055 16.635 1.245 ;
 RECT 15.935 1.385 16.075 1.625 ;
 RECT 16.775 1.385 17.005 1.455 ;
 RECT 15.935 1.245 17.005 1.385 ;
 RECT 16.465 0.915 16.765 1.055 ;
 RECT 15.905 1.625 16.16 1.92 ;
 RECT 13.14 1.56 13.28 2.11 ;
 RECT 12.09 1.405 12.32 1.42 ;
 RECT 12.09 1.56 12.32 1.615 ;
 RECT 12.09 1.42 13.28 1.56 ;
 RECT 13.14 2.11 15.465 2.245 ;
 RECT 13.14 2.245 15.46 2.25 ;
 RECT 15.235 2.035 15.465 2.11 ;
 RECT 17.005 2.205 17.145 2.39 ;
 RECT 12.86 1.895 13 2.39 ;
 RECT 12.86 2.39 17.145 2.53 ;
 RECT 11.735 1.755 13 1.895 ;
 RECT 11.735 1.895 11.875 2.34 ;
 RECT 10.465 2.3 10.695 2.34 ;
 RECT 10.465 2.48 10.695 2.51 ;
 RECT 10.465 2.34 11.875 2.48 ;
 RECT 17.005 2.065 21.03 2.205 ;
 RECT 20.89 2.205 21.03 2.52 ;
 RECT 25.23 2.48 25.37 2.52 ;
 RECT 20.89 2.52 25.37 2.66 ;
 RECT 25.23 2.27 25.46 2.48 ;
 RECT 8.615 1.04 8.755 1.475 ;
 RECT 8.455 1.475 8.755 1.635 ;
 RECT 8.615 1.775 8.755 2.18 ;
 RECT 8.545 0.9 8.82 1.04 ;
 RECT 9.195 1.21 9.335 1.635 ;
 RECT 8.615 1.685 9.335 1.775 ;
 RECT 8.455 1.635 9.335 1.685 ;
 RECT 3.87 2.105 5.09 2.245 ;
 RECT 4.43 1.225 7.08 1.25 ;
 RECT 6.375 1.365 6.515 2.25 ;
 END
END RDFFNSRASRQX2

MACRO RDFFNSRASRX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 27.84 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.965 0.75 21.285 1.085 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 26.125 1.435 26.465 1.8 ;
 RECT 24.445 1.99 26.31 2.13 ;
 RECT 22.215 2.22 24.585 2.36 ;
 RECT 26.17 1.8 26.31 1.99 ;
 RECT 24.445 1.435 24.585 1.99 ;
 RECT 22.215 1.39 22.355 2.22 ;
 RECT 23.6 1.37 23.74 2.22 ;
 RECT 24.445 2.13 24.585 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.165 1.135 0.46 1.41 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.825 0.08 2.105 0.295 ;
 RECT 24.565 0.08 24.805 0.26 ;
 RECT 5.755 0.31 6.045 0.45 ;
 RECT 9.44 0.615 9.71 0.755 ;
 RECT 13.365 0.275 14.39 0.415 ;
 RECT 17.725 0.335 17.99 0.495 ;
 RECT 14.25 0.75 15.195 0.89 ;
 RECT 0 -0.08 27.84 0.08 ;
 RECT 0.335 0.08 0.475 0.775 ;
 RECT 1.305 0.08 1.445 0.97 ;
 RECT 4.65 0.08 4.885 0.46 ;
 RECT 19.37 0.08 19.51 0.82 ;
 RECT 22.215 0.08 22.355 0.36 ;
 RECT 23.43 0.08 23.57 0.35 ;
 RECT 5.835 0.08 5.975 0.31 ;
 RECT 9.505 0.08 9.645 0.615 ;
 RECT 13.365 0.415 13.505 0.945 ;
 RECT 13.365 0.08 13.505 0.275 ;
 RECT 17.78 0.08 17.92 0.335 ;
 RECT 15.055 0.89 15.195 1.11 ;
 RECT 14.25 0.415 14.39 0.75 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.155 1.155 17.43 1.445 ;
 RECT 17.29 0.915 17.43 1.155 ;
 RECT 18.295 1.84 18.435 1.885 ;
 RECT 18.295 0.915 18.435 1.7 ;
 RECT 17.29 1.84 17.43 1.885 ;
 RECT 17.29 1.7 18.435 1.84 ;
 RECT 17.29 1.445 17.43 1.7 ;
 END
 ANTENNADIFFAREA 0.7 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 17.635 2.6 17.9 2.8 ;
 RECT 19.225 2.6 19.49 2.8 ;
 RECT 9.25 2.215 9.525 2.355 ;
 RECT 0 2.8 27.84 2.96 ;
 RECT 0.335 1.74 0.475 2.8 ;
 RECT 1.98 2.34 2.23 2.8 ;
 RECT 5.355 2.07 5.495 2.8 ;
 RECT 1.305 1.98 1.445 2.8 ;
 RECT 5.835 1.98 5.975 2.8 ;
 RECT 6.865 2 7.005 2.8 ;
 RECT 12.275 2.335 12.545 2.8 ;
 RECT 9.315 2.355 9.455 2.8 ;
 RECT 9.315 2.195 9.455 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.155 1.475 1.59 1.73 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.81 0.51 18.95 1.48 ;
 RECT 18.76 1.48 19 1.765 ;
 RECT 18.81 1.905 18.95 1.915 ;
 RECT 18.81 1.775 20.01 1.905 ;
 RECT 19.87 1.905 20.01 1.91 ;
 RECT 19.87 0.56 20.01 1.765 ;
 RECT 18.76 1.765 20.01 1.775 ;
 END
 ANTENNADIFFAREA 0.568 ;
 END Q

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.73 2.255 10.04 2.465 ;
 RECT 9.77 2.12 10.04 2.255 ;
 RECT 9.77 2.465 10.04 2.47 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.035 0.745 4.36 0.76 ;
 RECT 4.035 0.485 4.36 0.605 ;
 RECT 8.965 0.9 10.02 1.04 ;
 RECT 9.88 0.22 10.02 0.245 ;
 RECT 9.875 0.245 12.025 0.255 ;
 RECT 9.875 0.255 12.03 0.385 ;
 RECT 11.89 1.09 13.88 1.23 ;
 RECT 14.085 1.56 14.315 1.6 ;
 RECT 13.74 1.42 14.315 1.56 ;
 RECT 14.085 1.39 14.315 1.42 ;
 RECT 4.035 0.605 9.105 0.745 ;
 RECT 8.965 0.745 9.105 0.9 ;
 RECT 9.88 0.385 10.02 0.9 ;
 RECT 11.89 0.385 12.03 1.09 ;
 RECT 13.74 1.23 13.88 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.23 1.795 7.49 2.05 ;
 RECT 6.655 1.795 6.885 1.83 ;
 RECT 6.655 1.655 7.49 1.795 ;
 RECT 6.655 1.62 6.885 1.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 OBS
 LAYER PO ;
 RECT 19.65 1.43 19.75 2.575 ;
 RECT 20.255 0.22 20.485 0.255 ;
 RECT 20.255 0.355 20.485 0.43 ;
 RECT 19.65 0.255 20.485 0.355 ;
 RECT 14.22 0.73 14.32 1.39 ;
 RECT 14.085 1.39 14.32 1.6 ;
 RECT 14.22 1.6 14.32 2.39 ;
 RECT 2.405 0.285 2.505 1.52 ;
 RECT 1.905 1.52 2.505 1.62 ;
 RECT 2.405 0.185 11.295 0.195 ;
 RECT 4.46 0.095 11.295 0.185 ;
 RECT 2.405 0.195 4.56 0.285 ;
 RECT 11.195 0.195 11.295 1.29 ;
 RECT 12.09 1.39 12.285 1.405 ;
 RECT 3.225 1.565 3.325 2.675 ;
 RECT 2.34 1.62 2.44 2.675 ;
 RECT 1.905 1.44 2.15 1.52 ;
 RECT 1.905 1.62 2.15 1.69 ;
 RECT 4.46 0.285 4.56 1.24 ;
 RECT 11.195 1.29 12.285 1.39 ;
 RECT 2.34 2.675 3.325 2.775 ;
 RECT 12.09 1.405 12.32 1.615 ;
 RECT 22.475 1.245 22.575 2.02 ;
 RECT 22.345 1.035 22.575 1.245 ;
 RECT 12.585 0.105 15.41 0.205 ;
 RECT 12.585 0.205 12.685 1.91 ;
 RECT 15.31 0.205 15.41 1.265 ;
 RECT 11.765 1.71 11.865 1.91 ;
 RECT 10.68 1.61 11.865 1.71 ;
 RECT 10.68 0.475 10.78 1.61 ;
 RECT 11.23 1.71 11.33 2.425 ;
 RECT 7.345 0.475 7.445 0.895 ;
 RECT 11.765 1.91 12.685 2.01 ;
 RECT 7.345 0.375 10.78 0.475 ;
 RECT 7.22 0.895 7.45 1.105 ;
 RECT 12.895 0.455 14.825 0.535 ;
 RECT 14.595 0.535 14.825 0.6 ;
 RECT 14.595 0.39 14.825 0.435 ;
 RECT 12.975 0.435 14.825 0.455 ;
 RECT 12.895 0.535 13.125 0.665 ;
 RECT 13.75 0.535 13.98 0.835 ;
 RECT 13.75 0.835 13.85 2.39 ;
 RECT 22.78 0.215 22.88 0.995 ;
 RECT 22.78 0.995 23.02 1.205 ;
 RECT 22.78 1.205 22.88 2 ;
 RECT 25.175 0.375 25.275 0.99 ;
 RECT 25.175 0.99 25.425 1.2 ;
 RECT 25.175 1.2 25.275 2.27 ;
 RECT 25.175 2.27 25.46 2.48 ;
 RECT 10.16 0.655 10.26 2.305 ;
 RECT 10.465 2.3 10.695 2.305 ;
 RECT 10.465 2.405 10.695 2.51 ;
 RECT 10.16 2.305 10.695 2.405 ;
 RECT 22 0.21 22.1 0.755 ;
 RECT 22 0.855 22.1 2.2 ;
 RECT 24.865 1.125 24.965 2.2 ;
 RECT 21.035 0.755 22.57 0.84 ;
 RECT 21.035 0.84 22.565 0.855 ;
 RECT 22.47 0.215 22.57 0.755 ;
 RECT 21.035 0.855 21.265 1.05 ;
 RECT 22 2.2 24.965 2.3 ;
 RECT 23.69 1.06 23.79 1.14 ;
 RECT 23.69 0.38 23.79 0.96 ;
 RECT 23.69 1.14 23.96 1.24 ;
 RECT 23.86 1.24 23.96 1.84 ;
 RECT 23.27 0.935 23.5 0.96 ;
 RECT 23.27 0.96 23.79 1.06 ;
 RECT 23.27 1.06 23.5 1.145 ;
 RECT 24.055 0.22 24.285 0.28 ;
 RECT 24.055 0.38 24.285 0.43 ;
 RECT 23.69 0.28 24.285 0.38 ;
 RECT 7.945 1.575 8.045 2.485 ;
 RECT 8.455 1.575 8.685 1.685 ;
 RECT 7.945 1.475 8.685 1.575 ;
 RECT 25.875 0.195 25.975 2.665 ;
 RECT 24.865 0.095 25.975 0.195 ;
 RECT 24.865 0.195 24.965 0.945 ;
 RECT 21.24 1.78 21.34 2.665 ;
 RECT 21.24 1.57 21.525 1.78 ;
 RECT 21.24 2.665 25.975 2.765 ;
 RECT 12.17 0.795 12.335 0.925 ;
 RECT 11.49 0.885 11.72 0.925 ;
 RECT 11.49 1.025 11.72 1.095 ;
 RECT 11.49 0.925 12.335 1.025 ;
 RECT 12.17 0.585 12.4 0.795 ;
 RECT 3.26 0.47 3.555 0.705 ;
 RECT 3.26 0.705 3.36 1.17 ;
 RECT 2.83 1.27 2.93 1.445 ;
 RECT 2.83 1.17 3.36 1.27 ;
 RECT 2.685 1.445 2.93 1.69 ;
 RECT 4.16 0.715 4.26 1.61 ;
 RECT 4.195 1.71 4.295 2.48 ;
 RECT 4.16 1.61 4.295 1.71 ;
 RECT 4.04 0.485 4.28 0.715 ;
 RECT 9.765 0.655 9.865 1.24 ;
 RECT 9.155 1.34 9.385 1.475 ;
 RECT 9.155 1.24 9.865 1.34 ;
 RECT 1.565 0.49 1.665 1.495 ;
 RECT 1.37 1.495 1.665 1.745 ;
 RECT 1.565 1.745 1.665 2.37 ;
 RECT 3.72 1.33 3.86 1.475 ;
 RECT 3.72 1.71 3.82 2.475 ;
 RECT 3.76 0.65 3.86 1.33 ;
 RECT 3.72 1.475 3.95 1.71 ;
 RECT 1.09 0.46 1.19 1.125 ;
 RECT 1.09 1.225 1.19 2.465 ;
 RECT 0.205 1.225 0.435 1.385 ;
 RECT 0.205 1.125 1.19 1.225 ;
 RECT 8.87 0.655 8.97 1.18 ;
 RECT 8.87 1.28 8.97 1.655 ;
 RECT 7.955 0.66 8.055 1.18 ;
 RECT 8.87 1.655 9.83 1.755 ;
 RECT 9.73 1.755 9.83 2.255 ;
 RECT 8.87 1.755 8.97 2.51 ;
 RECT 7.955 1.18 8.97 1.28 ;
 RECT 9.73 2.255 9.96 2.465 ;
 RECT 16.19 0.77 16.29 2.155 ;
 RECT 16.19 0.55 16.29 0.56 ;
 RECT 16.19 0.56 16.445 0.77 ;
 RECT 16.825 0.43 16.925 1.245 ;
 RECT 17.555 0.39 17.655 1.4 ;
 RECT 17.555 1.5 17.655 2.37 ;
 RECT 18.045 0.51 18.145 1.4 ;
 RECT 18.045 1.5 18.145 2.37 ;
 RECT 16.76 0.22 16.99 0.29 ;
 RECT 16.76 0.39 16.99 0.43 ;
 RECT 16.76 0.29 17.655 0.39 ;
 RECT 17.555 1.4 18.145 1.5 ;
 RECT 16.775 1.245 17.005 1.455 ;
 RECT 4.98 2.445 5.24 2.655 ;
 RECT 5.14 1.79 5.24 2.445 ;
 RECT 15.25 1.445 15.35 2.035 ;
 RECT 15.235 2.035 15.465 2.245 ;
 RECT 15.72 0.55 15.82 2.69 ;
 RECT 6.65 1.58 6.75 1.62 ;
 RECT 6.39 1.01 6.49 1.48 ;
 RECT 6.65 1.83 6.75 2.69 ;
 RECT 6.65 1.62 6.885 1.83 ;
 RECT 6.39 1.48 6.75 1.58 ;
 RECT 6.65 2.69 15.82 2.79 ;
 RECT 6.09 0.98 6.19 1.615 ;
 RECT 5.95 1.615 6.19 1.825 ;
 RECT 6.09 1.825 6.19 2.51 ;
 RECT 19.07 1.33 19.75 1.43 ;
 RECT 19.07 1.13 19.32 1.33 ;
 RECT 19.07 1.43 19.17 2.575 ;
 RECT 19.65 0.355 19.75 1.33 ;
 RECT 19.07 0.385 19.17 1.13 ;
 LAYER CO ;
 RECT 0.84 2.115 0.97 2.245 ;
 RECT 17.785 0.36 17.915 0.49 ;
 RECT 19.875 0.63 20.005 0.76 ;
 RECT 23.94 0.595 24.07 0.725 ;
 RECT 3.375 0.525 3.505 0.655 ;
 RECT 4.42 1.825 4.55 1.955 ;
 RECT 24.45 1.49 24.58 1.62 ;
 RECT 16.415 1.705 16.545 1.835 ;
 RECT 17.7 2.64 17.83 2.77 ;
 RECT 24.08 1.405 24.21 1.535 ;
 RECT 7.7 0.905 7.83 1.035 ;
 RECT 5.84 0.315 5.97 0.445 ;
 RECT 8.175 0.905 8.305 1.035 ;
 RECT 11.45 0.595 11.58 0.725 ;
 RECT 9.51 0.62 9.64 0.75 ;
 RECT 23.605 1.445 23.735 1.575 ;
 RECT 0.34 1.825 0.47 1.955 ;
 RECT 14.475 1.035 14.605 1.165 ;
 RECT 15.06 0.91 15.19 1.04 ;
 RECT 6.87 2.11 7 2.24 ;
 RECT 19.375 0.62 19.505 0.75 ;
 RECT 5.36 2.135 5.49 2.265 ;
 RECT 2.975 2.105 3.105 2.235 ;
 RECT 3.94 2.11 4.07 2.24 ;
 RECT 1.895 0.145 2.025 0.275 ;
 RECT 10.945 1.9 11.075 2.03 ;
 RECT 0.34 2.345 0.47 2.475 ;
 RECT 2.05 2.345 2.18 2.475 ;
 RECT 23 0.435 23.13 0.565 ;
 RECT 17.295 1.705 17.425 1.835 ;
 RECT 6.65 1.23 6.78 1.36 ;
 RECT 15.47 1.705 15.6 1.835 ;
 RECT 5.84 2.075 5.97 2.205 ;
 RECT 3.48 0.88 3.61 1.01 ;
 RECT 13.5 1.835 13.63 1.965 ;
 RECT 0.255 1.215 0.385 1.345 ;
 RECT 9.78 2.295 9.91 2.425 ;
 RECT 19.14 1.17 19.27 1.3 ;
 RECT 16.825 1.285 16.955 1.415 ;
 RECT 14.645 0.43 14.775 0.56 ;
 RECT 16.265 0.6 16.395 0.73 ;
 RECT 16.81 0.26 16.94 0.39 ;
 RECT 5.03 2.485 5.16 2.615 ;
 RECT 15.285 2.075 15.415 2.205 ;
 RECT 6.705 1.66 6.835 1.79 ;
 RECT 6 1.655 6.13 1.785 ;
 RECT 20.305 0.26 20.435 0.39 ;
 RECT 25.245 1.03 25.375 1.16 ;
 RECT 12.945 0.495 13.075 0.625 ;
 RECT 14.135 1.43 14.265 1.56 ;
 RECT 12.22 0.625 12.35 0.755 ;
 RECT 12.14 1.445 12.27 1.575 ;
 RECT 22.395 1.075 22.525 1.205 ;
 RECT 7.27 0.935 7.4 1.065 ;
 RECT 23.32 0.975 23.45 1.105 ;
 RECT 13.8 0.665 13.93 0.795 ;
 RECT 22.84 1.035 22.97 1.165 ;
 RECT 25.28 2.31 25.41 2.44 ;
 RECT 10.515 2.34 10.645 2.47 ;
 RECT 21.085 0.88 21.215 1.01 ;
 RECT 24.105 0.26 24.235 0.39 ;
 RECT 8.505 1.515 8.635 1.645 ;
 RECT 21.345 1.61 21.475 1.74 ;
 RECT 11.54 0.925 11.67 1.055 ;
 RECT 3.01 0.88 3.14 1.01 ;
 RECT 11.45 1.87 11.58 2 ;
 RECT 4.89 2.11 5.02 2.24 ;
 RECT 4.705 0.32 4.835 0.45 ;
 RECT 22.22 0.135 22.35 0.265 ;
 RECT 1.965 1.495 2.095 1.625 ;
 RECT 1.915 0.745 2.045 0.875 ;
 RECT 1.785 1.995 1.915 2.125 ;
 RECT 8.62 1.995 8.75 2.125 ;
 RECT 0.34 0.59 0.47 0.72 ;
 RECT 8.175 2.07 8.305 2.2 ;
 RECT 10.945 0.595 11.075 0.725 ;
 RECT 2.74 1.49 2.87 1.62 ;
 RECT 9.205 1.28 9.335 1.41 ;
 RECT 18.815 1.725 18.945 1.855 ;
 RECT 0.34 2.085 0.47 2.215 ;
 RECT 6.38 2.045 6.51 2.175 ;
 RECT 1.43 1.55 1.56 1.68 ;
 RECT 13.37 0.765 13.5 0.895 ;
 RECT 1.31 0.74 1.44 0.87 ;
 RECT 24.615 0.12 24.745 0.25 ;
 RECT 4.095 0.53 4.225 0.66 ;
 RECT 18.815 0.62 18.945 0.75 ;
 RECT 12.345 2.38 12.475 2.51 ;
 RECT 8.62 0.905 8.75 1.035 ;
 RECT 21.75 1.425 21.88 1.555 ;
 RECT 0.34 0.33 0.47 0.46 ;
 RECT 16.535 0.92 16.665 1.05 ;
 RECT 22.22 1.475 22.35 1.605 ;
 RECT 10.42 0.875 10.55 1.005 ;
 RECT 2.625 0.79 2.755 0.92 ;
 RECT 14.44 1.835 14.57 1.965 ;
 RECT 3.47 2.07 3.6 2.2 ;
 RECT 26.175 1.475 26.305 1.605 ;
 RECT 18.3 1.705 18.43 1.835 ;
 RECT 19.875 1.71 20.005 1.84 ;
 RECT 17.295 0.975 17.425 1.105 ;
 RECT 0.84 0.74 0.97 0.87 ;
 RECT 2.56 1.825 2.69 1.955 ;
 RECT 10.42 1.945 10.55 2.075 ;
 RECT 1.31 2.05 1.44 2.18 ;
 RECT 21.5 0.505 21.63 0.635 ;
 RECT 7.695 2.015 7.825 2.145 ;
 RECT 23.435 0.12 23.565 0.25 ;
 RECT 23 1.485 23.13 1.615 ;
 RECT 25.395 1.465 25.525 1.595 ;
 RECT 15.94 1.705 16.07 1.835 ;
 RECT 25.395 0.595 25.525 0.725 ;
 RECT 3.77 1.525 3.9 1.655 ;
 RECT 9.32 2.225 9.45 2.355 ;
 RECT 18.3 0.975 18.43 1.105 ;
 RECT 19.29 2.64 19.42 2.77 ;
 LAYER M1 ;
 RECT 25.195 1.18 25.425 1.2 ;
 RECT 24.055 0.29 24.425 0.43 ;
 RECT 24.285 0.43 24.425 0.71 ;
 RECT 24.055 0.22 24.285 0.29 ;
 RECT 25.705 0.85 25.845 1.385 ;
 RECT 25.39 1.525 25.53 1.73 ;
 RECT 24.285 0.71 25.845 0.85 ;
 RECT 25.39 0.51 25.53 0.71 ;
 RECT 25.39 1.385 25.845 1.525 ;
 RECT 21.435 1.195 21.885 1.225 ;
 RECT 21.745 1.225 21.885 1.61 ;
 RECT 21.57 0.64 21.71 1.015 ;
 RECT 21.295 1.57 21.525 1.61 ;
 RECT 21.295 1.75 21.525 1.78 ;
 RECT 21.435 1.015 21.745 1.055 ;
 RECT 21.285 1.61 21.885 1.75 ;
 RECT 21.45 0.5 21.71 0.64 ;
 RECT 22.345 1.035 22.575 1.055 ;
 RECT 22.345 1.195 22.575 1.245 ;
 RECT 21.435 1.055 22.575 1.195 ;
 RECT 23.315 1.145 23.455 1.345 ;
 RECT 22.995 1.485 23.135 1.76 ;
 RECT 23.315 0.73 23.455 0.935 ;
 RECT 22.995 0.355 23.135 0.59 ;
 RECT 22.995 1.345 23.455 1.485 ;
 RECT 23.27 0.935 23.5 1.145 ;
 RECT 22.995 0.59 23.455 0.73 ;
 RECT 20.255 0.36 20.485 0.43 ;
 RECT 21.85 0.36 21.99 0.565 ;
 RECT 20.255 0.22 21.99 0.36 ;
 RECT 22.59 0.705 22.73 0.75 ;
 RECT 22.715 0.995 23.02 1.205 ;
 RECT 22.715 0.89 22.855 0.995 ;
 RECT 22.59 0.75 22.855 0.89 ;
 RECT 21.85 0.565 22.73 0.705 ;
 RECT 15.49 0.775 15.63 1.405 ;
 RECT 16.215 0.56 16.445 0.635 ;
 RECT 14.47 1.405 15.63 1.545 ;
 RECT 14.47 1.545 14.61 1.83 ;
 RECT 13.425 1.83 14.675 1.97 ;
 RECT 14.47 1.17 14.61 1.405 ;
 RECT 14.4 1.03 14.68 1.17 ;
 RECT 18.41 0.36 18.55 0.635 ;
 RECT 15.49 0.635 18.55 0.775 ;
 RECT 19.09 0.36 19.23 1.13 ;
 RECT 19.09 1.13 19.32 1.34 ;
 RECT 18.41 0.22 19.23 0.36 ;
 RECT 14.595 0.28 16.99 0.42 ;
 RECT 14.595 0.42 14.825 0.6 ;
 RECT 16.76 0.22 16.99 0.28 ;
 RECT 16.76 0.42 16.99 0.43 ;
 RECT 11.445 0.525 11.585 0.885 ;
 RECT 11.445 1.095 11.585 2.065 ;
 RECT 11.445 0.885 11.72 1.095 ;
 RECT 8.965 2.055 9.105 2.34 ;
 RECT 8.17 2.34 9.105 2.48 ;
 RECT 9.485 1.66 9.625 1.915 ;
 RECT 8.965 1.915 9.625 2.055 ;
 RECT 8.17 1.04 8.31 2.34 ;
 RECT 8.17 0.895 8.31 0.9 ;
 RECT 8.1 0.9 8.375 1.04 ;
 RECT 9.485 1.52 11.08 1.66 ;
 RECT 10.94 0.525 11.08 1.52 ;
 RECT 10.94 1.66 11.08 2.11 ;
 RECT 10.415 0.765 10.555 1.52 ;
 RECT 10.415 1.66 10.555 2.145 ;
 RECT 13.75 0.57 13.98 0.95 ;
 RECT 12.17 0.585 13.125 0.63 ;
 RECT 12.17 0.63 12.4 0.795 ;
 RECT 12.195 0.49 13.125 0.585 ;
 RECT 12.895 0.455 13.125 0.49 ;
 RECT 12.895 0.63 13.125 0.665 ;
 RECT 3.755 0.66 3.895 0.92 ;
 RECT 3.3 0.52 3.895 0.66 ;
 RECT 3.755 0.92 7.45 1.06 ;
 RECT 7.22 0.895 7.45 0.92 ;
 RECT 7.22 1.06 7.45 1.105 ;
 RECT 1.865 0.88 2.005 1.475 ;
 RECT 1.825 1.63 1.965 1.99 ;
 RECT 1.825 1.475 2.17 1.63 ;
 RECT 1.715 1.99 1.965 2.13 ;
 RECT 1.865 0.74 2.185 0.88 ;
 RECT 3.31 1.82 4.89 1.96 ;
 RECT 4.75 1.79 4.89 1.82 ;
 RECT 3.395 1.96 3.675 2.215 ;
 RECT 3.475 0.805 3.615 1.22 ;
 RECT 3.31 1.22 3.615 1.36 ;
 RECT 3.31 1.36 3.45 1.82 ;
 RECT 5.95 1.615 6.18 1.65 ;
 RECT 5.95 1.79 6.18 1.825 ;
 RECT 4.75 1.65 6.185 1.79 ;
 RECT 0.615 0.875 0.755 1.195 ;
 RECT 0.615 1.335 0.755 2.11 ;
 RECT 0.615 2.25 0.755 2.255 ;
 RECT 0.615 2.11 1.04 2.25 ;
 RECT 0.615 0.735 1.04 0.875 ;
 RECT 1.585 0.6 1.725 1.195 ;
 RECT 0.615 1.195 1.725 1.335 ;
 RECT 3.005 0.97 3.155 1.085 ;
 RECT 3.015 1.085 3.155 2.035 ;
 RECT 3.005 0.36 3.145 0.97 ;
 RECT 2.33 0.22 3.145 0.36 ;
 RECT 2.33 0.36 2.47 0.46 ;
 RECT 2.97 2.17 3.11 2.305 ;
 RECT 2.97 2.035 3.155 2.17 ;
 RECT 1.585 0.46 2.47 0.6 ;
 RECT 2.62 1.67 2.76 1.82 ;
 RECT 2.62 1.96 2.76 2.51 ;
 RECT 2.62 0.5 2.76 1.44 ;
 RECT 2.62 1.44 2.875 1.67 ;
 RECT 2.49 1.82 2.76 1.96 ;
 RECT 4.98 2.445 5.21 2.51 ;
 RECT 4.98 2.65 5.21 2.655 ;
 RECT 2.62 2.51 5.21 2.65 ;
 RECT 12.86 1.895 13 2.39 ;
 RECT 17.005 2.205 17.145 2.39 ;
 RECT 12.86 2.39 17.145 2.53 ;
 RECT 11.735 1.755 13 1.895 ;
 RECT 11.735 1.895 11.875 2.34 ;
 RECT 10.465 2.3 10.695 2.34 ;
 RECT 10.465 2.48 10.695 2.51 ;
 RECT 10.465 2.34 11.875 2.48 ;
 RECT 20.89 2.205 21.03 2.52 ;
 RECT 17.005 2.065 21.03 2.205 ;
 RECT 25.23 2.48 25.37 2.52 ;
 RECT 20.89 2.52 25.37 2.66 ;
 RECT 25.23 2.27 25.46 2.48 ;
 RECT 16.3 1.7 16.595 1.84 ;
 RECT 16.3 1.84 16.44 2.075 ;
 RECT 15.605 1.84 15.745 2.075 ;
 RECT 15.41 1.7 15.745 1.84 ;
 RECT 15.605 2.075 16.44 2.215 ;
 RECT 16.495 1.055 16.635 1.245 ;
 RECT 15.935 1.385 16.075 1.625 ;
 RECT 16.775 1.385 17.005 1.455 ;
 RECT 15.935 1.245 17.005 1.385 ;
 RECT 16.465 0.915 16.765 1.055 ;
 RECT 15.905 1.625 16.16 1.92 ;
 RECT 13.14 1.56 13.28 2.11 ;
 RECT 12.09 1.405 12.32 1.42 ;
 RECT 12.09 1.56 12.32 1.615 ;
 RECT 12.09 1.42 13.28 1.56 ;
 RECT 13.14 2.11 15.465 2.245 ;
 RECT 13.14 2.245 15.46 2.25 ;
 RECT 15.235 2.035 15.465 2.11 ;
 RECT 8.615 1.775 8.755 2.18 ;
 RECT 8.615 1.04 8.755 1.475 ;
 RECT 8.455 1.475 8.755 1.635 ;
 RECT 8.545 0.9 8.82 1.04 ;
 RECT 8.615 1.685 9.34 1.775 ;
 RECT 8.455 1.635 9.34 1.685 ;
 RECT 9.2 1.21 9.34 1.635 ;
 RECT 3.87 2.105 5.09 2.245 ;
 RECT 4.43 1.225 7.08 1.25 ;
 RECT 6.375 1.365 6.515 2.25 ;
 RECT 4.43 1.365 4.57 1.5 ;
 RECT 3.6 1.64 4.105 1.675 ;
 RECT 3.6 1.5 4.57 1.64 ;
 RECT 7.69 1.04 7.83 1.25 ;
 RECT 7.69 1.39 7.83 2.215 ;
 RECT 7.69 0.885 7.83 0.9 ;
 RECT 4.43 1.25 7.83 1.365 ;
 RECT 6.94 1.365 7.83 1.39 ;
 RECT 7.625 0.9 7.9 1.04 ;
 RECT 23.935 0.73 24.075 1.04 ;
 RECT 24.075 1.18 24.215 1.605 ;
 RECT 23.87 0.59 24.145 0.73 ;
 RECT 25.195 0.99 25.425 1.04 ;
 RECT 23.935 1.04 25.425 1.18 ;
 END
END RDFFNSRASRX1

MACRO RDFFNSRASRX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 30.08 BY 2.88 ;
 PIN SAVE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 23.185 0.84 23.48 1.08 ;
 RECT 23.185 0.755 23.415 0.84 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SAVE

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 28.275 1.435 28.615 1.8 ;
 RECT 26.595 1.99 28.46 2.13 ;
 RECT 24.365 2.22 26.735 2.36 ;
 RECT 26.595 1.435 26.735 1.99 ;
 RECT 28.32 1.8 28.46 1.99 ;
 RECT 24.365 1.39 24.505 2.22 ;
 RECT 25.75 1.37 25.89 2.22 ;
 RECT 26.595 2.13 26.735 2.22 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.175 1.135 0.46 1.42 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.825 0.08 2.105 0.295 ;
 RECT 26.715 0.08 26.955 0.26 ;
 RECT 5.755 0.31 6.045 0.45 ;
 RECT 9.44 0.59 9.71 0.73 ;
 RECT 13.365 0.275 14.39 0.415 ;
 RECT 19.05 0.335 19.315 0.495 ;
 RECT 18.045 0.335 18.31 0.495 ;
 RECT 14.25 0.75 15.195 0.89 ;
 RECT 0 -0.08 30.08 0.08 ;
 RECT 1.305 0.08 1.445 0.97 ;
 RECT 0.335 0.08 0.475 0.775 ;
 RECT 4.65 0.08 4.885 0.46 ;
 RECT 20.565 0.08 20.705 0.82 ;
 RECT 21.63 0.08 21.77 0.82 ;
 RECT 24.365 0.08 24.505 0.36 ;
 RECT 25.58 0.08 25.72 0.35 ;
 RECT 5.835 0.08 5.975 0.31 ;
 RECT 9.505 0.08 9.645 0.59 ;
 RECT 13.365 0.415 13.505 0.945 ;
 RECT 13.365 0.08 13.505 0.275 ;
 RECT 19.105 0.08 19.245 0.335 ;
 RECT 18.1 0.08 18.24 0.335 ;
 RECT 15.055 0.89 15.195 1.11 ;
 RECT 14.25 0.415 14.39 0.75 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 9.245 2.215 9.475 2.355 ;
 RECT 0 2.8 30.08 2.96 ;
 RECT 1.98 2.34 2.23 2.8 ;
 RECT 0.335 1.74 0.475 2.8 ;
 RECT 1.305 1.98 1.445 2.8 ;
 RECT 6.865 2 7.005 2.8 ;
 RECT 5.835 1.98 5.975 2.8 ;
 RECT 5.355 2.07 5.495 2.8 ;
 RECT 12.275 2.335 12.545 2.8 ;
 RECT 20.48 2.57 20.62 2.8 ;
 RECT 19.02 2.57 19.16 2.8 ;
 RECT 18.015 2.57 18.155 2.8 ;
 RECT 21.545 2.57 21.685 2.8 ;
 RECT 9.29 2.355 9.43 2.8 ;
 RECT 9.29 2.195 9.43 2.215 ;
 END
 END VDD

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.355 1.475 1.725 1.775 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN NRESTORE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.78 2.26 10.36 2.47 ;
 RECT 10.115 2.12 10.36 2.26 ;
 END
 ANTENNAGATEAREA 0.126 ;
 END NRESTORE

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.04 0.745 4.36 0.76 ;
 RECT 4.04 0.485 4.36 0.605 ;
 RECT 8.965 0.89 10.02 1.03 ;
 RECT 9.875 0.245 12.025 0.255 ;
 RECT 9.875 0.255 12.03 0.385 ;
 RECT 11.89 1.09 13.88 1.23 ;
 RECT 14.085 1.56 14.315 1.6 ;
 RECT 13.74 1.42 14.315 1.56 ;
 RECT 14.085 1.39 14.315 1.42 ;
 RECT 4.04 0.605 9.105 0.745 ;
 RECT 8.965 0.745 9.105 0.89 ;
 RECT 9.88 0.385 10.02 0.89 ;
 RECT 11.89 0.385 12.03 1.09 ;
 RECT 13.74 1.23 13.88 1.42 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END RSTB

 PIN SETB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.23 1.795 7.49 2.055 ;
 RECT 6.655 1.795 6.885 1.83 ;
 RECT 6.655 1.655 7.49 1.795 ;
 RECT 6.655 1.62 6.885 1.655 ;
 END
 ANTENNAGATEAREA 0.114 ;
 END SETB

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.405 1.155 17.76 1.445 ;
 RECT 17.61 0.915 17.75 1.155 ;
 RECT 18.615 1.84 18.755 1.885 ;
 RECT 18.615 0.915 18.755 1.7 ;
 RECT 19.59 1.84 19.73 1.885 ;
 RECT 19.59 0.915 19.73 1.7 ;
 RECT 17.61 1.7 19.73 1.84 ;
 RECT 17.61 1.84 17.75 1.885 ;
 RECT 17.61 1.445 17.75 1.7 ;
 END
 ANTENNADIFFAREA 1.145 ;
 END QN

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 20.005 0.51 20.145 1.48 ;
 RECT 21.065 1.905 21.205 1.91 ;
 RECT 21.065 0.56 21.205 1.765 ;
 RECT 22.13 1.905 22.27 1.91 ;
 RECT 22.13 0.56 22.27 1.765 ;
 RECT 20.005 1.905 20.145 1.915 ;
 RECT 20.005 1.48 20.28 1.765 ;
 RECT 20.005 1.765 22.27 1.905 ;
 END
 ANTENNADIFFAREA 0.909 ;
 END Q

 OBS
 LAYER PO ;
 RECT 22.405 0.22 22.635 0.275 ;
 RECT 22.405 0.375 22.635 0.43 ;
 RECT 21.91 0.275 22.635 0.375 ;
 RECT 14.22 0.73 14.32 1.39 ;
 RECT 14.085 1.39 14.32 1.6 ;
 RECT 14.22 1.6 14.32 2.39 ;
 RECT 2.405 0.285 2.505 1.52 ;
 RECT 1.905 1.52 2.505 1.62 ;
 RECT 2.405 0.185 11.295 0.195 ;
 RECT 4.46 0.095 11.295 0.185 ;
 RECT 2.405 0.195 4.56 0.285 ;
 RECT 11.195 0.195 11.295 1.29 ;
 RECT 12.09 1.39 12.285 1.405 ;
 RECT 3.225 1.565 3.325 2.675 ;
 RECT 2.34 1.62 2.44 2.675 ;
 RECT 1.905 1.44 2.15 1.52 ;
 RECT 1.905 1.62 2.15 1.69 ;
 RECT 4.46 0.285 4.56 1.24 ;
 RECT 11.195 1.29 12.285 1.39 ;
 RECT 2.34 2.675 3.325 2.775 ;
 RECT 12.09 1.405 12.32 1.615 ;
 RECT 24.625 1.245 24.725 2.02 ;
 RECT 24.495 1.035 24.725 1.245 ;
 RECT 12.585 0.105 15.41 0.205 ;
 RECT 12.585 0.205 12.685 1.91 ;
 RECT 15.31 0.205 15.41 1.265 ;
 RECT 11.765 1.71 11.865 1.91 ;
 RECT 10.68 1.61 11.865 1.71 ;
 RECT 10.68 0.475 10.78 1.61 ;
 RECT 11.23 1.71 11.33 2.425 ;
 RECT 7.345 0.475 7.445 0.895 ;
 RECT 11.765 1.91 12.685 2.01 ;
 RECT 7.345 0.375 10.78 0.475 ;
 RECT 7.22 0.895 7.45 1.105 ;
 RECT 12.895 0.455 14.825 0.535 ;
 RECT 14.595 0.535 14.825 0.6 ;
 RECT 14.595 0.39 14.825 0.435 ;
 RECT 12.975 0.435 14.825 0.455 ;
 RECT 12.895 0.535 13.125 0.665 ;
 RECT 13.75 0.535 13.98 0.835 ;
 RECT 13.75 0.835 13.85 2.39 ;
 RECT 24.93 0.215 25.03 0.995 ;
 RECT 24.93 0.995 25.17 1.205 ;
 RECT 24.93 1.205 25.03 2 ;
 RECT 27.325 0.375 27.425 0.99 ;
 RECT 27.325 0.99 27.575 1.2 ;
 RECT 27.325 1.2 27.425 2.27 ;
 RECT 27.325 2.27 27.61 2.48 ;
 RECT 10.195 0.655 10.295 2.305 ;
 RECT 10.58 2.3 10.81 2.305 ;
 RECT 10.58 2.405 10.81 2.51 ;
 RECT 10.195 2.305 10.815 2.405 ;
 RECT 24.15 0.21 24.25 0.755 ;
 RECT 24.15 0.855 24.25 2.2 ;
 RECT 27.015 1.125 27.115 2.2 ;
 RECT 23.185 0.755 24.72 0.84 ;
 RECT 23.185 0.84 24.715 0.855 ;
 RECT 24.62 0.215 24.72 0.755 ;
 RECT 23.185 0.855 23.415 0.965 ;
 RECT 24.15 2.2 27.115 2.3 ;
 RECT 25.84 1.06 25.94 1.14 ;
 RECT 25.84 0.38 25.94 0.96 ;
 RECT 25.84 1.14 26.11 1.24 ;
 RECT 26.01 1.24 26.11 1.84 ;
 RECT 25.42 0.935 25.65 0.96 ;
 RECT 25.42 0.96 25.94 1.06 ;
 RECT 25.42 1.06 25.65 1.145 ;
 RECT 26.205 0.22 26.435 0.28 ;
 RECT 26.205 0.38 26.435 0.43 ;
 RECT 25.84 0.28 26.435 0.38 ;
 RECT 7.945 1.575 8.045 2.485 ;
 RECT 8.455 1.575 8.685 1.685 ;
 RECT 7.945 1.475 8.685 1.575 ;
 RECT 28.025 0.195 28.125 2.665 ;
 RECT 27.015 0.095 28.125 0.195 ;
 RECT 27.015 0.195 27.115 0.945 ;
 RECT 23.39 1.665 23.49 2.665 ;
 RECT 23.39 1.45 23.49 1.455 ;
 RECT 23.39 1.455 23.675 1.665 ;
 RECT 23.39 2.665 28.125 2.765 ;
 RECT 12.17 0.795 12.335 0.925 ;
 RECT 11.49 0.885 11.72 0.925 ;
 RECT 11.49 1.025 11.72 1.095 ;
 RECT 11.49 0.925 12.335 1.025 ;
 RECT 12.17 0.585 12.4 0.795 ;
 RECT 1.565 0.49 1.665 1.495 ;
 RECT 1.37 1.495 1.665 1.745 ;
 RECT 1.565 1.745 1.665 2.37 ;
 RECT 3.72 1.33 3.86 1.475 ;
 RECT 3.72 1.71 3.82 2.475 ;
 RECT 3.76 0.65 3.86 1.33 ;
 RECT 3.72 1.475 3.95 1.71 ;
 RECT 4.16 0.715 4.26 1.61 ;
 RECT 4.195 1.71 4.295 2.48 ;
 RECT 4.16 1.61 4.295 1.71 ;
 RECT 4.04 0.485 4.28 0.715 ;
 RECT 3.26 0.705 3.36 1.165 ;
 RECT 2.83 1.27 2.93 1.445 ;
 RECT 3.26 0.47 3.555 0.705 ;
 RECT 2.83 1.17 3.37 1.265 ;
 RECT 3.06 1.165 3.37 1.17 ;
 RECT 2.83 1.265 3.205 1.27 ;
 RECT 2.685 1.445 2.93 1.69 ;
 RECT 1.09 0.27 1.19 1.165 ;
 RECT 1.09 1.265 1.19 2.465 ;
 RECT 0.205 1.265 0.435 1.39 ;
 RECT 0.205 1.165 1.19 1.265 ;
 RECT 9.765 0.655 9.865 1.155 ;
 RECT 9.15 1.255 9.38 1.405 ;
 RECT 9.15 1.155 9.865 1.255 ;
 RECT 8.87 0.655 8.97 1.18 ;
 RECT 8.87 1.28 8.97 1.655 ;
 RECT 7.955 0.66 8.055 1.18 ;
 RECT 9.88 1.445 9.98 1.655 ;
 RECT 9.88 1.755 9.98 2.26 ;
 RECT 8.87 1.755 8.97 2.51 ;
 RECT 7.955 1.18 8.97 1.28 ;
 RECT 8.87 1.655 9.98 1.755 ;
 RECT 9.78 2.26 10.01 2.47 ;
 RECT 16.19 0.77 16.29 2.155 ;
 RECT 16.19 0.55 16.29 0.56 ;
 RECT 16.19 0.56 16.445 0.77 ;
 RECT 17.875 0.39 17.975 1.4 ;
 RECT 17.875 1.5 17.975 2.37 ;
 RECT 16.825 0.43 16.925 1.245 ;
 RECT 16.76 0.3 17.975 0.39 ;
 RECT 16.76 0.29 17.96 0.3 ;
 RECT 19.37 0.51 19.47 1.4 ;
 RECT 19.37 1.5 19.47 2.37 ;
 RECT 18.88 0.515 18.98 1.4 ;
 RECT 18.88 1.5 18.98 2.37 ;
 RECT 17.875 1.4 19.47 1.5 ;
 RECT 18.365 0.51 18.465 1.4 ;
 RECT 18.365 1.5 18.465 2.37 ;
 RECT 16.76 0.22 16.99 0.29 ;
 RECT 16.76 0.39 16.99 0.43 ;
 RECT 16.775 1.245 17.005 1.455 ;
 RECT 4.98 2.445 5.24 2.655 ;
 RECT 5.14 1.79 5.24 2.445 ;
 RECT 15.25 1.445 15.35 2.035 ;
 RECT 15.235 2.035 15.465 2.245 ;
 RECT 15.72 0.55 15.82 2.69 ;
 RECT 6.65 1.83 6.75 2.69 ;
 RECT 6.65 1.58 6.75 1.62 ;
 RECT 6.39 1.01 6.49 1.48 ;
 RECT 6.65 1.62 6.885 1.83 ;
 RECT 6.65 2.69 15.82 2.79 ;
 RECT 6.39 1.48 6.75 1.58 ;
 RECT 6.09 0.98 6.19 1.615 ;
 RECT 5.95 1.615 6.19 1.825 ;
 RECT 6.09 1.825 6.19 2.51 ;
 RECT 20.265 1.33 22.01 1.43 ;
 RECT 20.265 1.43 20.365 2.575 ;
 RECT 20.265 1.13 20.54 1.33 ;
 RECT 20.845 1.43 20.945 2.575 ;
 RECT 21.33 1.43 21.43 2.575 ;
 RECT 21.91 0.375 22.01 1.33 ;
 RECT 20.265 0.385 20.365 1.13 ;
 RECT 20.845 0.385 20.945 1.33 ;
 RECT 21.33 0.385 21.43 1.33 ;
 RECT 21.91 1.43 22.01 2.575 ;
 LAYER CO ;
 RECT 4.42 1.825 4.55 1.955 ;
 RECT 10.42 1.805 10.55 1.935 ;
 RECT 26.6 1.49 26.73 1.62 ;
 RECT 7.695 2.015 7.825 2.145 ;
 RECT 4.705 0.32 4.835 0.45 ;
 RECT 26.09 0.595 26.22 0.725 ;
 RECT 27.545 0.595 27.675 0.725 ;
 RECT 10.945 0.595 11.075 0.725 ;
 RECT 1.785 1.995 1.915 2.125 ;
 RECT 1.31 2.05 1.44 2.18 ;
 RECT 3.01 0.88 3.14 1.01 ;
 RECT 24.37 0.135 24.5 0.265 ;
 RECT 3.77 1.525 3.9 1.655 ;
 RECT 2.74 1.49 2.87 1.62 ;
 RECT 11.45 1.87 11.58 2 ;
 RECT 0.34 0.59 0.47 0.72 ;
 RECT 3.375 0.525 3.505 0.655 ;
 RECT 8.62 1.995 8.75 2.125 ;
 RECT 4.89 2.11 5.02 2.24 ;
 RECT 8.175 2.07 8.305 2.2 ;
 RECT 1.965 1.495 2.095 1.625 ;
 RECT 20.36 1.17 20.49 1.3 ;
 RECT 0.255 1.22 0.385 1.35 ;
 RECT 9.2 1.235 9.33 1.365 ;
 RECT 9.83 2.3 9.96 2.43 ;
 RECT 16.825 1.285 16.955 1.415 ;
 RECT 14.645 0.43 14.775 0.56 ;
 RECT 16.265 0.6 16.395 0.73 ;
 RECT 16.81 0.26 16.94 0.39 ;
 RECT 5.03 2.485 5.16 2.615 ;
 RECT 15.285 2.075 15.415 2.205 ;
 RECT 6.705 1.66 6.835 1.79 ;
 RECT 6 1.655 6.13 1.785 ;
 RECT 22.455 0.26 22.585 0.39 ;
 RECT 27.395 1.03 27.525 1.16 ;
 RECT 12.945 0.495 13.075 0.625 ;
 RECT 14.135 1.43 14.265 1.56 ;
 RECT 12.22 0.625 12.35 0.755 ;
 RECT 12.14 1.445 12.27 1.575 ;
 RECT 24.545 1.075 24.675 1.205 ;
 RECT 7.27 0.935 7.4 1.065 ;
 RECT 25.47 0.975 25.6 1.105 ;
 RECT 13.8 0.665 13.93 0.795 ;
 RECT 24.99 1.035 25.12 1.165 ;
 RECT 27.43 2.31 27.56 2.44 ;
 RECT 10.63 2.34 10.76 2.47 ;
 RECT 23.235 0.795 23.365 0.925 ;
 RECT 26.255 0.26 26.385 0.39 ;
 RECT 8.505 1.515 8.635 1.645 ;
 RECT 23.495 1.495 23.625 1.625 ;
 RECT 11.54 0.925 11.67 1.055 ;
 RECT 12.345 2.38 12.475 2.51 ;
 RECT 10.945 1.9 11.075 2.03 ;
 RECT 16.415 1.705 16.545 1.835 ;
 RECT 15.06 0.91 15.19 1.04 ;
 RECT 26.23 1.405 26.36 1.535 ;
 RECT 15.47 1.705 15.6 1.835 ;
 RECT 8.175 0.905 8.305 1.035 ;
 RECT 3.94 2.11 4.07 2.24 ;
 RECT 9.51 0.595 9.64 0.725 ;
 RECT 0.34 2.345 0.47 2.475 ;
 RECT 0.34 1.825 0.47 1.955 ;
 RECT 13.5 1.835 13.63 1.965 ;
 RECT 2.05 2.345 2.18 2.475 ;
 RECT 6.65 1.23 6.78 1.36 ;
 RECT 0.34 0.33 0.47 0.46 ;
 RECT 1.31 0.74 1.44 0.87 ;
 RECT 5.84 2.075 5.97 2.205 ;
 RECT 2.625 0.79 2.755 0.92 ;
 RECT 28.325 1.475 28.455 1.605 ;
 RECT 18.105 0.36 18.235 0.49 ;
 RECT 21.55 2.64 21.68 2.77 ;
 RECT 20.57 0.62 20.7 0.75 ;
 RECT 19.595 0.975 19.725 1.105 ;
 RECT 18.62 1.705 18.75 1.835 ;
 RECT 18.02 2.64 18.15 2.77 ;
 RECT 20.01 1.725 20.14 1.855 ;
 RECT 21.635 0.62 21.765 0.75 ;
 RECT 19.11 0.36 19.24 0.49 ;
 RECT 18.62 0.975 18.75 1.105 ;
 RECT 21.07 0.63 21.2 0.76 ;
 RECT 22.135 0.63 22.265 0.76 ;
 RECT 21.07 1.71 21.2 1.84 ;
 RECT 17.615 0.975 17.745 1.105 ;
 RECT 19.025 2.64 19.155 2.77 ;
 RECT 20.485 2.64 20.615 2.77 ;
 RECT 17.615 1.705 17.745 1.835 ;
 RECT 22.135 1.71 22.265 1.84 ;
 RECT 19.595 1.705 19.725 1.835 ;
 RECT 20.01 0.62 20.14 0.75 ;
 RECT 1.915 0.745 2.045 0.875 ;
 RECT 0.34 2.085 0.47 2.215 ;
 RECT 6.38 2.045 6.51 2.175 ;
 RECT 1.43 1.55 1.56 1.68 ;
 RECT 14.475 1.035 14.605 1.165 ;
 RECT 7.7 0.905 7.83 1.035 ;
 RECT 11.45 0.595 11.58 0.725 ;
 RECT 25.755 1.445 25.885 1.575 ;
 RECT 6.87 2.11 7 2.24 ;
 RECT 5.84 0.315 5.97 0.445 ;
 RECT 2.975 2.105 3.105 2.235 ;
 RECT 3.48 0.88 3.61 1.01 ;
 RECT 16.535 0.92 16.665 1.05 ;
 RECT 5.36 2.135 5.49 2.265 ;
 RECT 26.765 0.12 26.895 0.25 ;
 RECT 1.895 0.145 2.025 0.275 ;
 RECT 25.15 0.435 25.28 0.565 ;
 RECT 8.62 0.905 8.75 1.035 ;
 RECT 0.84 0.74 0.97 0.87 ;
 RECT 4.095 0.53 4.225 0.66 ;
 RECT 25.585 0.12 25.715 0.25 ;
 RECT 2.56 1.825 2.69 1.955 ;
 RECT 9.295 2.225 9.425 2.355 ;
 RECT 0.84 2.115 0.97 2.245 ;
 RECT 24.37 1.475 24.5 1.605 ;
 RECT 14.44 1.835 14.57 1.965 ;
 RECT 27.545 1.465 27.675 1.595 ;
 RECT 23.9 1.425 24.03 1.555 ;
 RECT 13.37 0.765 13.5 0.895 ;
 RECT 23.65 0.505 23.78 0.635 ;
 RECT 10.42 0.875 10.55 1.005 ;
 RECT 25.15 1.485 25.28 1.615 ;
 RECT 3.47 2.07 3.6 2.2 ;
 RECT 15.94 1.705 16.07 1.835 ;
 LAYER M1 ;
 RECT 26.085 1.04 27.575 1.18 ;
 RECT 27.345 1.18 27.575 1.2 ;
 RECT 26.205 0.29 26.575 0.43 ;
 RECT 26.435 0.43 26.575 0.71 ;
 RECT 26.205 0.22 26.435 0.29 ;
 RECT 27.855 0.85 27.995 1.385 ;
 RECT 27.54 1.525 27.68 1.73 ;
 RECT 26.435 0.71 27.995 0.85 ;
 RECT 27.54 0.51 27.68 0.71 ;
 RECT 27.54 1.385 27.995 1.525 ;
 RECT 23.895 1.195 24.035 1.455 ;
 RECT 23.72 0.64 23.86 1.055 ;
 RECT 23.445 1.595 23.675 1.665 ;
 RECT 23.895 1.595 24.035 1.665 ;
 RECT 23.445 1.455 24.035 1.595 ;
 RECT 23.6 0.5 23.86 0.64 ;
 RECT 24.495 1.035 24.725 1.055 ;
 RECT 23.72 1.055 24.725 1.195 ;
 RECT 24.495 1.195 24.725 1.245 ;
 RECT 25.465 1.145 25.605 1.345 ;
 RECT 25.145 1.485 25.285 1.76 ;
 RECT 25.465 0.73 25.605 0.935 ;
 RECT 25.145 0.355 25.285 0.59 ;
 RECT 25.145 1.345 25.605 1.485 ;
 RECT 25.42 0.935 25.65 1.145 ;
 RECT 25.145 0.59 25.605 0.73 ;
 RECT 22.405 0.36 22.635 0.43 ;
 RECT 24 0.36 24.14 0.565 ;
 RECT 22.405 0.22 24.14 0.36 ;
 RECT 24.74 0.705 24.88 0.75 ;
 RECT 24.865 0.995 25.17 1.205 ;
 RECT 24.865 0.89 25.005 0.995 ;
 RECT 24.74 0.75 25.005 0.89 ;
 RECT 24 0.565 24.88 0.705 ;
 RECT 13.75 0.57 13.98 0.95 ;
 RECT 16.76 0.22 16.99 0.28 ;
 RECT 16.76 0.42 16.99 0.43 ;
 RECT 14.595 0.28 16.99 0.42 ;
 RECT 14.595 0.42 14.825 0.6 ;
 RECT 15.49 0.775 15.63 1.405 ;
 RECT 16.215 0.56 16.445 0.635 ;
 RECT 14.47 1.405 15.63 1.545 ;
 RECT 14.47 1.545 14.61 1.83 ;
 RECT 13.425 1.83 14.675 1.97 ;
 RECT 14.47 1.17 14.61 1.405 ;
 RECT 14.4 1.03 14.68 1.17 ;
 RECT 19.605 0.36 19.745 0.635 ;
 RECT 15.49 0.635 19.745 0.775 ;
 RECT 20.285 1.13 20.54 1.34 ;
 RECT 20.285 0.36 20.425 1.13 ;
 RECT 19.605 0.22 20.425 0.36 ;
 RECT 12.17 0.585 13.125 0.63 ;
 RECT 12.895 0.63 13.125 0.665 ;
 RECT 12.895 0.455 13.125 0.49 ;
 RECT 12.195 0.49 13.125 0.585 ;
 RECT 12.17 0.63 12.4 0.795 ;
 RECT 11.445 0.525 11.585 0.885 ;
 RECT 11.445 1.095 11.585 2.065 ;
 RECT 11.445 0.885 11.72 1.095 ;
 RECT 8.965 2.055 9.105 2.34 ;
 RECT 8.17 2.34 9.105 2.48 ;
 RECT 9.525 1.6 9.665 1.915 ;
 RECT 8.965 1.915 9.665 2.055 ;
 RECT 8.17 1.04 8.31 2.34 ;
 RECT 8.17 0.895 8.31 0.9 ;
 RECT 8.1 0.9 8.375 1.04 ;
 RECT 10.415 0.765 10.555 1.46 ;
 RECT 10.415 1.6 10.555 1.8 ;
 RECT 10.94 0.525 11.08 1.46 ;
 RECT 10.94 1.6 11.08 2.11 ;
 RECT 9.525 1.46 11.08 1.6 ;
 RECT 10.35 1.8 10.62 1.94 ;
 RECT 3.755 0.66 3.895 0.905 ;
 RECT 3.3 0.52 3.895 0.66 ;
 RECT 3.755 0.905 7.455 1.045 ;
 RECT 7.22 0.895 7.45 0.905 ;
 RECT 7.22 1.045 7.45 1.105 ;
 RECT 3.31 1.82 4.89 1.96 ;
 RECT 4.75 1.79 4.89 1.82 ;
 RECT 3.395 1.96 3.675 2.215 ;
 RECT 3.475 0.805 3.615 1.22 ;
 RECT 3.31 1.22 3.615 1.36 ;
 RECT 3.31 1.36 3.45 1.82 ;
 RECT 5.95 1.615 6.18 1.65 ;
 RECT 5.95 1.79 6.18 1.825 ;
 RECT 4.75 1.65 6.185 1.79 ;
 RECT 0.615 1.335 0.755 2.11 ;
 RECT 0.615 2.25 0.755 2.255 ;
 RECT 0.615 0.875 0.755 1.195 ;
 RECT 0.615 2.11 1.04 2.25 ;
 RECT 0.615 0.735 1.04 0.875 ;
 RECT 0.615 1.195 1.725 1.335 ;
 RECT 1.585 0.6 1.725 1.195 ;
 RECT 3.005 0.97 3.155 1.08 ;
 RECT 3.015 1.08 3.155 2.035 ;
 RECT 3.005 0.36 3.145 0.97 ;
 RECT 2.33 0.22 3.145 0.36 ;
 RECT 2.33 0.36 2.47 0.46 ;
 RECT 2.97 2.17 3.11 2.305 ;
 RECT 2.97 2.035 3.155 2.17 ;
 RECT 1.585 0.46 2.47 0.6 ;
 RECT 1.865 0.88 2.005 1.475 ;
 RECT 1.715 1.99 2.005 2.13 ;
 RECT 1.865 1.63 2.005 1.99 ;
 RECT 1.865 1.475 2.17 1.63 ;
 RECT 1.865 0.74 2.185 0.88 ;
 RECT 2.62 1.67 2.76 1.82 ;
 RECT 2.62 1.96 2.76 2.51 ;
 RECT 2.62 0.5 2.76 1.44 ;
 RECT 2.62 1.44 2.875 1.67 ;
 RECT 2.49 1.82 2.76 1.96 ;
 RECT 4.98 2.445 5.21 2.51 ;
 RECT 4.98 2.65 5.21 2.655 ;
 RECT 2.62 2.51 5.21 2.65 ;
 RECT 12.86 1.895 13 2.39 ;
 RECT 17.005 2.205 17.145 2.39 ;
 RECT 12.86 2.39 17.145 2.53 ;
 RECT 11.735 1.755 13 1.895 ;
 RECT 11.735 1.895 11.875 2.34 ;
 RECT 10.58 2.3 10.81 2.34 ;
 RECT 10.58 2.34 11.875 2.48 ;
 RECT 10.58 2.48 10.81 2.51 ;
 RECT 17.005 2.065 23.18 2.205 ;
 RECT 23.04 2.205 23.18 2.52 ;
 RECT 27.38 2.48 27.52 2.52 ;
 RECT 23.04 2.52 27.52 2.66 ;
 RECT 27.38 2.27 27.61 2.48 ;
 RECT 15.41 1.7 15.745 1.84 ;
 RECT 15.605 1.84 15.745 2.075 ;
 RECT 16.3 1.84 16.44 2.075 ;
 RECT 16.3 1.7 16.595 1.84 ;
 RECT 15.605 2.075 16.44 2.215 ;
 RECT 16.495 1.055 16.635 1.245 ;
 RECT 15.935 1.385 16.075 1.625 ;
 RECT 15.935 1.245 17.005 1.385 ;
 RECT 16.775 1.385 17.005 1.455 ;
 RECT 16.465 0.915 16.765 1.055 ;
 RECT 15.905 1.625 16.16 1.92 ;
 RECT 13.14 1.56 13.28 2.11 ;
 RECT 12.09 1.405 12.32 1.42 ;
 RECT 12.09 1.42 13.28 1.56 ;
 RECT 12.09 1.56 12.32 1.615 ;
 RECT 13.14 2.11 15.465 2.245 ;
 RECT 15.235 2.035 15.465 2.11 ;
 RECT 13.14 2.245 15.46 2.25 ;
 RECT 8.615 1.775 8.755 2.18 ;
 RECT 8.615 1.04 8.755 1.475 ;
 RECT 8.455 1.475 8.755 1.635 ;
 RECT 8.545 0.9 8.82 1.04 ;
 RECT 9.065 1.41 9.205 1.635 ;
 RECT 8.615 1.685 9.205 1.775 ;
 RECT 8.455 1.635 9.205 1.685 ;
 RECT 9.065 1.195 9.38 1.41 ;
 RECT 3.87 2.105 5.09 2.245 ;
 RECT 4.43 1.225 7.08 1.25 ;
 RECT 6.375 1.365 6.515 2.25 ;
 RECT 4.43 1.365 4.57 1.5 ;
 RECT 3.6 1.64 4.105 1.675 ;
 RECT 3.6 1.5 4.57 1.64 ;
 RECT 7.69 1.04 7.83 1.25 ;
 RECT 7.69 1.39 7.83 2.215 ;
 RECT 7.69 0.885 7.83 0.9 ;
 RECT 4.43 1.25 7.83 1.365 ;
 RECT 6.94 1.365 7.83 1.39 ;
 RECT 7.625 0.9 7.9 1.04 ;
 RECT 26.085 0.73 26.225 1.04 ;
 RECT 26.225 1.18 26.365 1.605 ;
 RECT 26.02 0.59 26.295 0.73 ;
 RECT 27.345 0.99 27.575 1.04 ;
 END
END RDFFNSRASRX2

MACRO AND2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.77 0.84 1.1 1.08 ;
 END
 ANTENNAGATEAREA 0.062 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.26 1.945 1.535 2.365 ;
 END
 ANTENNAGATEAREA 0.062 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.185 1.105 2.425 1.345 ;
 RECT 2.185 1.345 2.325 2.565 ;
 RECT 2.185 0.275 2.325 1.105 ;
 END
 ANTENNADIFFAREA 0.464 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 0.77 1.495 0.91 2.8 ;
 RECT 1.71 1.495 1.85 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 RECT 1.71 0.08 1.85 0.555 ;
 RECT 0.31 0.08 0.45 0.755 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 1.81 1.12 2.065 1.35 ;
 RECT 1.965 0.105 2.065 1.12 ;
 RECT 1.965 1.35 2.065 2.75 ;
 RECT 1.025 0.105 1.125 0.845 ;
 RECT 1.025 1.075 1.125 2.03 ;
 RECT 0.895 0.845 1.125 1.075 ;
 RECT 1.495 0.105 1.595 1.925 ;
 RECT 1.305 1.925 1.595 2.155 ;
 LAYER CO ;
 RECT 2.19 2.33 2.32 2.46 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 1.355 1.98 1.485 2.11 ;
 RECT 0.945 0.895 1.075 1.025 ;
 RECT 1.86 1.17 1.99 1.3 ;
 RECT 2.19 0.325 2.32 0.455 ;
 RECT 1.715 0.325 1.845 0.455 ;
 RECT 0.775 0.325 0.905 0.455 ;
 RECT 1.715 1.545 1.845 1.675 ;
 RECT 2.19 2.065 2.32 2.195 ;
 RECT 2.19 1.805 2.32 1.935 ;
 RECT 2.19 1.545 2.32 1.675 ;
 RECT 1.715 1.545 1.845 1.675 ;
 RECT 1.245 1.545 1.375 1.675 ;
 RECT 0.775 1.545 0.905 1.675 ;
 LAYER M1 ;
 RECT 1.24 1.5 1.38 1.725 ;
 RECT 1.24 0.32 1.38 1.5 ;
 RECT 0.725 0.32 1.38 0.46 ;
 RECT 1.81 1.12 2.04 1.35 ;
 RECT 1.24 1.21 2.035 1.35 ;
 END
END AND2X1

MACRO AND2X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.88 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.115 0.96 1.45 ;
 END
 ANTENNAGATEAREA 0.062 ;
 END IN1

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.045 0.84 2.38 1.215 ;
 RECT 2.045 1.215 2.185 2.565 ;
 RECT 2.045 0.475 2.185 0.84 ;
 END
 ANTENNADIFFAREA 0.578 ;
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.88 0.08 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 1.57 0.08 1.71 0.825 ;
 RECT 2.52 0.08 2.66 0.775 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 1.945 1.395 2.365 ;
 END
 ANTENNAGATEAREA 0.062 ;
 END IN2

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.88 2.96 ;
 RECT 0.205 1.495 0.345 2.8 ;
 RECT 1.57 1.495 1.71 2.8 ;
 RECT 0.63 1.595 0.77 2.8 ;
 RECT 2.53 1.495 2.67 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.885 0.565 0.985 1.12 ;
 RECT 0.885 1.35 0.985 2.055 ;
 RECT 0.755 1.12 0.985 1.35 ;
 RECT 1.635 1.19 2.405 1.29 ;
 RECT 2.305 0.375 2.405 1.19 ;
 RECT 1.825 0.375 1.925 1.12 ;
 RECT 1.635 1.12 1.925 1.19 ;
 RECT 1.635 1.29 1.925 1.35 ;
 RECT 2.305 1.29 2.405 2.75 ;
 RECT 1.825 1.35 1.925 2.75 ;
 RECT 1.355 0.565 1.455 1.93 ;
 RECT 1.165 1.93 1.455 2.16 ;
 LAYER CO ;
 RECT 2.05 2.325 2.18 2.455 ;
 RECT 2.535 2.36 2.665 2.49 ;
 RECT 2.535 2.08 2.665 2.21 ;
 RECT 2.535 1.81 2.665 1.94 ;
 RECT 1.575 2.33 1.705 2.46 ;
 RECT 1.575 1.805 1.705 1.935 ;
 RECT 2.525 0.595 2.655 0.725 ;
 RECT 2.535 1.545 2.665 1.675 ;
 RECT 2.535 1.545 2.665 1.675 ;
 RECT 2.05 1.545 2.18 1.675 ;
 RECT 0.635 0.785 0.765 0.915 ;
 RECT 0.635 1.67 0.765 1.8 ;
 RECT 1.105 1.545 1.235 1.675 ;
 RECT 1.215 1.97 1.345 2.1 ;
 RECT 2.05 1.805 2.18 1.935 ;
 RECT 0.805 1.17 0.935 1.3 ;
 RECT 2.05 2.065 2.18 2.195 ;
 RECT 1.575 1.545 1.705 1.675 ;
 RECT 1.575 0.595 1.705 0.725 ;
 RECT 2.05 0.595 2.18 0.725 ;
 RECT 1.685 1.17 1.815 1.3 ;
 RECT 1.575 2.065 1.705 2.195 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 0.21 1.545 0.34 1.675 ;
 RECT 0.21 1.805 0.34 1.935 ;
 RECT 0.21 2.065 0.34 2.195 ;
 LAYER M1 ;
 RECT 0.585 0.78 1.24 0.92 ;
 RECT 1.1 1.5 1.24 1.725 ;
 RECT 1.1 0.51 1.24 1.5 ;
 RECT 1.635 1.12 1.865 1.35 ;
 RECT 1.1 1.21 1.865 1.35 ;
 END
END AND2X2

MACRO AND2X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.06 1.06 2.395 1.125 ;
 RECT 2.06 0.78 2.395 0.92 ;
 RECT 3.05 1.06 3.19 2.565 ;
 RECT 2.06 0.92 3.19 1.06 ;
 RECT 3.05 0.505 3.19 0.92 ;
 RECT 2.06 1.125 2.2 2.565 ;
 RECT 2.06 0.54 2.2 0.78 ;
 END
 ANTENNADIFFAREA 1.156 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 RECT 0.205 1.495 0.345 2.8 ;
 RECT 0.64 1.6 0.78 2.8 ;
 RECT 1.58 1.495 1.72 2.8 ;
 RECT 2.545 1.495 2.685 2.8 ;
 RECT 3.535 1.495 3.675 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.52 1.135 0.965 1.4 ;
 END
 ANTENNAGATEAREA 0.062 ;
 END IN1

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 0.22 0.08 0.36 0.755 ;
 RECT 1.58 0.08 1.72 0.945 ;
 RECT 2.535 0.08 2.675 0.77 ;
 RECT 3.53 0.08 3.67 0.765 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.035 1.93 1.405 2.365 ;
 END
 ANTENNAGATEAREA 0.062 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 0.76 1.135 0.995 1.365 ;
 RECT 0.895 0.535 0.995 1.135 ;
 RECT 0.895 1.365 0.995 2.045 ;
 RECT 1.84 0.365 1.94 1.12 ;
 RECT 1.645 1.12 1.94 1.19 ;
 RECT 3.305 0.365 3.405 1.19 ;
 RECT 1.645 1.19 3.405 1.29 ;
 RECT 3.305 1.29 3.405 2.75 ;
 RECT 2.825 0.365 2.925 1.19 ;
 RECT 2.825 1.29 2.925 2.75 ;
 RECT 1.645 1.29 1.94 1.35 ;
 RECT 1.84 1.35 1.94 2.75 ;
 RECT 2.32 0.365 2.42 1.19 ;
 RECT 2.32 1.29 2.42 2.75 ;
 RECT 1.365 0.535 1.465 1.93 ;
 RECT 1.175 1.93 1.465 2.16 ;
 LAYER CO ;
 RECT 1.585 2.355 1.715 2.485 ;
 RECT 1.585 2.075 1.715 2.205 ;
 RECT 1.585 1.805 1.715 1.935 ;
 RECT 3.54 2.335 3.67 2.465 ;
 RECT 3.54 2.075 3.67 2.205 ;
 RECT 3.54 1.81 3.67 1.94 ;
 RECT 3.055 2.325 3.185 2.455 ;
 RECT 2.55 2.34 2.68 2.47 ;
 RECT 2.55 2.065 2.68 2.195 ;
 RECT 2.55 1.805 2.68 1.935 ;
 RECT 2.065 2.375 2.195 2.505 ;
 RECT 3.535 0.585 3.665 0.715 ;
 RECT 3.54 1.545 3.67 1.675 ;
 RECT 3.055 1.545 3.185 1.675 ;
 RECT 3.055 2.065 3.185 2.195 ;
 RECT 3.055 0.585 3.185 0.715 ;
 RECT 3.055 1.805 3.185 1.935 ;
 RECT 2.065 1.545 2.195 1.675 ;
 RECT 1.225 1.97 1.355 2.1 ;
 RECT 0.21 2.065 0.34 2.195 ;
 RECT 2.55 1.545 2.68 1.675 ;
 RECT 0.645 0.775 0.775 0.905 ;
 RECT 2.065 1.805 2.195 1.935 ;
 RECT 1.695 1.17 1.825 1.3 ;
 RECT 2.54 0.585 2.67 0.715 ;
 RECT 0.645 1.65 0.775 1.78 ;
 RECT 2.065 0.68 2.195 0.81 ;
 RECT 0.81 1.185 0.94 1.315 ;
 RECT 0.21 1.805 0.34 1.935 ;
 RECT 2.065 2.065 2.195 2.195 ;
 RECT 0.21 1.545 0.34 1.675 ;
 RECT 1.585 1.545 1.715 1.675 ;
 RECT 1.585 0.755 1.715 0.885 ;
 RECT 1.585 1.545 1.715 1.675 ;
 RECT 1.115 1.545 1.245 1.675 ;
 RECT 2.55 1.545 2.68 1.675 ;
 RECT 0.225 0.315 0.355 0.445 ;
 RECT 0.225 0.575 0.355 0.705 ;
 LAYER M1 ;
 RECT 1.11 1.5 1.25 1.725 ;
 RECT 1.11 0.75 1.25 1.5 ;
 RECT 0.595 0.77 1.25 0.91 ;
 RECT 1.645 1.12 1.845 1.35 ;
 RECT 1.11 1.21 1.845 1.35 ;
 END
END AND2X4

MACRO AND3X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.88 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.395 2.1 1.72 2.36 ;
 END
 ANTENNAGATEAREA 0.051 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.52 2.42 0.92 2.66 ;
 END
 ANTENNAGATEAREA 0.051 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.48 0.835 1.92 1.075 ;
 END
 ANTENNAGATEAREA 0.051 ;
 END IN3

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.44 0.475 2.75 0.85 ;
 RECT 2.61 0.85 2.75 2.59 ;
 END
 ANTENNADIFFAREA 0.577 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.88 2.96 ;
 RECT 2.06 1.52 2.2 2.8 ;
 RECT 1.115 1.53 1.255 2.8 ;
 RECT 0.23 1.51 0.37 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.88 0.08 ;
 RECT 2.06 0.08 2.2 0.77 ;
 RECT 0.23 0.08 0.37 0.845 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 1.84 0.34 1.94 0.835 ;
 RECT 1.84 1.065 1.94 1.935 ;
 RECT 1.71 0.835 1.94 1.065 ;
 RECT 0.9 0.335 1 2.43 ;
 RECT 0.685 2.43 1 2.65 ;
 RECT 0.685 2.65 0.915 2.66 ;
 RECT 2.315 0.335 2.415 1.15 ;
 RECT 2.315 1.38 2.415 2.755 ;
 RECT 2.12 1.15 2.415 1.38 ;
 RECT 1.37 0.335 1.47 2.115 ;
 RECT 1.37 2.115 1.6 2.345 ;
 LAYER CO ;
 RECT 2.615 2.345 2.745 2.475 ;
 RECT 0.235 0.405 0.365 0.535 ;
 RECT 0.235 0.665 0.365 0.795 ;
 RECT 0.235 1.56 0.365 1.69 ;
 RECT 0.235 2.08 0.365 2.21 ;
 RECT 0.235 1.82 0.365 1.95 ;
 RECT 1.42 2.165 1.55 2.295 ;
 RECT 2.065 1.57 2.195 1.7 ;
 RECT 2.17 1.2 2.3 1.33 ;
 RECT 0.65 0.56 0.78 0.69 ;
 RECT 0.735 2.48 0.865 2.61 ;
 RECT 2.615 2.075 2.745 2.205 ;
 RECT 2.615 1.555 2.745 1.685 ;
 RECT 0.65 1.555 0.78 1.685 ;
 RECT 1.12 1.58 1.25 1.71 ;
 RECT 2.065 0.56 2.195 0.69 ;
 RECT 2.615 1.815 2.745 1.945 ;
 RECT 1.75 0.885 1.88 1.015 ;
 RECT 2.615 0.56 2.745 0.69 ;
 RECT 1.59 1.51 1.72 1.64 ;
 LAYER M1 ;
 RECT 0.6 0.555 1.215 0.7 ;
 RECT 1.075 0.555 1.215 1.355 ;
 RECT 0.645 1.235 0.785 1.735 ;
 RECT 1.585 1.235 1.725 1.69 ;
 RECT 2.12 1.19 2.35 1.38 ;
 RECT 0.64 1.235 2.35 1.375 ;
 END
END AND3X1

MACRO AND3X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 1.995 0.34 2.265 0.48 ;
 RECT 0.23 0.08 0.37 0.85 ;
 RECT 3.09 0.08 3.23 0.555 ;
 RECT 2.06 0.08 2.2 0.34 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.52 2.1 0.875 2.36 ;
 END
 ANTENNAGATEAREA 0.052 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 2.06 1.525 2.2 2.8 ;
 RECT 1.115 1.535 1.255 2.8 ;
 RECT 0.23 1.515 0.37 2.8 ;
 RECT 3.09 1.745 3.23 2.8 ;
 END
 END VDD

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.705 0.835 2.04 1.08 ;
 END
 ANTENNAGATEAREA 0.052 ;
 END IN3

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.615 1.155 3.015 1.4 ;
 RECT 2.615 1.4 2.755 2.595 ;
 RECT 2.615 0.27 2.755 1.155 ;
 END
 ANTENNADIFFAREA 0.556 ;
 END Q

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.395 1.8 1.805 2.075 ;
 END
 ANTENNAGATEAREA 0.052 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 1.84 0.105 1.94 0.84 ;
 RECT 1.84 1.07 1.94 1.96 ;
 RECT 1.71 0.84 1.94 1.07 ;
 RECT 0.9 0.105 1 2.105 ;
 RECT 0.685 2.105 1 2.335 ;
 RECT 2.18 1.215 2.97 1.315 ;
 RECT 2.18 1.155 2.495 1.215 ;
 RECT 2.87 0.105 2.97 1.215 ;
 RECT 2.18 1.315 2.495 1.385 ;
 RECT 2.395 0.105 2.495 1.155 ;
 RECT 2.87 1.315 2.97 2.76 ;
 RECT 2.395 1.385 2.495 2.76 ;
 RECT 1.37 0.105 1.47 1.835 ;
 RECT 1.37 1.835 1.6 2.065 ;
 LAYER CO ;
 RECT 3.095 2.4 3.225 2.53 ;
 RECT 3.095 2.14 3.225 2.27 ;
 RECT 3.095 1.845 3.225 1.975 ;
 RECT 3.095 0.345 3.225 0.475 ;
 RECT 2.62 1.56 2.75 1.69 ;
 RECT 0.65 1.56 0.78 1.69 ;
 RECT 2.62 1.82 2.75 1.95 ;
 RECT 0.235 1.825 0.365 1.955 ;
 RECT 2.62 2.08 2.75 2.21 ;
 RECT 1.77 0.89 1.9 1.02 ;
 RECT 1.12 1.585 1.25 1.715 ;
 RECT 1.59 1.495 1.72 1.625 ;
 RECT 2.065 1.575 2.195 1.705 ;
 RECT 0.65 0.495 0.78 0.625 ;
 RECT 2.065 0.345 2.195 0.475 ;
 RECT 2.62 0.415 2.75 0.545 ;
 RECT 1.42 1.885 1.55 2.015 ;
 RECT 0.735 2.155 0.865 2.285 ;
 RECT 0.235 0.41 0.365 0.54 ;
 RECT 0.235 0.67 0.365 0.8 ;
 RECT 2.62 2.35 2.75 2.48 ;
 RECT 0.235 1.565 0.365 1.695 ;
 RECT 0.235 2.085 0.365 2.215 ;
 RECT 2.23 1.205 2.36 1.335 ;
 LAYER M1 ;
 RECT 0.6 0.485 1.215 0.63 ;
 RECT 1.075 0.47 1.215 1.36 ;
 RECT 0.645 1.24 0.785 1.74 ;
 RECT 1.52 1.49 1.79 1.63 ;
 RECT 1.52 1.24 1.79 1.63 ;
 RECT 2.18 1.195 2.41 1.385 ;
 RECT 0.64 1.24 2.41 1.38 ;
 END
END AND3X2

MACRO AND3X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.58 1.425 3.72 2.59 ;
 RECT 3.58 1.12 3.955 1.425 ;
 RECT 2.615 1.12 2.755 2.59 ;
 RECT 2.615 0.265 2.755 0.98 ;
 RECT 2.615 0.98 3.72 1.12 ;
 RECT 3.58 0.265 3.72 0.98 ;
 END
 ANTENNADIFFAREA 1.112 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 2.06 1.52 2.2 2.8 ;
 RECT 1.115 1.53 1.255 2.8 ;
 RECT 0.23 1.51 0.37 2.8 ;
 RECT 3.09 1.52 3.23 2.8 ;
 RECT 4.055 1.755 4.195 2.8 ;
 END
 END VDD

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.725 0.845 2.05 1.08 ;
 END
 ANTENNAGATEAREA 0.052 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 0.23 0.08 0.37 0.845 ;
 RECT 2.06 0.08 2.2 0.55 ;
 RECT 3.09 0.08 3.23 0.55 ;
 RECT 4.055 0.08 4.195 0.55 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.395 2.08 1.72 2.36 ;
 END
 ANTENNAGATEAREA 0.052 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.52 1.8 0.935 2.125 ;
 END
 ANTENNAGATEAREA 0.052 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 1.37 0.1 1.47 2.115 ;
 RECT 1.37 2.115 1.6 2.345 ;
 RECT 0.9 0.1 1 1.885 ;
 RECT 0.685 1.885 1 2.115 ;
 RECT 2.245 1.21 3.935 1.31 ;
 RECT 3.36 0.1 3.46 1.21 ;
 RECT 3.835 0.1 3.935 1.21 ;
 RECT 2.87 0.1 2.97 1.21 ;
 RECT 2.395 0.1 2.495 1.15 ;
 RECT 2.245 1.15 2.495 1.21 ;
 RECT 2.245 1.31 2.495 1.38 ;
 RECT 3.835 1.31 3.935 2.755 ;
 RECT 3.36 1.31 3.46 2.755 ;
 RECT 2.87 1.31 2.97 2.755 ;
 RECT 2.395 1.38 2.495 2.755 ;
 RECT 1.84 0.1 1.94 0.845 ;
 RECT 1.84 1.075 1.94 1.955 ;
 RECT 1.73 0.845 1.96 1.075 ;
 LAYER CO ;
 RECT 3.095 2.135 3.225 2.265 ;
 RECT 3.585 2.345 3.715 2.475 ;
 RECT 4.06 0.32 4.19 0.45 ;
 RECT 4.06 2.395 4.19 2.525 ;
 RECT 4.06 2.135 4.19 2.265 ;
 RECT 3.585 2.075 3.715 2.205 ;
 RECT 3.585 1.815 3.715 1.945 ;
 RECT 3.585 0.39 3.715 0.52 ;
 RECT 4.06 1.84 4.19 1.97 ;
 RECT 3.585 1.555 3.715 1.685 ;
 RECT 1.78 0.895 1.91 1.025 ;
 RECT 0.235 0.405 0.365 0.535 ;
 RECT 2.065 0.32 2.195 0.45 ;
 RECT 2.62 1.815 2.75 1.945 ;
 RECT 2.62 0.39 2.75 0.52 ;
 RECT 0.65 1.525 0.78 1.655 ;
 RECT 0.735 1.935 0.865 2.065 ;
 RECT 3.095 1.84 3.225 1.97 ;
 RECT 2.62 2.345 2.75 2.475 ;
 RECT 3.095 2.395 3.225 2.525 ;
 RECT 2.295 1.2 2.425 1.33 ;
 RECT 3.095 1.57 3.225 1.7 ;
 RECT 0.235 1.82 0.365 1.95 ;
 RECT 1.12 1.58 1.25 1.71 ;
 RECT 0.235 1.56 0.365 1.69 ;
 RECT 2.62 1.555 2.75 1.685 ;
 RECT 3.095 0.32 3.225 0.45 ;
 RECT 0.235 2.08 0.365 2.21 ;
 RECT 2.62 2.075 2.75 2.205 ;
 RECT 1.59 1.49 1.72 1.62 ;
 RECT 1.42 2.165 1.55 2.295 ;
 RECT 2.065 1.57 2.195 1.7 ;
 RECT 0.235 0.665 0.365 0.795 ;
 RECT 0.65 0.47 0.78 0.6 ;
 LAYER M1 ;
 RECT 1.075 0.465 1.215 1.355 ;
 RECT 0.6 0.46 1.215 0.605 ;
 RECT 1.585 1.235 1.725 1.67 ;
 RECT 0.58 1.52 0.85 1.66 ;
 RECT 0.645 1.235 0.785 1.66 ;
 RECT 2.245 1.19 2.475 1.38 ;
 RECT 0.64 1.235 2.415 1.375 ;
 END
END AND3X4

MACRO NOR3X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 2.88 ;
 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.87 1.12 4.205 1.36 ;
 RECT 3.87 1.36 4.01 2.56 ;
 RECT 3.87 0.31 4.01 1.12 ;
 END
 ANTENNADIFFAREA 0.646 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 2.39 1.565 2.53 2.8 ;
 RECT 3.39 1.515 3.53 2.8 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 4.365 1.39 4.505 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.275 1.04 1.625 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.69 1.04 1.135 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.12 0.745 2.36 1.095 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 2.3 0.08 2.44 0.555 ;
 RECT 1.34 0.08 1.48 0.505 ;
 RECT 3.4 0.08 3.54 0.875 ;
 RECT 0.31 0.08 0.45 0.755 ;
 RECT 4.37 0.08 4.51 0.875 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 3.495 1.12 3.755 1.21 ;
 RECT 3.495 1.31 3.755 1.35 ;
 RECT 3.495 1.21 4.245 1.31 ;
 RECT 4.145 0.155 4.245 1.21 ;
 RECT 4.145 1.31 4.245 2.75 ;
 RECT 3.655 0.155 3.755 1.12 ;
 RECT 3.655 1.35 3.755 2.75 ;
 RECT 1.4 1.14 1.705 1.37 ;
 RECT 1.605 0.105 1.705 1.14 ;
 RECT 1.605 1.37 1.705 2.755 ;
 RECT 0.89 1.12 1.22 1.35 ;
 RECT 1.12 0.105 1.22 1.12 ;
 RECT 1.12 1.35 1.22 2.76 ;
 RECT 2.715 0.105 2.815 1.12 ;
 RECT 2.715 1.35 2.815 2.18 ;
 RECT 2.61 1.12 2.84 1.35 ;
 RECT 2.085 0.105 2.185 0.745 ;
 RECT 2.085 0.975 2.185 2.76 ;
 RECT 2.085 0.745 2.315 0.975 ;
 LAYER CO ;
 RECT 3.875 2.28 4.005 2.41 ;
 RECT 3.395 1.585 3.525 1.715 ;
 RECT 3.395 1.845 3.525 1.975 ;
 RECT 3.395 2.11 3.525 2.24 ;
 RECT 4.37 1.5 4.5 1.63 ;
 RECT 4.37 1.775 4.5 1.905 ;
 RECT 4.37 2.065 4.5 2.195 ;
 RECT 2.395 1.84 2.525 1.97 ;
 RECT 2.395 2.1 2.525 2.23 ;
 RECT 4.375 0.405 4.505 0.535 ;
 RECT 4.375 0.68 4.505 0.81 ;
 RECT 4.37 2.34 4.5 2.47 ;
 RECT 3.875 1.5 4.005 1.63 ;
 RECT 3.405 0.405 3.535 0.535 ;
 RECT 3.395 2.375 3.525 2.505 ;
 RECT 3.545 1.17 3.675 1.3 ;
 RECT 2.135 0.795 2.265 0.925 ;
 RECT 2.95 1.545 3.08 1.675 ;
 RECT 1.345 0.325 1.475 0.455 ;
 RECT 2.305 0.325 2.435 0.455 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 0.94 1.17 1.07 1.3 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 3.405 0.68 3.535 0.81 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 2.66 1.17 2.79 1.3 ;
 RECT 3.875 1.76 4.005 1.89 ;
 RECT 2.395 2.36 2.525 2.49 ;
 RECT 1.83 0.325 1.96 0.455 ;
 RECT 2.95 1.805 3.08 1.935 ;
 RECT 0.87 1.545 1 1.675 ;
 RECT 1.45 1.19 1.58 1.32 ;
 RECT 2.95 0.325 3.08 0.455 ;
 RECT 0.865 0.325 0.995 0.455 ;
 RECT 3.875 0.46 4.005 0.59 ;
 RECT 3.875 2.02 4.005 2.15 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 0.315 0.315 0.445 0.445 ;
 LAYER M1 ;
 RECT 0.86 0.26 1 0.685 ;
 RECT 1.82 0.825 1.96 1.255 ;
 RECT 1.82 1.395 1.96 1.54 ;
 RECT 1.82 0.505 1.96 0.685 ;
 RECT 0.86 0.685 1.96 0.825 ;
 RECT 0.725 1.54 1.96 1.68 ;
 RECT 1.815 0.275 1.975 0.505 ;
 RECT 2.645 1.12 2.8 1.255 ;
 RECT 1.82 1.255 2.8 1.395 ;
 RECT 2.945 0.275 3.085 1.185 ;
 RECT 2.945 1.325 3.085 2.05 ;
 RECT 2.945 1.185 3.685 1.325 ;
 RECT 3.53 1.12 3.685 1.185 ;
 RECT 3.53 1.325 3.685 1.35 ;
 END
END NOR3X2

MACRO NOR3X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.76 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.76 2.96 ;
 RECT 4.365 1.455 4.505 2.8 ;
 RECT 3.39 1.5 3.53 2.8 ;
 RECT 2.39 1.535 2.53 2.8 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 5.35 1.525 5.49 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.76 0.08 ;
 RECT 1.34 0.08 1.48 0.505 ;
 RECT 4.37 0.08 4.51 0.875 ;
 RECT 2.3 0.08 2.44 0.555 ;
 RECT 0.31 0.08 0.45 0.755 ;
 RECT 3.4 0.08 3.54 0.875 ;
 RECT 5.37 0.08 5.51 0.875 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.84 0.84 5.08 1.045 ;
 RECT 4.86 1.185 5 2.57 ;
 RECT 3.87 1.045 5.08 1.165 ;
 RECT 3.87 0.31 4.01 1.045 ;
 RECT 4.86 0.31 5 0.84 ;
 RECT 3.87 1.185 4.01 2.62 ;
 RECT 3.87 1.165 5 1.185 ;
 END
 ANTENNADIFFAREA 1.302 ;
 END QN

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.325 1.04 1.68 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.84 1.04 1.14 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.125 0.745 2.52 1.08 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN3

 OBS
 LAYER PO ;
 RECT 0.895 1.14 1.22 1.37 ;
 RECT 1.12 0.105 1.22 1.14 ;
 RECT 1.12 1.37 1.22 2.755 ;
 RECT 3.495 1.085 3.755 1.21 ;
 RECT 3.495 1.31 3.755 1.315 ;
 RECT 3.495 1.21 5.225 1.31 ;
 RECT 5.125 0.155 5.225 1.21 ;
 RECT 5.125 1.31 5.225 2.76 ;
 RECT 4.63 0.155 4.73 1.21 ;
 RECT 4.63 1.31 4.73 2.76 ;
 RECT 4.145 0.155 4.245 1.21 ;
 RECT 4.145 1.31 4.245 2.76 ;
 RECT 3.655 0.155 3.755 1.085 ;
 RECT 3.655 1.315 3.755 2.76 ;
 RECT 1.445 1.14 1.705 1.37 ;
 RECT 1.605 0.105 1.705 1.14 ;
 RECT 1.605 1.37 1.705 2.755 ;
 RECT 2.715 0.105 2.815 1.12 ;
 RECT 2.715 1.35 2.815 2.76 ;
 RECT 2.715 1.12 2.945 1.35 ;
 RECT 2.085 0.105 2.185 0.745 ;
 RECT 2.085 0.975 2.185 2.75 ;
 RECT 2.085 0.745 2.315 0.975 ;
 LAYER CO ;
 RECT 5.375 0.68 5.505 0.81 ;
 RECT 5.375 0.405 5.505 0.535 ;
 RECT 5.355 2.19 5.485 2.32 ;
 RECT 4.865 0.46 4.995 0.59 ;
 RECT 4.865 1.51 4.995 1.64 ;
 RECT 4.865 1.77 4.995 1.9 ;
 RECT 4.865 2.03 4.995 2.16 ;
 RECT 2.95 2.09 3.08 2.22 ;
 RECT 4.375 0.405 4.505 0.535 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 2.395 2.225 2.525 2.355 ;
 RECT 0.945 1.19 1.075 1.32 ;
 RECT 2.95 0.325 3.08 0.455 ;
 RECT 2.305 0.325 2.435 0.455 ;
 RECT 3.875 1.77 4.005 1.9 ;
 RECT 4.375 0.68 4.505 0.81 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 3.395 2.19 3.525 2.32 ;
 RECT 3.875 0.46 4.005 0.59 ;
 RECT 2.135 0.795 2.265 0.925 ;
 RECT 4.37 2.19 4.5 2.32 ;
 RECT 3.405 0.405 3.535 0.535 ;
 RECT 0.865 0.325 0.995 0.455 ;
 RECT 1.83 0.325 1.96 0.455 ;
 RECT 1.345 0.325 1.475 0.455 ;
 RECT 3.875 1.51 4.005 1.64 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 3.875 2.03 4.005 2.16 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 1.495 1.19 1.625 1.32 ;
 RECT 2.765 1.17 2.895 1.3 ;
 RECT 3.545 1.135 3.675 1.265 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 0.87 1.545 1 1.675 ;
 RECT 3.405 0.68 3.535 0.81 ;
 RECT 2.95 2.35 3.08 2.48 ;
 RECT 5.355 1.64 5.485 1.77 ;
 RECT 5.355 1.925 5.485 2.055 ;
 RECT 5.355 2.19 5.485 2.32 ;
 RECT 4.865 2.29 4.995 2.42 ;
 RECT 4.37 1.65 4.5 1.78 ;
 RECT 4.37 1.925 4.5 2.055 ;
 RECT 3.875 2.29 4.005 2.42 ;
 RECT 3.395 1.64 3.525 1.77 ;
 RECT 3.395 1.925 3.525 2.055 ;
 RECT 2.395 1.69 2.525 1.82 ;
 RECT 2.395 1.96 2.525 2.09 ;
 LAYER M1 ;
 RECT 0.86 0.26 1 0.685 ;
 RECT 1.82 0.825 1.96 1.255 ;
 RECT 1.82 1.395 1.96 1.54 ;
 RECT 1.82 0.505 1.96 0.685 ;
 RECT 0.86 0.685 1.96 0.825 ;
 RECT 0.725 1.54 1.96 1.68 ;
 RECT 1.815 0.275 1.975 0.505 ;
 RECT 1.82 1.255 2.935 1.395 ;
 RECT 2.72 1.12 2.935 1.255 ;
 RECT 3.085 0.46 3.225 1.185 ;
 RECT 3.085 1.325 3.225 1.78 ;
 RECT 2.945 1.92 3.085 2.55 ;
 RECT 2.945 1.78 3.225 1.92 ;
 RECT 2.88 0.32 3.225 0.46 ;
 RECT 3.085 1.185 3.725 1.325 ;
 RECT 3.495 1.085 3.725 1.185 ;
 END
END NOR3X4

MACRO AND4X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.96 0.755 2.265 1.08 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN3

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 0.835 1.055 1.085 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN1

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.28 1.865 2.545 2.365 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN4

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 3.725 0.08 3.865 0.505 ;
 RECT 0.365 0.08 0.505 0.91 ;
 RECT 2.67 0.08 2.81 0.505 ;
 RECT 4.72 0.08 4.86 0.505 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.22 0.835 3.485 0.905 ;
 RECT 3.22 1.075 3.36 2.57 ;
 RECT 3.22 1.045 3.485 1.075 ;
 RECT 4.25 1.045 4.39 2.585 ;
 RECT 3.22 0.905 4.39 1.045 ;
 RECT 4.25 0.27 4.39 0.905 ;
 RECT 3.22 0.27 3.36 0.835 ;
 END
 ANTENNADIFFAREA 1.194 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 1.675 1.555 1.905 1.695 ;
 RECT 2.73 1.515 2.87 2.8 ;
 RECT 0.37 1.495 0.51 2.8 ;
 RECT 3.73 1.515 3.87 2.8 ;
 RECT 4.725 1.515 4.865 2.8 ;
 RECT 0.78 1.51 0.92 2.8 ;
 RECT 1.72 1.695 1.86 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.86 1.58 2.38 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 1.975 0.26 2.075 0.775 ;
 RECT 1.975 0.775 2.21 1.005 ;
 RECT 1.975 1.005 2.075 1.915 ;
 RECT 2.45 0.265 2.55 1.865 ;
 RECT 2.32 1.865 2.55 2.095 ;
 RECT 1.035 0.255 1.135 0.845 ;
 RECT 0.825 0.845 1.135 1.075 ;
 RECT 1.035 1.075 1.135 1.92 ;
 RECT 2.845 1.2 4.605 1.3 ;
 RECT 4.505 0.105 4.605 1.2 ;
 RECT 4.02 0.1 4.12 1.2 ;
 RECT 3.49 0.105 3.59 1.2 ;
 RECT 3 0.105 3.1 1.15 ;
 RECT 2.845 1.15 3.1 1.2 ;
 RECT 2.845 1.3 3.1 1.38 ;
 RECT 4.505 1.3 4.605 2.76 ;
 RECT 4.02 1.3 4.12 2.76 ;
 RECT 3.49 1.3 3.59 2.76 ;
 RECT 3 1.38 3.1 2.76 ;
 RECT 1.505 0.26 1.605 1.86 ;
 RECT 1.375 1.86 1.605 2.09 ;
 LAYER CO ;
 RECT 4.73 2.39 4.86 2.52 ;
 RECT 4.73 2.115 4.86 2.245 ;
 RECT 4.73 1.835 4.86 1.965 ;
 RECT 4.255 2.34 4.385 2.47 ;
 RECT 3.735 2.385 3.865 2.515 ;
 RECT 3.735 2.095 3.865 2.225 ;
 RECT 3.735 1.825 3.865 1.955 ;
 RECT 3.225 2.355 3.355 2.485 ;
 RECT 2.735 2.38 2.865 2.51 ;
 RECT 2.735 2.11 2.865 2.24 ;
 RECT 2.735 1.835 2.865 1.965 ;
 RECT 4.73 1.565 4.86 1.695 ;
 RECT 4.725 0.325 4.855 0.455 ;
 RECT 4.255 1.56 4.385 1.69 ;
 RECT 4.255 0.325 4.385 0.455 ;
 RECT 4.255 1.82 4.385 1.95 ;
 RECT 4.255 2.08 4.385 2.21 ;
 RECT 0.875 0.895 1.005 1.025 ;
 RECT 1.425 1.91 1.555 2.04 ;
 RECT 3.73 0.325 3.86 0.455 ;
 RECT 0.37 0.47 0.5 0.6 ;
 RECT 2.015 0.825 2.145 0.955 ;
 RECT 3.735 1.565 3.865 1.695 ;
 RECT 0.375 2.065 0.505 2.195 ;
 RECT 0.785 1.56 0.915 1.69 ;
 RECT 0.375 1.805 0.505 1.935 ;
 RECT 0.375 1.545 0.505 1.675 ;
 RECT 2.895 1.2 3.025 1.33 ;
 RECT 3.225 1.82 3.355 1.95 ;
 RECT 3.225 2.08 3.355 2.21 ;
 RECT 1.255 1.51 1.385 1.64 ;
 RECT 0.37 0.73 0.5 0.86 ;
 RECT 1.725 1.56 1.855 1.69 ;
 RECT 2.37 1.915 2.5 2.045 ;
 RECT 2.735 1.565 2.865 1.695 ;
 RECT 0.785 0.485 0.915 0.615 ;
 RECT 3.225 0.325 3.355 0.455 ;
 RECT 2.195 1.505 2.325 1.635 ;
 RECT 3.225 1.56 3.355 1.69 ;
 RECT 2.675 0.325 2.805 0.455 ;
 RECT 1.725 1.56 1.855 1.69 ;
 LAYER M1 ;
 RECT 0.905 0.495 1.81 0.635 ;
 RECT 1.67 0.55 1.81 1.345 ;
 RECT 0.78 0.435 0.92 0.665 ;
 RECT 1.25 1.245 1.39 1.695 ;
 RECT 1.25 1.235 2.33 1.375 ;
 RECT 2.19 1.24 2.33 1.685 ;
 RECT 2.845 1.19 3.075 1.34 ;
 RECT 2.195 1.235 3.075 1.375 ;
 END
END AND4X4

MACRO AO21X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 3.14 1.585 3.28 2.8 ;
 RECT 2.725 1.785 2.865 2.8 ;
 RECT 0.115 1.825 0.255 2.8 ;
 RECT 1.055 1.825 1.195 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.12 0.46 1.4 ;
 END
 ANTENNAGATEAREA 0.075 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.64 1.155 0.96 1.4 ;
 END
 ANTENNAGATEAREA 0.075 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.195 1.155 1.56 1.4 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN3

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.255 1.08 2.395 2.44 ;
 RECT 2.255 0.84 2.52 1.08 ;
 RECT 2.255 0.49 2.395 0.84 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 2.725 0.08 2.865 0.735 ;
 RECT 3.14 0.08 3.28 0.78 ;
 RECT 1.365 0.08 1.505 0.715 ;
 RECT 0.115 0.08 0.255 0.71 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 1.15 0.305 1.25 1.165 ;
 RECT 1.67 1.38 1.77 2.35 ;
 RECT 1.15 1.165 1.38 1.28 ;
 RECT 1.15 1.28 1.77 1.38 ;
 RECT 0.37 1.39 0.47 2.24 ;
 RECT 0.37 0.305 0.47 1.18 ;
 RECT 0.23 1.18 0.47 1.39 ;
 RECT 0.68 1.27 0.94 1.435 ;
 RECT 0.68 0.305 0.78 1.225 ;
 RECT 0.84 1.435 0.94 2.24 ;
 RECT 0.68 1.225 0.91 1.27 ;
 RECT 2.51 0.315 2.61 0.985 ;
 RECT 2.51 1.085 2.61 2.74 ;
 RECT 1.84 0.875 2.07 0.985 ;
 RECT 1.84 0.985 2.61 1.085 ;
 LAYER CO ;
 RECT 2.73 1.84 2.86 1.97 ;
 RECT 2.73 2.1 2.86 2.23 ;
 RECT 2.26 1.735 2.39 1.865 ;
 RECT 2.26 2 2.39 2.13 ;
 RECT 1.89 1.96 2.02 2.09 ;
 RECT 0.12 1.88 0.25 2.01 ;
 RECT 3.145 1.895 3.275 2.025 ;
 RECT 1.2 1.205 1.33 1.335 ;
 RECT 0.73 1.265 0.86 1.395 ;
 RECT 2.73 0.555 2.86 0.685 ;
 RECT 2.26 2.26 2.39 2.39 ;
 RECT 1.06 1.88 1.19 2.01 ;
 RECT 1.37 0.535 1.5 0.665 ;
 RECT 0.59 1.88 0.72 2.01 ;
 RECT 0.12 0.525 0.25 0.655 ;
 RECT 3.145 2.155 3.275 2.285 ;
 RECT 0.9 0.535 1.03 0.665 ;
 RECT 3.145 0.34 3.275 0.47 ;
 RECT 1.89 1.7 2.02 1.83 ;
 RECT 2.26 0.555 2.39 0.685 ;
 RECT 1.89 0.915 2.02 1.045 ;
 RECT 3.145 1.635 3.275 1.765 ;
 RECT 1.42 1.75 1.55 1.88 ;
 RECT 3.145 0.6 3.275 0.73 ;
 RECT 2.73 2.36 2.86 2.49 ;
 RECT 0.28 1.22 0.41 1.35 ;
 LAYER M1 ;
 RECT 0.585 1.685 0.725 2.075 ;
 RECT 1.415 1.685 1.555 1.935 ;
 RECT 0.585 1.545 1.555 1.685 ;
 RECT 0.895 0.48 1.035 0.87 ;
 RECT 1.885 0.865 2.025 0.87 ;
 RECT 1.885 1.01 2.025 2.15 ;
 RECT 0.895 0.87 2.025 1.01 ;
 END
END AO21X1

MACRO AO21X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 1.16 0.48 1.415 ;
 END
 ANTENNAGATEAREA 0.075 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.4 3.335 2.44 ;
 RECT 3.195 1.16 3.48 1.4 ;
 RECT 2.255 1.105 2.395 2.44 ;
 RECT 2.255 0.965 3.335 1.105 ;
 RECT 2.255 0.51 2.395 0.965 ;
 RECT 3.195 1.105 3.335 1.16 ;
 RECT 3.195 0.51 3.335 0.965 ;
 END
 ANTENNADIFFAREA 0.93 ;
 END Q

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.195 1.155 1.56 1.4 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 3.61 0.08 3.75 0.78 ;
 RECT 2.725 0.08 2.865 0.76 ;
 RECT 0.115 0.08 0.255 0.675 ;
 RECT 1.365 0.08 1.505 0.655 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.16 1.01 1.455 ;
 END
 ANTENNAGATEAREA 0.075 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 3.61 1.585 3.75 2.8 ;
 RECT 2.725 1.8 2.865 2.8 ;
 RECT 0.115 1.685 0.255 2.8 ;
 RECT 1.055 1.95 1.195 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.37 1.39 0.47 2.36 ;
 RECT 0.37 0.265 0.47 1.18 ;
 RECT 0.23 1.18 0.47 1.39 ;
 RECT 1.15 0.335 1.25 1.165 ;
 RECT 1.67 1.38 1.77 2.475 ;
 RECT 1.15 1.165 1.38 1.28 ;
 RECT 1.15 1.28 1.77 1.38 ;
 RECT 0.68 1.27 0.94 1.435 ;
 RECT 0.68 0.265 0.78 1.225 ;
 RECT 0.84 1.435 0.94 2.36 ;
 RECT 0.68 1.225 0.91 1.27 ;
 RECT 2.98 1.235 3.08 2.74 ;
 RECT 2.51 1.235 2.61 2.74 ;
 RECT 2.98 0.335 3.08 1.135 ;
 RECT 2.51 0.335 2.61 1.135 ;
 RECT 1.97 1.085 2.07 1.135 ;
 RECT 1.97 1.135 3.08 1.235 ;
 RECT 1.84 0.875 2.07 1.085 ;
 LAYER CO ;
 RECT 0.12 1.74 0.25 1.87 ;
 RECT 2.73 1.86 2.86 1.99 ;
 RECT 2.73 2.12 2.86 2.25 ;
 RECT 2.26 1.74 2.39 1.87 ;
 RECT 2.26 2 2.39 2.13 ;
 RECT 3.2 1.74 3.33 1.87 ;
 RECT 3.2 2 3.33 2.13 ;
 RECT 3.2 0.57 3.33 0.7 ;
 RECT 3.2 2.26 3.33 2.39 ;
 RECT 1.42 1.77 1.55 1.9 ;
 RECT 3.615 0.6 3.745 0.73 ;
 RECT 2.26 0.57 2.39 0.7 ;
 RECT 3.615 1.635 3.745 1.765 ;
 RECT 0.12 0.485 0.25 0.615 ;
 RECT 3.615 2.155 3.745 2.285 ;
 RECT 1.89 1.83 2.02 1.96 ;
 RECT 1.89 0.915 2.02 1.045 ;
 RECT 0.59 1.69 0.72 1.82 ;
 RECT 0.12 2 0.25 2.13 ;
 RECT 3.615 1.895 3.745 2.025 ;
 RECT 1.2 1.205 1.33 1.335 ;
 RECT 0.9 0.485 1.03 0.615 ;
 RECT 1.37 0.475 1.5 0.605 ;
 RECT 0.28 1.22 0.41 1.35 ;
 RECT 0.73 1.265 0.86 1.395 ;
 RECT 3.615 0.34 3.745 0.47 ;
 RECT 2.26 2.26 2.39 2.39 ;
 RECT 1.89 2.09 2.02 2.22 ;
 RECT 2.73 2.38 2.86 2.51 ;
 RECT 1.06 2 1.19 2.13 ;
 RECT 2.73 0.57 2.86 0.7 ;
 LAYER M1 ;
 RECT 1.415 1.76 1.555 1.95 ;
 RECT 0.585 1.62 1.555 1.76 ;
 RECT 0.585 1.76 0.725 1.9 ;
 RECT 0.895 0.42 1.035 0.86 ;
 RECT 1.885 1 2.025 2.32 ;
 RECT 0.895 0.86 2.025 1 ;
 END
END AO21X2

MACRO AO221X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.535 0.79 2.855 1.035 ;
 RECT 2.6 1.035 2.84 1.05 ;
 END
 ANTENNAGATEAREA 0.104 ;
 END IN5

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.225 1.16 3.48 1.4 ;
 RECT 3.225 0.495 3.365 1.16 ;
 RECT 3.225 1.4 3.365 2.44 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 3.695 0.08 3.835 0.73 ;
 RECT 4.11 0.08 4.25 0.78 ;
 RECT 0.115 0.08 0.255 0.785 ;
 RECT 1.755 0.08 1.895 0.795 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.47 0.46 1.825 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.48 1.01 1.76 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.195 1.475 1.56 1.72 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN3

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 3.695 1.805 3.835 2.8 ;
 RECT 4.11 1.585 4.25 2.8 ;
 RECT 0.115 2.095 0.255 2.8 ;
 RECT 1.055 2.21 1.195 2.8 ;
 END
 END VDD

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.88 1.48 2.2 1.765 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN4

 OBS
 LAYER PO ;
 RECT 2.01 0.385 2.11 0.985 ;
 RECT 2.615 1.085 2.715 2.78 ;
 RECT 2.01 0.985 2.72 1.01 ;
 RECT 2.49 0.8 2.72 0.985 ;
 RECT 2.01 1.01 2.715 1.085 ;
 RECT 1.98 1.545 2.24 1.755 ;
 RECT 1.54 0.385 1.64 1.265 ;
 RECT 2.14 1.755 2.24 2.78 ;
 RECT 2.14 1.365 2.24 1.545 ;
 RECT 1.54 1.265 2.24 1.365 ;
 RECT 0.68 0.385 0.78 1.545 ;
 RECT 0.84 1.795 0.94 2.77 ;
 RECT 0.68 1.545 0.91 1.695 ;
 RECT 0.68 1.695 0.94 1.795 ;
 RECT 3.48 0.325 3.58 1.315 ;
 RECT 3.48 1.415 3.58 2.78 ;
 RECT 2.9 1.205 3.13 1.315 ;
 RECT 2.9 1.315 3.58 1.415 ;
 RECT 0.23 1.65 0.47 1.86 ;
 RECT 0.37 0.385 0.47 1.65 ;
 RECT 0.37 1.86 0.47 2.77 ;
 RECT 1.15 0.385 1.25 1.485 ;
 RECT 1.67 1.645 1.77 2.78 ;
 RECT 1.15 1.485 1.38 1.545 ;
 RECT 1.15 1.645 1.38 1.695 ;
 RECT 1.15 1.545 1.77 1.645 ;
 LAYER CO ;
 RECT 3.7 1.86 3.83 1.99 ;
 RECT 3.7 2.12 3.83 2.25 ;
 RECT 2.835 1.93 2.965 2.06 ;
 RECT 0.12 2.15 0.25 2.28 ;
 RECT 3.23 1.74 3.36 1.87 ;
 RECT 3.23 2 3.36 2.13 ;
 RECT 4.115 0.6 4.245 0.73 ;
 RECT 4.115 0.34 4.245 0.47 ;
 RECT 2.03 1.585 2.16 1.715 ;
 RECT 2.835 2.19 2.965 2.32 ;
 RECT 2.54 0.84 2.67 0.97 ;
 RECT 2.95 1.245 3.08 1.375 ;
 RECT 0.73 1.585 0.86 1.715 ;
 RECT 1.42 2.26 1.55 2.39 ;
 RECT 1.76 0.615 1.89 0.745 ;
 RECT 3.7 0.545 3.83 0.675 ;
 RECT 1.2 1.525 1.33 1.655 ;
 RECT 2.23 0.615 2.36 0.745 ;
 RECT 1.06 2.26 1.19 2.39 ;
 RECT 4.115 1.635 4.245 1.765 ;
 RECT 2.36 2.26 2.49 2.39 ;
 RECT 0.12 0.605 0.25 0.735 ;
 RECT 0.28 1.69 0.41 1.82 ;
 RECT 0.59 2.26 0.72 2.39 ;
 RECT 3.7 2.38 3.83 2.51 ;
 RECT 3.23 0.545 3.36 0.675 ;
 RECT 0.9 0.605 1.03 0.735 ;
 RECT 3.23 2.26 3.36 2.39 ;
 RECT 0.12 2.41 0.25 2.54 ;
 RECT 4.115 1.895 4.245 2.025 ;
 RECT 1.89 2.075 2.02 2.205 ;
 RECT 4.115 2.155 4.245 2.285 ;
 LAYER M1 ;
 RECT 0.585 2.07 0.725 2.445 ;
 RECT 1.885 2.07 2.025 2.255 ;
 RECT 0.585 1.93 2.025 2.07 ;
 RECT 2.355 2.205 2.495 2.485 ;
 RECT 1.415 2.21 1.555 2.485 ;
 RECT 1.415 2.485 2.495 2.625 ;
 RECT 0.895 0.555 1.035 1.195 ;
 RECT 2.225 0.565 2.365 1.195 ;
 RECT 2.83 1.335 3.085 1.425 ;
 RECT 0.895 1.195 3.085 1.335 ;
 RECT 2.83 1.425 2.97 2.37 ;
 END
END AO221X1

MACRO AO221X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.195 1.475 1.56 1.72 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN3

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 3.2 1.94 3.34 2.8 ;
 RECT 4.665 1.585 4.805 2.8 ;
 RECT 4.14 1.685 4.28 2.8 ;
 RECT 1.055 2.21 1.195 2.8 ;
 RECT 0.115 2.21 0.255 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.125 1.445 0.46 1.72 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.67 1.4 3.81 2.46 ;
 RECT 3.67 1.16 4.12 1.4 ;
 RECT 3.67 0.59 3.81 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END Q

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.64 0.79 2.04 1.035 ;
 RECT 1.64 1.035 1.88 1.05 ;
 END
 ANTENNAGATEAREA 0.104 ;
 END IN5

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.885 1.48 2.2 1.765 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN4

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.48 1.01 1.77 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END IN1

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 3.2 0.08 3.34 0.78 ;
 RECT 4.675 0.08 4.815 0.78 ;
 RECT 4.14 0.08 4.28 0.775 ;
 RECT 1.755 0.08 1.895 0.545 ;
 RECT 0.115 0.08 0.255 0.535 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 1.855 0.8 2.11 0.985 ;
 RECT 2.01 0.135 2.11 0.8 ;
 RECT 2.615 1.085 2.715 2.65 ;
 RECT 1.855 0.985 2.715 1.01 ;
 RECT 2.01 1.01 2.715 1.085 ;
 RECT 3.28 1.31 4.025 1.395 ;
 RECT 3.28 1.185 3.555 1.31 ;
 RECT 3.455 1.395 4.025 1.41 ;
 RECT 3.925 0.33 4.025 1.31 ;
 RECT 3.925 1.41 4.025 2.78 ;
 RECT 3.455 0.33 3.555 1.185 ;
 RECT 3.455 1.41 3.555 2.78 ;
 RECT 0.68 1.615 0.94 1.755 ;
 RECT 0.68 0.135 0.78 1.545 ;
 RECT 0.84 1.755 0.94 2.62 ;
 RECT 0.68 1.545 0.91 1.615 ;
 RECT 1.15 0.135 1.25 1.485 ;
 RECT 1.67 1.645 1.77 2.65 ;
 RECT 1.15 1.485 1.38 1.545 ;
 RECT 1.15 1.645 1.38 1.695 ;
 RECT 1.15 1.545 1.77 1.645 ;
 RECT 0.37 0.135 0.47 1.47 ;
 RECT 0.37 1.68 0.47 2.62 ;
 RECT 0.23 1.47 0.47 1.68 ;
 RECT 1.98 1.545 2.24 1.755 ;
 RECT 1.54 0.135 1.64 1.265 ;
 RECT 2.14 1.755 2.24 2.65 ;
 RECT 2.14 1.365 2.24 1.545 ;
 RECT 1.54 1.265 2.24 1.365 ;
 LAYER CO ;
 RECT 2.835 1.93 2.965 2.06 ;
 RECT 4.145 1.76 4.275 1.89 ;
 RECT 4.145 2.02 4.275 2.15 ;
 RECT 3.675 1.74 3.805 1.87 ;
 RECT 3.675 2 3.805 2.13 ;
 RECT 3.205 2 3.335 2.13 ;
 RECT 3.675 0.65 3.805 0.78 ;
 RECT 4.145 0.59 4.275 0.72 ;
 RECT 3.205 0.59 3.335 0.72 ;
 RECT 4.145 2.285 4.275 2.415 ;
 RECT 1.06 2.26 1.19 2.39 ;
 RECT 0.12 2.26 0.25 2.39 ;
 RECT 3.675 2.26 3.805 2.39 ;
 RECT 1.89 2.075 2.02 2.205 ;
 RECT 2.03 1.585 2.16 1.715 ;
 RECT 3.33 1.225 3.46 1.355 ;
 RECT 4.67 2.155 4.8 2.285 ;
 RECT 1.42 2.26 1.55 2.39 ;
 RECT 0.73 1.585 0.86 1.715 ;
 RECT 2.23 0.365 2.36 0.495 ;
 RECT 0.9 0.355 1.03 0.485 ;
 RECT 2.835 2.19 2.965 2.32 ;
 RECT 1.2 1.525 1.33 1.655 ;
 RECT 4.67 1.895 4.8 2.025 ;
 RECT 4.68 0.6 4.81 0.73 ;
 RECT 4.67 1.635 4.8 1.765 ;
 RECT 3.205 2.26 3.335 2.39 ;
 RECT 4.68 0.34 4.81 0.47 ;
 RECT 1.76 0.365 1.89 0.495 ;
 RECT 1.905 0.84 2.035 0.97 ;
 RECT 2.36 2.26 2.49 2.39 ;
 RECT 0.59 2.26 0.72 2.39 ;
 RECT 0.28 1.51 0.41 1.64 ;
 RECT 0.12 0.355 0.25 0.485 ;
 LAYER M1 ;
 RECT 2.355 2.205 2.495 2.485 ;
 RECT 1.415 2.21 1.555 2.485 ;
 RECT 1.415 2.485 2.495 2.625 ;
 RECT 0.585 2.07 0.725 2.445 ;
 RECT 1.885 2.07 2.025 2.255 ;
 RECT 0.585 1.93 2.025 2.07 ;
 RECT 2.225 0.315 2.365 1.195 ;
 RECT 0.895 1.195 2.97 1.22 ;
 RECT 2.83 1.36 2.97 2.37 ;
 RECT 0.895 0.305 1.035 1.195 ;
 RECT 3.325 1.175 3.465 1.22 ;
 RECT 3.325 1.36 3.465 1.405 ;
 RECT 0.895 1.22 3.475 1.335 ;
 RECT 2.83 1.335 3.475 1.36 ;
 END
END AO221X2

MACRO AO222X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.235 1.16 4.61 1.4 ;
 RECT 4.235 1.4 4.375 2.44 ;
 RECT 4.235 0.64 4.375 1.16 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END Q

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.48 0.475 1.72 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.48 1.08 1.79 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.48 1.72 1.77 ;
 END
 ANTENNAGATEAREA 0.083 ;
 END IN3

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.01 1.48 2.43 1.77 ;
 END
 ANTENNAGATEAREA 0.083 ;
 END IN4

 PIN IN6
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.64 0.685 1.995 1.055 ;
 END
 ANTENNAGATEAREA 0.083 ;
 END IN6

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.92 0.52 3.265 0.925 ;
 END
 ANTENNAGATEAREA 0.083 ;
 END IN5

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 3.765 0.08 3.905 0.885 ;
 RECT 4.65 0.08 4.79 0.93 ;
 RECT 0.125 0.08 0.265 0.535 ;
 RECT 1.685 0.08 1.825 0.535 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 4.65 1.645 4.79 2.8 ;
 RECT 3.765 1.95 3.905 2.8 ;
 RECT 0.125 2.235 0.265 2.8 ;
 RECT 1.065 2.215 1.205 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 2.71 1.085 2.81 2.635 ;
 RECT 1.94 0.955 2.04 0.985 ;
 RECT 1.94 0.985 2.81 1.085 ;
 RECT 1.94 0.135 2.04 0.745 ;
 RECT 1.81 0.745 2.04 0.955 ;
 RECT 1.47 0.135 1.57 1.265 ;
 RECT 2.15 1.755 2.25 2.635 ;
 RECT 2.15 1.365 2.25 1.545 ;
 RECT 1.47 1.265 2.25 1.365 ;
 RECT 2.15 1.545 2.38 1.755 ;
 RECT 1.475 1.645 1.78 1.755 ;
 RECT 1.68 1.755 1.78 2.635 ;
 RECT 1.16 0.135 1.26 1.545 ;
 RECT 1.16 1.545 1.78 1.645 ;
 RECT 0.69 1.615 0.95 1.825 ;
 RECT 0.69 0.135 0.79 1.615 ;
 RECT 0.85 1.825 0.95 2.65 ;
 RECT 0.38 0.135 0.48 1.475 ;
 RECT 0.38 1.685 0.48 2.65 ;
 RECT 0.24 1.475 0.48 1.685 ;
 RECT 4.02 0.335 4.12 1.085 ;
 RECT 4.02 1.295 4.12 2.74 ;
 RECT 3.89 1.085 4.12 1.295 ;
 RECT 3.18 0.915 3.28 2.635 ;
 RECT 2.24 0.135 2.34 0.705 ;
 RECT 3.05 0.805 3.28 0.915 ;
 RECT 2.24 0.705 3.28 0.805 ;
 LAYER CO ;
 RECT 3.94 1.125 4.07 1.255 ;
 RECT 3.77 0.705 3.9 0.835 ;
 RECT 3.77 2.26 3.9 2.39 ;
 RECT 3.77 2 3.9 2.13 ;
 RECT 4.655 0.73 4.785 0.86 ;
 RECT 4.655 0.47 4.785 0.6 ;
 RECT 4.655 1.695 4.785 1.825 ;
 RECT 4.655 2.215 4.785 2.345 ;
 RECT 4.655 1.955 4.785 2.085 ;
 RECT 1.86 0.785 1.99 0.915 ;
 RECT 2.2 1.585 2.33 1.715 ;
 RECT 1.525 1.585 1.655 1.715 ;
 RECT 0.74 1.655 0.87 1.785 ;
 RECT 0.29 1.515 0.42 1.645 ;
 RECT 3.1 0.745 3.23 0.875 ;
 RECT 2.93 2 3.06 2.13 ;
 RECT 1.9 2 2.03 2.13 ;
 RECT 4.24 2.26 4.37 2.39 ;
 RECT 4.24 2 4.37 2.13 ;
 RECT 2.46 0.355 2.59 0.485 ;
 RECT 3.4 2.26 3.53 2.39 ;
 RECT 2.37 2.26 2.5 2.39 ;
 RECT 1.43 2.26 1.56 2.39 ;
 RECT 1.69 0.355 1.82 0.485 ;
 RECT 0.91 0.355 1.04 0.485 ;
 RECT 1.07 2.29 1.2 2.42 ;
 RECT 0.6 2.115 0.73 2.245 ;
 RECT 0.13 0.355 0.26 0.485 ;
 RECT 4.24 0.705 4.37 0.835 ;
 RECT 4.24 1.74 4.37 1.87 ;
 RECT 0.13 2.295 0.26 2.425 ;
 RECT 4.24 1.48 4.37 1.61 ;
 LAYER M1 ;
 RECT 2.455 0.305 2.595 1.2 ;
 RECT 0.905 1.26 3.065 1.34 ;
 RECT 2.925 1.34 3.065 2.18 ;
 RECT 0.905 0.305 1.045 1.2 ;
 RECT 0.905 1.2 4.085 1.26 ;
 RECT 2.925 1.12 4.085 1.2 ;
 RECT 3.935 1.075 4.075 1.12 ;
 RECT 3.935 1.26 4.075 1.305 ;
 RECT 2.365 2.21 2.505 2.355 ;
 RECT 3.395 2.21 3.535 2.355 ;
 RECT 1.425 2.21 1.565 2.355 ;
 RECT 1.425 2.355 3.535 2.495 ;
 RECT 0.595 2.07 0.735 2.3 ;
 RECT 1.895 2.07 2.035 2.18 ;
 RECT 0.595 1.93 2.035 2.07 ;
 END
END AO222X1

MACRO AO222X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.92 0.52 3.37 0.925 ;
 END
 ANTENNAGATEAREA 0.083 ;
 END IN5

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 3.67 0.08 3.81 0.735 ;
 RECT 4.61 0.08 4.75 0.73 ;
 RECT 5.035 0.08 5.175 0.905 ;
 RECT 1.755 0.08 1.895 0.535 ;
 RECT 0.115 0.08 0.255 0.535 ;
 END
 END VSS

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.44 0.77 1.78 1.095 ;
 END
 ANTENNAGATEAREA 0.083 ;
 END IN4

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.14 1.16 4.44 1.4 ;
 RECT 4.14 1.4 4.28 2.46 ;
 RECT 4.14 0.64 4.28 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END Q

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.84 0.68 1.24 1.045 ;
 END
 ANTENNAGATEAREA 0.083 ;
 END IN3

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.165 1.475 0.46 1.825 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END IN2

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 5.025 1.645 5.165 2.8 ;
 RECT 3.67 1.95 3.81 2.8 ;
 RECT 4.61 1.95 4.75 2.8 ;
 RECT 0.115 2.21 0.255 2.8 ;
 RECT 1.055 2.21 1.195 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.48 1.01 1.79 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END IN1

 PIN IN6
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.925 0.815 2.205 1.095 ;
 END
 ANTENNAGATEAREA 0.083 ;
 END IN6

 OBS
 LAYER PO ;
 RECT 0.37 1.775 0.47 2.62 ;
 RECT 0.37 0.135 0.47 1.565 ;
 RECT 0.23 1.565 0.47 1.775 ;
 RECT 2.01 0.135 2.11 0.875 ;
 RECT 2.615 1.085 2.715 2.62 ;
 RECT 1.88 0.875 2.11 0.985 ;
 RECT 1.88 0.985 2.715 1.085 ;
 RECT 1.67 1.645 1.77 2.62 ;
 RECT 1.15 0.135 1.25 0.715 ;
 RECT 1.15 0.925 1.25 1.545 ;
 RECT 1.15 1.545 1.77 1.645 ;
 RECT 1.02 0.715 1.25 0.925 ;
 RECT 0.68 1.695 0.94 1.825 ;
 RECT 0.68 0.135 0.78 1.615 ;
 RECT 0.84 1.825 0.94 2.62 ;
 RECT 0.68 1.615 0.91 1.695 ;
 RECT 2.14 1.365 2.24 2.62 ;
 RECT 1.54 0.135 1.64 0.875 ;
 RECT 1.54 1.085 1.64 1.265 ;
 RECT 1.54 1.265 2.24 1.365 ;
 RECT 1.47 0.875 1.7 1.085 ;
 RECT 3.76 1.025 4.025 1.035 ;
 RECT 3.925 0.315 4.025 1.025 ;
 RECT 3.76 1.135 4.025 1.235 ;
 RECT 3.925 1.235 4.025 2.74 ;
 RECT 4.395 0.315 4.495 1.035 ;
 RECT 3.76 1.035 4.495 1.135 ;
 RECT 4.395 1.135 4.495 2.74 ;
 RECT 3.085 0.915 3.185 2.62 ;
 RECT 2.31 0.135 2.41 0.705 ;
 RECT 2.955 0.805 3.185 0.915 ;
 RECT 2.31 0.705 3.185 0.805 ;
 LAYER CO ;
 RECT 2.36 2 2.49 2.13 ;
 RECT 4.615 0.545 4.745 0.675 ;
 RECT 4.615 2.26 4.745 2.39 ;
 RECT 4.615 2 4.745 2.13 ;
 RECT 1.76 0.355 1.89 0.485 ;
 RECT 1.42 2.26 1.55 2.39 ;
 RECT 0.12 0.355 0.25 0.485 ;
 RECT 0.9 0.355 1.03 0.485 ;
 RECT 3.675 2 3.805 2.13 ;
 RECT 4.145 2.26 4.275 2.39 ;
 RECT 2.36 2.26 2.49 2.39 ;
 RECT 3.81 1.065 3.94 1.195 ;
 RECT 5.03 1.955 5.16 2.085 ;
 RECT 1.93 0.915 2.06 1.045 ;
 RECT 4.145 2 4.275 2.13 ;
 RECT 5.03 1.695 5.16 1.825 ;
 RECT 0.12 2.26 0.25 2.39 ;
 RECT 0.28 1.605 0.41 1.735 ;
 RECT 1.07 0.755 1.2 0.885 ;
 RECT 1.52 0.915 1.65 1.045 ;
 RECT 3.675 2.26 3.805 2.39 ;
 RECT 5.04 0.445 5.17 0.575 ;
 RECT 5.03 2.215 5.16 2.345 ;
 RECT 0.59 2.26 0.72 2.39 ;
 RECT 3.305 2.26 3.435 2.39 ;
 RECT 1.89 2 2.02 2.13 ;
 RECT 2.53 0.355 2.66 0.485 ;
 RECT 3.005 0.745 3.135 0.875 ;
 RECT 4.145 1.74 4.275 1.87 ;
 RECT 5.04 0.705 5.17 0.835 ;
 RECT 0.73 1.655 0.86 1.785 ;
 RECT 1.06 2.26 1.19 2.39 ;
 RECT 2.835 2 2.965 2.13 ;
 RECT 4.145 1.48 4.275 1.61 ;
 RECT 3.675 0.55 3.805 0.68 ;
 RECT 4.145 0.705 4.275 0.835 ;
 LAYER M1 ;
 RECT 2.355 1.945 2.495 2.52 ;
 RECT 3.3 2.21 3.44 2.52 ;
 RECT 1.415 2.21 1.555 2.52 ;
 RECT 1.415 2.52 3.44 2.66 ;
 RECT 2.525 0.305 2.665 1.34 ;
 RECT 1.155 1.34 3.65 1.48 ;
 RECT 3.51 1.2 3.65 1.34 ;
 RECT 2.83 1.48 2.97 2.18 ;
 RECT 0.56 0.49 0.7 1.2 ;
 RECT 0.56 0.35 1.08 0.49 ;
 RECT 0.56 1.2 1.295 1.34 ;
 RECT 3.805 1.015 3.945 1.06 ;
 RECT 3.805 1.2 3.945 1.245 ;
 RECT 3.51 1.06 3.96 1.2 ;
 RECT 0.585 2.07 0.725 2.44 ;
 RECT 1.885 2.07 2.025 2.18 ;
 RECT 0.585 1.93 2.025 2.07 ;
 END
END AO222X2

MACRO AO22X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.655 1.44 0.965 1.76 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN1

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 3.195 0.08 3.335 0.765 ;
 RECT 3.61 0.08 3.75 0.78 ;
 RECT 0.115 0.08 0.255 0.98 ;
 RECT 1.755 0.08 1.895 0.965 ;
 END
 END VSS

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.15 1.48 1.56 1.72 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN3

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 3.61 1.585 3.75 2.8 ;
 RECT 3.195 2.02 3.335 2.8 ;
 RECT 1.055 2.21 1.195 2.8 ;
 RECT 0.115 2.21 0.255 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.44 0.475 1.76 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.725 1.16 3 1.4 ;
 RECT 2.725 1.4 2.865 2.44 ;
 RECT 2.725 0.685 2.865 1.16 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END Q

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.88 1.48 2.205 1.765 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN4

 OBS
 LAYER PO ;
 RECT 2.98 1.085 3.08 2.74 ;
 RECT 2.98 0.315 3.08 0.985 ;
 RECT 2.31 0.875 2.54 0.985 ;
 RECT 2.31 0.985 3.08 1.085 ;
 RECT 1.98 1.545 2.24 1.755 ;
 RECT 1.54 0.565 1.64 1.265 ;
 RECT 2.14 1.755 2.24 2.62 ;
 RECT 2.14 1.365 2.24 1.545 ;
 RECT 1.54 1.265 2.24 1.365 ;
 RECT 0.68 0.565 0.78 1.545 ;
 RECT 0.84 1.795 0.94 2.62 ;
 RECT 0.68 1.545 0.91 1.695 ;
 RECT 0.68 1.695 0.94 1.795 ;
 RECT 1.15 0.565 1.25 1.475 ;
 RECT 1.67 1.645 1.77 2.62 ;
 RECT 1.15 1.475 1.38 1.545 ;
 RECT 1.15 1.645 1.38 1.695 ;
 RECT 1.15 1.545 1.77 1.645 ;
 RECT 0.37 1.71 0.47 2.62 ;
 RECT 0.37 0.565 0.47 1.5 ;
 RECT 0.23 1.5 0.47 1.71 ;
 LAYER CO ;
 RECT 3.2 2.08 3.33 2.21 ;
 RECT 2.73 1.74 2.86 1.87 ;
 RECT 2.73 2 2.86 2.13 ;
 RECT 1.76 0.785 1.89 0.915 ;
 RECT 1.89 2.08 2.02 2.21 ;
 RECT 2.03 1.585 2.16 1.715 ;
 RECT 2.36 0.915 2.49 1.045 ;
 RECT 0.73 1.585 0.86 1.715 ;
 RECT 3.615 2.155 3.745 2.285 ;
 RECT 3.615 1.895 3.745 2.025 ;
 RECT 1.2 1.525 1.33 1.655 ;
 RECT 3.2 0.555 3.33 0.685 ;
 RECT 0.59 2.08 0.72 2.21 ;
 RECT 0.28 1.54 0.41 1.67 ;
 RECT 3.615 1.635 3.745 1.765 ;
 RECT 0.12 0.785 0.25 0.915 ;
 RECT 3.615 0.6 3.745 0.73 ;
 RECT 1.06 2.26 1.19 2.39 ;
 RECT 0.9 0.785 1.03 0.915 ;
 RECT 3.2 2.34 3.33 2.47 ;
 RECT 3.615 0.34 3.745 0.47 ;
 RECT 2.73 2.26 2.86 2.39 ;
 RECT 2.73 0.735 2.86 0.865 ;
 RECT 1.42 2.26 1.55 2.39 ;
 RECT 2.36 2.26 2.49 2.39 ;
 RECT 0.12 2.26 0.25 2.39 ;
 LAYER M1 ;
 RECT 0.585 2.07 0.725 2.265 ;
 RECT 1.885 2.07 2.025 2.26 ;
 RECT 0.585 1.93 2.025 2.07 ;
 RECT 0.895 0.735 1.035 1.14 ;
 RECT 1.415 2.21 1.555 2.485 ;
 RECT 2.355 0.865 2.495 1.14 ;
 RECT 2.355 1.28 2.495 2.485 ;
 RECT 0.895 1.14 2.495 1.28 ;
 RECT 1.415 2.485 2.495 2.625 ;
 END
END AO22X1

MACRO AO22X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.195 1.475 1.56 1.72 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN3

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.88 1.48 2.2 1.765 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN4

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.56 0.965 3.805 1.13 ;
 RECT 3.665 0.455 3.805 0.825 ;
 RECT 3.665 1.13 3.805 2.44 ;
 RECT 2.725 0.965 2.865 2.44 ;
 RECT 2.725 0.825 3.805 0.965 ;
 RECT 2.725 0.455 2.865 0.825 ;
 END
 ANTENNADIFFAREA 0.93 ;
 END Q

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.47 0.94 1.755 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.48 0.47 1.72 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 3.195 0.08 3.335 0.65 ;
 RECT 4.08 0.08 4.22 0.78 ;
 RECT 0.115 0.08 0.255 0.8 ;
 RECT 1.755 0.08 1.895 0.795 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 3.195 1.68 3.335 2.8 ;
 RECT 4.08 1.585 4.22 2.8 ;
 RECT 0.115 2.21 0.255 2.8 ;
 RECT 1.055 2.21 1.195 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 1.98 1.545 2.24 1.755 ;
 RECT 1.54 0.395 1.64 1.265 ;
 RECT 2.14 1.755 2.24 2.62 ;
 RECT 2.14 1.365 2.24 1.545 ;
 RECT 1.54 1.265 2.24 1.365 ;
 RECT 0.37 0.395 0.47 1.48 ;
 RECT 0.37 1.72 0.47 2.62 ;
 RECT 0.23 1.48 0.47 1.72 ;
 RECT 3.45 1.085 3.55 2.74 ;
 RECT 2.98 1.085 3.08 2.74 ;
 RECT 2.31 0.985 3.55 1.085 ;
 RECT 3.45 0.205 3.55 0.985 ;
 RECT 2.98 0.205 3.08 0.985 ;
 RECT 2.31 0.875 2.54 0.985 ;
 RECT 0.68 0.395 0.78 1.545 ;
 RECT 0.84 1.795 0.94 2.62 ;
 RECT 0.68 1.545 0.91 1.695 ;
 RECT 0.68 1.695 0.94 1.795 ;
 RECT 1.15 0.395 1.25 1.485 ;
 RECT 1.67 1.645 1.77 2.62 ;
 RECT 1.15 1.485 1.38 1.545 ;
 RECT 1.15 1.645 1.38 1.695 ;
 RECT 1.15 1.545 1.77 1.645 ;
 LAYER CO ;
 RECT 3.67 1.74 3.8 1.87 ;
 RECT 2.73 1.74 2.86 1.87 ;
 RECT 3.2 1.74 3.33 1.87 ;
 RECT 3.2 2 3.33 2.13 ;
 RECT 3.67 2 3.8 2.13 ;
 RECT 2.73 2 2.86 2.13 ;
 RECT 3.67 0.515 3.8 0.645 ;
 RECT 3.67 2.26 3.8 2.39 ;
 RECT 1.06 2.26 1.19 2.39 ;
 RECT 3.2 0.46 3.33 0.59 ;
 RECT 1.2 1.525 1.33 1.655 ;
 RECT 2.73 2.26 2.86 2.39 ;
 RECT 4.085 2.155 4.215 2.285 ;
 RECT 0.12 2.26 0.25 2.39 ;
 RECT 2.36 2.26 2.49 2.39 ;
 RECT 1.76 0.615 1.89 0.745 ;
 RECT 4.085 1.895 4.215 2.025 ;
 RECT 2.03 1.585 2.16 1.715 ;
 RECT 1.89 2.08 2.02 2.21 ;
 RECT 0.12 0.615 0.25 0.745 ;
 RECT 4.085 0.6 4.215 0.73 ;
 RECT 4.085 1.635 4.215 1.765 ;
 RECT 4.085 0.34 4.215 0.47 ;
 RECT 0.59 2.26 0.72 2.39 ;
 RECT 3.2 2.26 3.33 2.39 ;
 RECT 1.42 2.26 1.55 2.39 ;
 RECT 0.9 0.615 1.03 0.745 ;
 RECT 0.285 1.54 0.415 1.67 ;
 RECT 2.36 0.915 2.49 1.045 ;
 RECT 2.73 0.515 2.86 0.645 ;
 RECT 0.73 1.585 0.86 1.715 ;
 LAYER M1 ;
 RECT 0.585 2.07 0.725 2.445 ;
 RECT 1.885 2.07 2.025 2.26 ;
 RECT 0.585 1.93 2.025 2.07 ;
 RECT 0.895 0.56 1.035 1.04 ;
 RECT 1.415 2.21 1.555 2.485 ;
 RECT 2.355 0.865 2.495 1.04 ;
 RECT 2.355 1.18 2.495 2.485 ;
 RECT 1.415 2.485 2.495 2.625 ;
 RECT 0.895 1.04 2.495 1.18 ;
 END
END AO22X2

MACRO AOI21X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 3.625 1.585 3.765 2.8 ;
 RECT 2.735 2.05 2.875 2.8 ;
 RECT 0.115 2.21 0.255 2.8 ;
 RECT 1.055 2.21 1.195 2.8 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.205 1.4 3.345 2.44 ;
 RECT 3.205 1.16 3.48 1.4 ;
 RECT 3.205 0.495 3.345 1.16 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END QN

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.63 1.46 0.92 1.72 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.445 0.47 1.72 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN2

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.185 1.475 1.56 1.72 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 2.735 0.08 2.875 0.735 ;
 RECT 3.62 0.08 3.76 0.78 ;
 RECT 1.365 0.08 1.505 0.965 ;
 RECT 0.115 0.08 0.255 0.965 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 2.52 0.55 2.62 2.1 ;
 RECT 2.39 2.1 2.62 2.31 ;
 RECT 0.68 1.545 0.92 1.695 ;
 RECT 0.68 0.565 0.78 1.545 ;
 RECT 0.84 1.795 0.94 2.62 ;
 RECT 0.68 1.695 0.94 1.795 ;
 RECT 0.37 0.565 0.47 1.5 ;
 RECT 0.37 1.71 0.47 2.62 ;
 RECT 0.24 1.5 0.47 1.71 ;
 RECT 2.99 1.38 3.09 2.76 ;
 RECT 2.99 0.33 3.09 1.17 ;
 RECT 2.81 1.17 3.09 1.38 ;
 RECT 1.15 1.485 1.39 1.545 ;
 RECT 1.15 0.565 1.25 1.485 ;
 RECT 1.68 1.645 1.78 2.62 ;
 RECT 1.16 1.645 1.39 1.695 ;
 RECT 1.15 1.545 1.78 1.645 ;
 LAYER CO ;
 RECT 3.21 1.74 3.34 1.87 ;
 RECT 3.21 2 3.34 2.13 ;
 RECT 2.74 2.11 2.87 2.24 ;
 RECT 0.29 1.54 0.42 1.67 ;
 RECT 1.37 0.785 1.5 0.915 ;
 RECT 1.9 2.27 2.03 2.4 ;
 RECT 3.63 2.155 3.76 2.285 ;
 RECT 1.43 2.27 1.56 2.4 ;
 RECT 0.12 2.26 0.25 2.39 ;
 RECT 3.21 2.26 3.34 2.39 ;
 RECT 3.63 1.635 3.76 1.765 ;
 RECT 3.21 0.55 3.34 0.68 ;
 RECT 3.625 0.6 3.755 0.73 ;
 RECT 1.21 1.525 1.34 1.655 ;
 RECT 0.12 0.785 0.25 0.915 ;
 RECT 0.9 0.785 1.03 0.915 ;
 RECT 3.625 0.34 3.755 0.47 ;
 RECT 2.27 0.77 2.4 0.9 ;
 RECT 3.63 1.895 3.76 2.025 ;
 RECT 2.74 2.37 2.87 2.5 ;
 RECT 2.74 0.55 2.87 0.68 ;
 RECT 2.27 1.59 2.4 1.72 ;
 RECT 1.06 2.26 1.19 2.39 ;
 RECT 0.74 1.585 0.87 1.715 ;
 RECT 2.86 1.21 2.99 1.34 ;
 RECT 0.59 2.26 0.72 2.39 ;
 RECT 2.44 2.14 2.57 2.27 ;
 LAYER M1 ;
 RECT 0.585 2.07 0.725 2.445 ;
 RECT 1.425 2.07 1.565 2.46 ;
 RECT 0.585 1.93 1.565 2.07 ;
 RECT 0.895 0.735 1.035 1.165 ;
 RECT 1.895 1.305 2.035 2.14 ;
 RECT 1.895 2.14 2.59 2.28 ;
 RECT 1.895 2.28 2.035 2.455 ;
 RECT 2.435 2.09 2.575 2.14 ;
 RECT 2.435 2.28 2.575 2.32 ;
 RECT 0.895 1.165 2.035 1.305 ;
 RECT 2.265 0.715 2.405 1.205 ;
 RECT 2.265 1.345 2.405 1.77 ;
 RECT 2.855 1.16 2.995 1.205 ;
 RECT 2.855 1.345 2.995 1.39 ;
 RECT 2.265 1.205 2.995 1.345 ;
 END
END AOI21X1

MACRO AOI21X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 4.09 0.08 4.23 0.78 ;
 RECT 2.735 0.08 2.875 0.925 ;
 RECT 3.675 0.08 3.815 0.875 ;
 RECT 0.115 0.08 0.255 0.805 ;
 RECT 1.365 0.08 1.505 0.795 ;
 END
 END VSS

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.745 2.115 2.2 2.415 ;
 END
 ANTENNAGATEAREA 0.086 ;
 END IN3

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.16 0.475 1.4 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.64 1.465 0.96 1.72 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 4.09 1.585 4.23 2.8 ;
 RECT 2.735 2.055 2.875 2.8 ;
 RECT 3.675 2.035 3.815 2.8 ;
 RECT 0.115 2.21 0.255 2.8 ;
 RECT 1.055 2.21 1.195 2.8 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.205 1.4 3.345 2.44 ;
 RECT 3.205 1.155 3.48 1.4 ;
 RECT 3.205 0.63 3.345 1.155 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END QN

 OBS
 LAYER PO ;
 RECT 2.52 0.525 2.62 0.985 ;
 RECT 2.52 1.085 2.62 2.195 ;
 RECT 1.85 0.875 2.08 0.985 ;
 RECT 1.85 0.985 2.62 1.085 ;
 RECT 0.68 1.545 0.92 1.695 ;
 RECT 0.68 0.395 0.78 1.545 ;
 RECT 0.84 1.795 0.94 2.62 ;
 RECT 0.68 1.695 0.94 1.795 ;
 RECT 1.15 0.395 1.25 1.27 ;
 RECT 1.68 1.37 1.78 2.23 ;
 RECT 1.68 2.23 1.98 2.46 ;
 RECT 1.15 1.27 1.78 1.37 ;
 RECT 0.37 1.39 0.47 2.62 ;
 RECT 0.37 0.395 0.47 1.16 ;
 RECT 0.255 1.16 0.47 1.39 ;
 RECT 3.46 1.35 3.56 2.76 ;
 RECT 2.99 1.38 3.09 2.76 ;
 RECT 2.99 0.305 3.09 1.17 ;
 RECT 2.81 1.17 3.09 1.25 ;
 RECT 2.81 1.25 3.56 1.35 ;
 RECT 2.81 1.35 3.09 1.38 ;
 RECT 3.46 0.305 3.56 1.25 ;
 LAYER CO ;
 RECT 2.27 1.77 2.4 1.9 ;
 RECT 3.21 1.74 3.34 1.87 ;
 RECT 2.74 2.11 2.87 2.24 ;
 RECT 3.68 2.11 3.81 2.24 ;
 RECT 3.21 2 3.34 2.13 ;
 RECT 3.68 0.685 3.81 0.815 ;
 RECT 3.68 2.37 3.81 2.5 ;
 RECT 2.74 0.73 2.87 0.86 ;
 RECT 3.21 0.69 3.34 0.82 ;
 RECT 2.27 0.745 2.4 0.875 ;
 RECT 2.27 1.51 2.4 1.64 ;
 RECT 0.74 1.585 0.87 1.715 ;
 RECT 4.095 2.155 4.225 2.285 ;
 RECT 0.295 1.21 0.425 1.34 ;
 RECT 0.12 2.26 0.25 2.39 ;
 RECT 4.095 1.895 4.225 2.025 ;
 RECT 0.59 2.26 0.72 2.39 ;
 RECT 0.9 0.615 1.03 0.745 ;
 RECT 3.21 2.26 3.34 2.39 ;
 RECT 1.43 1.58 1.56 1.71 ;
 RECT 4.095 1.635 4.225 1.765 ;
 RECT 2.74 2.37 2.87 2.5 ;
 RECT 1.06 2.26 1.19 2.39 ;
 RECT 2.86 1.21 2.99 1.34 ;
 RECT 4.095 0.34 4.225 0.47 ;
 RECT 0.12 0.615 0.25 0.745 ;
 RECT 1.81 2.28 1.94 2.41 ;
 RECT 1.9 0.915 2.03 1.045 ;
 RECT 1.37 0.615 1.5 0.745 ;
 RECT 4.095 0.6 4.225 0.73 ;
 RECT 1.9 1.575 2.03 1.705 ;
 LAYER M1 ;
 RECT 0.585 2.07 0.725 2.445 ;
 RECT 1.425 1.515 1.565 1.93 ;
 RECT 0.585 1.93 1.565 2.07 ;
 RECT 2.265 0.685 2.405 1.205 ;
 RECT 2.265 1.345 2.405 1.955 ;
 RECT 2.855 1.16 2.995 1.205 ;
 RECT 2.855 1.345 2.995 1.39 ;
 RECT 2.265 1.205 2.995 1.345 ;
 RECT 0.895 0.545 1.035 0.94 ;
 RECT 1.71 0.865 2.035 0.94 ;
 RECT 1.71 1.08 2.035 1.11 ;
 RECT 1.895 1.11 2.035 1.76 ;
 RECT 0.895 0.94 2.035 1.08 ;
 END
END AOI21X2

MACRO AOI221X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.96 1.28 2.2 1.72 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN4

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.48 0.46 1.825 ;
 END
 ANTENNAGATEAREA 0.065 ;
 END IN2

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.195 1.475 1.56 1.72 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN3

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.57 0.22 0.93 0.475 ;
 END
 ANTENNAGATEAREA 0.065 ;
 END IN1

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 3.695 0.08 3.835 0.685 ;
 RECT 4.64 0.08 4.78 0.855 ;
 RECT 0.115 0.08 0.255 0.855 ;
 RECT 1.755 0.08 1.895 0.855 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 4.58 1.585 4.72 2.8 ;
 RECT 3.695 1.89 3.835 2.8 ;
 RECT 1.055 2.21 1.195 2.8 ;
 RECT 0.115 2.21 0.255 2.8 ;
 END
 END VDD

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.05 0.225 2.525 0.48 ;
 END
 ANTENNAGATEAREA 0.116 ;
 END IN5

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.165 1.08 4.305 2.44 ;
 RECT 4.165 0.84 4.44 1.08 ;
 RECT 4.165 0.41 4.305 0.84 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END QN

 OBS
 LAYER PO ;
 RECT 3.48 0.255 3.58 1.285 ;
 RECT 2.9 1.285 3.58 1.385 ;
 RECT 3.48 1.385 3.58 2.39 ;
 RECT 2.9 1.255 3.13 1.285 ;
 RECT 2.9 1.385 3.13 1.465 ;
 RECT 1.54 0.45 1.64 1.265 ;
 RECT 2.14 1.505 2.24 2.62 ;
 RECT 1.98 1.365 2.24 1.505 ;
 RECT 1.54 1.265 2.24 1.365 ;
 RECT 1.15 0.45 1.25 1.485 ;
 RECT 1.67 1.645 1.77 2.62 ;
 RECT 1.15 1.485 1.38 1.545 ;
 RECT 1.15 1.645 1.38 1.695 ;
 RECT 1.15 1.545 1.77 1.645 ;
 RECT 0.23 1.65 0.47 1.86 ;
 RECT 0.37 0.45 0.47 1.65 ;
 RECT 0.37 1.86 0.47 2.62 ;
 RECT 2.615 1.085 2.715 2.77 ;
 RECT 2.01 0.455 2.11 0.985 ;
 RECT 2.01 0.985 2.715 1.085 ;
 RECT 2.005 0.245 2.235 0.455 ;
 RECT 0.84 1.795 0.94 2.62 ;
 RECT 0.68 0.475 0.78 1.695 ;
 RECT 0.68 1.695 0.94 1.795 ;
 RECT 0.68 0.265 0.91 0.475 ;
 RECT 3.95 1.18 4.05 2.74 ;
 RECT 3.95 0.255 4.05 0.97 ;
 RECT 3.835 0.97 4.065 1.18 ;
 LAYER CO ;
 RECT 4.645 0.395 4.775 0.525 ;
 RECT 2.95 1.295 3.08 1.425 ;
 RECT 3.23 2.03 3.36 2.16 ;
 RECT 1.2 1.525 1.33 1.655 ;
 RECT 1.06 2.26 1.19 2.39 ;
 RECT 2.36 2.205 2.49 2.335 ;
 RECT 3.7 0.475 3.83 0.605 ;
 RECT 0.9 0.67 1.03 0.8 ;
 RECT 0.12 0.67 0.25 0.8 ;
 RECT 0.28 1.69 0.41 1.82 ;
 RECT 4.585 2.155 4.715 2.285 ;
 RECT 3.23 0.475 3.36 0.605 ;
 RECT 3.7 1.97 3.83 2.1 ;
 RECT 1.76 0.67 1.89 0.8 ;
 RECT 4.17 2.26 4.3 2.39 ;
 RECT 2.03 1.335 2.16 1.465 ;
 RECT 4.585 1.635 4.715 1.765 ;
 RECT 0.59 2.26 0.72 2.39 ;
 RECT 0.12 2.26 0.25 2.39 ;
 RECT 1.89 2.075 2.02 2.205 ;
 RECT 1.42 2.26 1.55 2.39 ;
 RECT 2.835 2.19 2.965 2.32 ;
 RECT 2.055 0.285 2.185 0.415 ;
 RECT 4.645 0.655 4.775 0.785 ;
 RECT 3.885 1.01 4.015 1.14 ;
 RECT 4.17 2 4.3 2.13 ;
 RECT 2.23 0.67 2.36 0.8 ;
 RECT 4.585 1.895 4.715 2.025 ;
 RECT 0.73 0.305 0.86 0.435 ;
 RECT 4.17 0.475 4.3 0.605 ;
 LAYER M1 ;
 RECT 0.585 2.07 0.725 2.445 ;
 RECT 1.885 2.07 2.025 2.255 ;
 RECT 0.585 1.93 2.025 2.07 ;
 RECT 2.355 2.145 2.495 2.485 ;
 RECT 1.415 2.21 1.555 2.485 ;
 RECT 1.415 2.485 2.495 2.625 ;
 RECT 3.225 0.42 3.365 1.005 ;
 RECT 3.225 1.145 3.365 2.23 ;
 RECT 3.225 1.005 4.02 1.145 ;
 RECT 3.88 0.96 4.02 1.005 ;
 RECT 3.88 1.145 4.02 1.19 ;
 RECT 0.895 0.62 1.035 0.995 ;
 RECT 2.225 0.62 2.365 0.995 ;
 RECT 2.83 1.135 2.97 1.245 ;
 RECT 2.83 1.475 2.97 2.37 ;
 RECT 0.895 0.995 2.97 1.135 ;
 RECT 2.83 1.245 3.085 1.475 ;
 END
END AOI221X1

MACRO AOI221X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.76 1.16 2.255 1.515 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN4

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.63 0.34 3.055 0.665 ;
 END
 ANTENNAGATEAREA 0.116 ;
 END IN5

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.455 0.47 1.73 ;
 END
 ANTENNAGATEAREA 0.065 ;
 END IN2

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.12 1.16 1.51 1.44 ;
 END
 ANTENNAGATEAREA 0.068 ;
 END IN3

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.51 2.245 0.915 2.66 ;
 END
 ANTENNAGATEAREA 0.065 ;
 END IN1

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 3.695 0.08 3.835 0.96 ;
 RECT 4.635 0.08 4.775 0.775 ;
 RECT 5.05 0.08 5.19 0.88 ;
 RECT 1.755 0.08 1.895 0.695 ;
 RECT 0.115 0.08 0.255 0.71 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 3.695 2.06 3.835 2.8 ;
 RECT 5.05 1.585 5.19 2.8 ;
 RECT 4.635 2.055 4.775 2.8 ;
 RECT 0.115 2.09 0.255 2.8 ;
 RECT 1.055 2.095 1.195 2.8 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.165 1.425 4.305 2.44 ;
 RECT 4.165 1.16 4.6 1.425 ;
 RECT 4.165 0.59 4.305 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END QN

 OBS
 LAYER PO ;
 RECT 1.54 0.295 1.64 1.265 ;
 RECT 2.155 1.505 2.255 2.385 ;
 RECT 1.965 1.365 2.255 1.505 ;
 RECT 1.54 1.265 2.255 1.365 ;
 RECT 3.48 0.555 3.58 2.025 ;
 RECT 3.33 2.025 3.58 2.235 ;
 RECT 0.37 0.295 0.47 1.49 ;
 RECT 0.37 1.7 0.47 2.505 ;
 RECT 0.23 1.49 0.47 1.7 ;
 RECT 2.01 0.295 2.11 0.985 ;
 RECT 2.63 0.655 2.73 0.985 ;
 RECT 2.63 1.085 2.73 2.78 ;
 RECT 2.01 0.985 2.73 1.085 ;
 RECT 2.63 0.435 2.975 0.655 ;
 RECT 0.68 0.295 0.78 1.695 ;
 RECT 0.84 1.795 0.94 2.405 ;
 RECT 0.66 2.405 0.94 2.615 ;
 RECT 0.68 1.695 0.94 1.795 ;
 RECT 1.15 0.295 1.25 1.155 ;
 RECT 1.685 1.645 1.785 2.385 ;
 RECT 1.15 1.365 1.25 1.545 ;
 RECT 1.15 1.545 1.785 1.645 ;
 RECT 1.12 1.155 1.35 1.365 ;
 RECT 3.825 1.135 4.52 1.18 ;
 RECT 4.42 1.18 4.52 2.74 ;
 RECT 4.42 0.335 4.52 1.08 ;
 RECT 3.875 1.08 4.52 1.135 ;
 RECT 3.95 0.335 4.05 1.08 ;
 RECT 3.95 1.345 4.05 2.74 ;
 RECT 3.825 1.18 4.055 1.345 ;
 LAYER CO ;
 RECT 2.85 1.93 2.98 2.06 ;
 RECT 4.17 1.74 4.3 1.87 ;
 RECT 3.7 2.11 3.83 2.24 ;
 RECT 4.64 2.11 4.77 2.24 ;
 RECT 4.64 0.585 4.77 0.715 ;
 RECT 4.64 2.37 4.77 2.5 ;
 RECT 3.23 0.775 3.36 0.905 ;
 RECT 1.06 2.145 1.19 2.275 ;
 RECT 0.12 2.145 0.25 2.275 ;
 RECT 5.055 0.42 5.185 0.55 ;
 RECT 1.17 1.195 1.3 1.325 ;
 RECT 5.055 0.68 5.185 0.81 ;
 RECT 3.875 1.175 4.005 1.305 ;
 RECT 0.12 0.515 0.25 0.645 ;
 RECT 0.71 2.445 0.84 2.575 ;
 RECT 2.375 2.01 2.505 2.14 ;
 RECT 0.9 0.515 1.03 0.645 ;
 RECT 5.055 1.635 5.185 1.765 ;
 RECT 2.85 2.19 2.98 2.32 ;
 RECT 2.795 0.485 2.925 0.615 ;
 RECT 5.055 2.155 5.185 2.285 ;
 RECT 1.905 1.775 2.035 1.905 ;
 RECT 1.435 2.03 1.565 2.16 ;
 RECT 5.055 1.895 5.185 2.025 ;
 RECT 4.17 2.26 4.3 2.39 ;
 RECT 3.7 2.37 3.83 2.5 ;
 RECT 0.59 1.93 0.72 2.06 ;
 RECT 0.28 1.53 0.41 1.66 ;
 RECT 1.76 0.515 1.89 0.645 ;
 RECT 2.015 1.335 2.145 1.465 ;
 RECT 4.17 2 4.3 2.13 ;
 RECT 4.17 0.665 4.3 0.795 ;
 RECT 3.38 2.065 3.51 2.195 ;
 RECT 3.7 0.775 3.83 0.905 ;
 RECT 2.23 0.525 2.36 0.655 ;
 RECT 3.23 1.52 3.36 1.65 ;
 LAYER M1 ;
 RECT 2.37 1.945 2.51 2.25 ;
 RECT 1.43 1.96 1.57 2.25 ;
 RECT 1.43 2.25 2.51 2.39 ;
 RECT 0.75 1.8 0.89 1.925 ;
 RECT 0.75 1.77 2.085 1.8 ;
 RECT 0.75 1.66 2.04 1.77 ;
 RECT 1.855 1.8 2.085 1.91 ;
 RECT 0.515 1.925 0.89 2.065 ;
 RECT 0.895 0.465 1.035 0.87 ;
 RECT 2.225 0.475 2.365 0.87 ;
 RECT 2.845 1.01 2.985 2.06 ;
 RECT 2.845 2.06 3.53 2.2 ;
 RECT 2.845 2.2 2.985 2.37 ;
 RECT 3.375 2.015 3.515 2.06 ;
 RECT 3.375 2.2 3.515 2.245 ;
 RECT 0.895 0.87 2.985 1.01 ;
 RECT 3.225 0.72 3.365 1.17 ;
 RECT 3.225 1.31 3.365 1.7 ;
 RECT 3.87 1.125 4.01 1.17 ;
 RECT 3.87 1.31 4.01 1.355 ;
 RECT 3.225 1.17 4.025 1.31 ;
 END
END AOI221X2

MACRO AOI222X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 0.84 0.475 1.22 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 4.14 0.08 4.28 0.74 ;
 RECT 5.025 0.08 5.165 0.785 ;
 RECT 2.53 0.08 2.67 0.65 ;
 RECT 0.94 0.08 1.08 0.555 ;
 END
 END VSS

 PIN IN6
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.52 2.275 2.9 2.66 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN6

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 4.14 2.205 4.28 2.8 ;
 RECT 5.025 1.585 5.165 2.8 ;
 RECT 0.115 1.71 0.255 2.8 ;
 RECT 1.055 1.76 1.195 2.8 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.565 1.16 4.95 1.405 ;
 RECT 4.61 1.405 4.75 2.215 ;
 RECT 4.61 0.665 4.75 1.16 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END QN

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2 2.27 2.38 2.66 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN4

 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.11 1.13 3.5 1.455 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN5

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.375 2.27 1.785 2.66 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN3

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.485 2.12 0.915 2.41 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 3.085 0.245 3.185 1.15 ;
 RECT 3.085 1.38 3.185 2.395 ;
 RECT 3.085 1.15 3.375 1.38 ;
 RECT 1.975 0.245 2.075 1.19 ;
 RECT 1.67 1.29 1.77 2.29 ;
 RECT 1.67 1.19 2.075 1.29 ;
 RECT 1.56 2.29 1.77 2.52 ;
 RECT 0.37 1.22 0.47 2.16 ;
 RECT 1.195 0.15 1.295 0.62 ;
 RECT 0.37 0.72 0.47 1.01 ;
 RECT 0.23 1.01 0.47 1.22 ;
 RECT 0.37 0.62 1.295 0.72 ;
 RECT 2.315 0.245 2.415 1.47 ;
 RECT 2.14 1.57 2.24 2.27 ;
 RECT 2.14 1.47 2.415 1.57 ;
 RECT 2.14 2.27 2.35 2.5 ;
 RECT 2.785 0.245 2.885 1.39 ;
 RECT 2.615 1.49 2.715 2.3 ;
 RECT 2.615 1.39 2.885 1.49 ;
 RECT 2.615 2.3 2.825 2.53 ;
 RECT 1.505 0.245 1.605 0.9 ;
 RECT 0.84 1 0.94 2.105 ;
 RECT 0.68 2.105 0.94 2.315 ;
 RECT 0.84 0.9 1.605 1 ;
 RECT 4.395 0.33 4.495 1.09 ;
 RECT 4.395 1.3 4.495 2.74 ;
 RECT 4.24 1.09 4.495 1.3 ;
 RECT 3.925 0.61 4.025 2.12 ;
 RECT 3.765 0.4 4.025 0.61 ;
 LAYER CO ;
 RECT 3.205 1.2 3.335 1.33 ;
 RECT 4.615 1.505 4.745 1.635 ;
 RECT 1.6 2.34 1.73 2.47 ;
 RECT 5.03 0.34 5.16 0.47 ;
 RECT 4.29 1.13 4.42 1.26 ;
 RECT 2.655 2.35 2.785 2.48 ;
 RECT 0.12 1.77 0.25 1.9 ;
 RECT 3.675 0.77 3.805 0.9 ;
 RECT 4.145 0.555 4.275 0.685 ;
 RECT 5.03 2.155 5.16 2.285 ;
 RECT 5.03 1.635 5.16 1.765 ;
 RECT 4.615 0.72 4.745 0.85 ;
 RECT 3.675 1.515 3.805 1.645 ;
 RECT 4.615 2.025 4.745 2.155 ;
 RECT 5.03 1.895 5.16 2.025 ;
 RECT 0.73 2.145 0.86 2.275 ;
 RECT 1.89 1.71 2.02 1.84 ;
 RECT 1.42 1.82 1.55 1.95 ;
 RECT 2.36 1.82 2.49 1.95 ;
 RECT 1.06 1.81 1.19 1.94 ;
 RECT 2.835 1.695 2.965 1.825 ;
 RECT 4.145 2.26 4.275 2.39 ;
 RECT 3.815 0.44 3.945 0.57 ;
 RECT 5.03 0.6 5.16 0.73 ;
 RECT 0.945 0.37 1.075 0.5 ;
 RECT 1.725 0.465 1.855 0.595 ;
 RECT 4.615 1.765 4.745 1.895 ;
 RECT 3.305 0.465 3.435 0.595 ;
 RECT 0.28 1.05 0.41 1.18 ;
 RECT 3.305 1.82 3.435 1.95 ;
 RECT 2.535 0.465 2.665 0.595 ;
 RECT 0.59 1.635 0.72 1.765 ;
 RECT 2.18 2.32 2.31 2.45 ;
 LAYER M1 ;
 RECT 1.72 0.41 1.86 0.79 ;
 RECT 2.83 0.93 2.97 1.69 ;
 RECT 2.83 1.83 2.97 1.835 ;
 RECT 2.775 1.69 3.015 1.83 ;
 RECT 3.3 0.555 3.44 0.79 ;
 RECT 3.3 0.435 4 0.555 ;
 RECT 3.76 0.555 4 0.575 ;
 RECT 3.3 0.415 3.99 0.435 ;
 RECT 1.72 0.79 3.44 0.93 ;
 RECT 3.67 0.715 3.81 1.1 ;
 RECT 3.67 1.24 3.81 1.695 ;
 RECT 4.285 1.08 4.425 1.1 ;
 RECT 4.285 1.24 4.425 1.31 ;
 RECT 3.67 1.1 4.425 1.24 ;
 RECT 2.355 1.77 2.495 1.99 ;
 RECT 3.3 1.68 3.44 1.99 ;
 RECT 1.415 1.68 1.555 1.99 ;
 RECT 1.415 1.99 3.44 2.13 ;
 RECT 0.585 1.535 0.725 1.845 ;
 RECT 1.885 1.535 2.025 1.705 ;
 RECT 1.84 1.705 2.07 1.845 ;
 RECT 0.585 1.395 2.025 1.535 ;
 END
END AOI222X1

MACRO AOI222X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.08 BY 2.88 ;
 PIN IN5
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.915 0.54 3.165 0.925 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN5

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.835 0.585 1.26 0.915 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN3

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.48 0.46 1.77 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.64 1.36 0.98 1.745 ;
 END
 ANTENNAGATEAREA 0.061 ;
 END IN1

 PIN IN6
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.88 0.585 2.205 0.92 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN6

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.08 0.08 ;
 RECT 1.71 0.305 1.94 0.445 ;
 RECT 4.14 0.08 4.28 0.9 ;
 RECT 5.08 0.08 5.22 0.695 ;
 RECT 5.57 0.08 5.71 0.93 ;
 RECT 0.115 0.08 0.255 0.49 ;
 RECT 1.755 0.08 1.895 0.305 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.08 2.96 ;
 RECT 5.495 1.585 5.635 2.8 ;
 RECT 4.14 2.065 4.28 2.8 ;
 RECT 5.08 2.065 5.22 2.8 ;
 RECT 1.055 2.195 1.195 2.8 ;
 RECT 0.115 2.17 0.255 2.8 ;
 END
 END VDD

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.415 0.585 1.73 0.93 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END IN4

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.61 1.14 4.945 1.415 ;
 RECT 4.61 1.415 4.75 2.44 ;
 RECT 4.61 0.605 4.75 1.14 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END QN

 OBS
 LAYER PO ;
 RECT 2.14 1.415 2.24 2.625 ;
 RECT 1.54 0.09 1.64 0.585 ;
 RECT 1.54 0.795 1.64 1.315 ;
 RECT 1.54 1.315 2.24 1.415 ;
 RECT 1.43 0.585 1.675 0.795 ;
 RECT 0.37 0.09 0.47 1.545 ;
 RECT 0.37 1.755 0.47 2.62 ;
 RECT 0.23 1.545 0.47 1.755 ;
 RECT 1.67 1.695 1.77 2.625 ;
 RECT 1.15 0.09 1.25 0.595 ;
 RECT 1.15 0.805 1.25 1.595 ;
 RECT 1.15 1.595 1.77 1.695 ;
 RECT 1.02 0.595 1.25 0.805 ;
 RECT 0.68 0.09 0.78 1.38 ;
 RECT 0.84 1.59 0.94 2.62 ;
 RECT 0.68 1.38 0.94 1.59 ;
 RECT 3.925 0.535 4.025 2.12 ;
 RECT 3.75 0.325 4.025 0.535 ;
 RECT 4.395 0.27 4.495 0.965 ;
 RECT 4.865 1.065 4.965 2.74 ;
 RECT 4.395 1.275 4.495 2.74 ;
 RECT 4.865 0.27 4.965 0.965 ;
 RECT 4.395 0.965 4.965 1.065 ;
 RECT 4.235 1.065 4.495 1.275 ;
 RECT 3.085 0.915 3.185 2.625 ;
 RECT 2.31 0.09 2.41 0.755 ;
 RECT 2.955 0.705 3.185 0.755 ;
 RECT 2.955 0.855 3.185 0.915 ;
 RECT 2.31 0.755 3.185 0.855 ;
 RECT 2.01 0.09 2.11 0.615 ;
 RECT 2.01 0.825 2.11 1.035 ;
 RECT 2.615 1.135 2.715 2.625 ;
 RECT 1.88 0.615 2.11 0.825 ;
 RECT 2.01 1.035 2.715 1.135 ;
 LAYER CO ;
 RECT 3.675 1.53 3.805 1.66 ;
 RECT 4.145 2.38 4.275 2.51 ;
 RECT 3.8 0.365 3.93 0.495 ;
 RECT 0.12 2.235 0.25 2.365 ;
 RECT 5.575 0.47 5.705 0.6 ;
 RECT 5.5 1.635 5.63 1.765 ;
 RECT 4.145 0.715 4.275 0.845 ;
 RECT 1.06 2.245 1.19 2.375 ;
 RECT 0.12 0.31 0.25 0.44 ;
 RECT 2.53 0.31 2.66 0.44 ;
 RECT 2.36 2.265 2.49 2.395 ;
 RECT 2.835 1.95 2.965 2.08 ;
 RECT 5.575 0.73 5.705 0.86 ;
 RECT 1.495 0.625 1.625 0.755 ;
 RECT 0.28 1.585 0.41 1.715 ;
 RECT 3.305 2.265 3.435 2.395 ;
 RECT 4.615 2 4.745 2.13 ;
 RECT 4.615 2.26 4.745 2.39 ;
 RECT 3.675 0.715 3.805 0.845 ;
 RECT 0.9 0.31 1.03 0.44 ;
 RECT 5.5 1.895 5.63 2.025 ;
 RECT 1.93 0.655 2.06 0.785 ;
 RECT 1.89 1.955 2.02 2.085 ;
 RECT 5.5 2.155 5.63 2.285 ;
 RECT 0.73 1.42 0.86 1.55 ;
 RECT 4.285 1.105 4.415 1.235 ;
 RECT 3.005 0.745 3.135 0.875 ;
 RECT 4.615 1.74 4.745 1.87 ;
 RECT 5.085 2.12 5.215 2.25 ;
 RECT 4.145 2.12 4.275 2.25 ;
 RECT 5.085 0.51 5.215 0.64 ;
 RECT 5.085 2.38 5.215 2.51 ;
 RECT 4.615 0.655 4.745 0.785 ;
 RECT 0.59 2.22 0.72 2.35 ;
 RECT 1.07 0.635 1.2 0.765 ;
 RECT 1.42 2.265 1.55 2.395 ;
 RECT 1.76 0.31 1.89 0.44 ;
 LAYER M1 ;
 RECT 0.585 2.055 0.725 2.4 ;
 RECT 1.885 1.89 2.025 1.915 ;
 RECT 1.885 2.055 2.025 2.215 ;
 RECT 0.585 1.915 2.025 2.055 ;
 RECT 2.355 2.205 2.495 2.515 ;
 RECT 3.3 2.21 3.44 2.515 ;
 RECT 1.415 2.215 1.555 2.515 ;
 RECT 1.415 2.515 3.44 2.655 ;
 RECT 3.67 0.66 3.81 1.095 ;
 RECT 3.67 1.235 3.81 1.72 ;
 RECT 3.67 1.095 4.425 1.235 ;
 RECT 4.28 1.055 4.42 1.095 ;
 RECT 4.28 1.235 4.42 1.285 ;
 RECT 0.4 0.445 0.54 1.07 ;
 RECT 0.4 0.305 1.085 0.445 ;
 RECT 2.525 0.36 2.665 1.07 ;
 RECT 2.525 1.21 2.665 1.245 ;
 RECT 0.4 1.07 2.665 1.21 ;
 RECT 2.83 1.385 2.97 2.145 ;
 RECT 2.525 1.245 2.97 1.385 ;
 RECT 3.745 0.36 3.985 0.5 ;
 RECT 2.525 0.22 3.985 0.36 ;
 END
END AOI222X2

MACRO AOI22X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 3.195 0.08 3.335 0.665 ;
 RECT 4.08 0.08 4.22 0.78 ;
 RECT 1.755 0.08 1.895 0.865 ;
 RECT 0.115 0.08 0.255 0.865 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 4.08 1.585 4.22 2.8 ;
 RECT 3.195 2.31 3.335 2.8 ;
 RECT 0.115 2.21 0.255 2.8 ;
 RECT 1.055 2.21 1.195 2.8 ;
 END
 END VDD

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.89 1.48 2.2 1.765 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END IN4

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.155 0.46 1.4 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END IN2

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.175 0.32 1.565 0.76 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END IN3

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.435 0.96 1.72 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END IN1

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.56 0.78 3.805 1.02 ;
 RECT 3.665 0.62 3.805 0.78 ;
 RECT 3.665 1.02 3.805 1.985 ;
 END
 ANTENNADIFFAREA 0.465 ;
 END QN

 OBS
 LAYER PO ;
 RECT 3.45 1.38 3.55 2.76 ;
 RECT 3.45 0.265 3.55 1.17 ;
 RECT 3.27 1.17 3.55 1.38 ;
 RECT 0.68 0.45 0.78 1.545 ;
 RECT 0.84 1.795 0.94 2.62 ;
 RECT 0.68 1.545 0.91 1.695 ;
 RECT 0.68 1.695 0.94 1.795 ;
 RECT 1.98 1.545 2.24 1.755 ;
 RECT 1.54 0.45 1.64 1.265 ;
 RECT 2.14 1.755 2.24 2.62 ;
 RECT 2.14 1.365 2.24 1.545 ;
 RECT 1.54 1.265 2.24 1.365 ;
 RECT 1.67 1.645 1.77 2.62 ;
 RECT 1.15 0.54 1.25 1.545 ;
 RECT 1.15 1.545 1.77 1.645 ;
 RECT 1.13 0.33 1.36 0.54 ;
 RECT 0.37 1.39 0.47 2.62 ;
 RECT 0.37 0.45 0.47 1.18 ;
 RECT 0.23 1.18 0.47 1.39 ;
 RECT 2.98 0.555 3.08 0.985 ;
 RECT 2.98 1.085 3.08 1.94 ;
 RECT 2.31 0.875 2.54 0.985 ;
 RECT 2.31 0.985 3.08 1.085 ;
 LAYER CO ;
 RECT 3.67 1.8 3.8 1.93 ;
 RECT 3.32 1.21 3.45 1.34 ;
 RECT 3.67 0.68 3.8 0.81 ;
 RECT 3.67 1.54 3.8 1.67 ;
 RECT 2.36 2.26 2.49 2.39 ;
 RECT 4.085 1.635 4.215 1.765 ;
 RECT 0.59 2.26 0.72 2.39 ;
 RECT 0.73 1.585 0.86 1.715 ;
 RECT 1.76 0.67 1.89 0.8 ;
 RECT 0.12 0.67 0.25 0.8 ;
 RECT 0.12 2.26 0.25 2.39 ;
 RECT 4.085 1.895 4.215 2.025 ;
 RECT 2.36 0.915 2.49 1.045 ;
 RECT 3.2 2.37 3.33 2.5 ;
 RECT 3.2 0.485 3.33 0.615 ;
 RECT 2.03 1.585 2.16 1.715 ;
 RECT 4.085 0.34 4.215 0.47 ;
 RECT 1.89 2.16 2.02 2.29 ;
 RECT 4.085 0.6 4.215 0.73 ;
 RECT 1.18 0.37 1.31 0.5 ;
 RECT 0.9 0.67 1.03 0.8 ;
 RECT 2.73 0.695 2.86 0.825 ;
 RECT 2.73 1.56 2.86 1.69 ;
 RECT 1.06 2.26 1.19 2.39 ;
 RECT 0.28 1.22 0.41 1.35 ;
 RECT 1.42 2.26 1.55 2.39 ;
 RECT 4.085 2.155 4.215 2.285 ;
 LAYER M1 ;
 RECT 0.585 2.07 0.725 2.445 ;
 RECT 1.885 2.07 2.025 2.345 ;
 RECT 0.585 1.93 2.025 2.07 ;
 RECT 2.725 0.645 2.865 1.205 ;
 RECT 2.725 1.345 2.865 1.74 ;
 RECT 3.315 1.16 3.455 1.205 ;
 RECT 3.315 1.345 3.455 1.39 ;
 RECT 2.725 1.205 3.455 1.345 ;
 RECT 0.895 0.615 1.035 1.04 ;
 RECT 1.415 2.21 1.555 2.485 ;
 RECT 2.355 1.18 2.495 2.485 ;
 RECT 2.355 0.865 2.495 1.04 ;
 RECT 1.415 2.485 2.495 2.625 ;
 RECT 0.895 1.04 2.495 1.18 ;
 END
END AOI22X1

MACRO AOI22X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.17 1.48 1.575 1.72 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END IN3

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.31 0.79 1.615 1.045 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END IN4

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.16 1.48 0.44 1.745 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.48 1.03 1.72 ;
 END
 ANTENNAGATEAREA 0.056 ;
 END IN1

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 4.59 0.08 4.73 0.78 ;
 RECT 3.225 0.08 3.365 0.78 ;
 RECT 4.165 0.08 4.305 0.775 ;
 RECT 1.755 0.08 1.895 0.735 ;
 RECT 0.115 0.08 0.255 0.735 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.695 1.4 3.835 2.44 ;
 RECT 3.695 1.16 4.12 1.4 ;
 RECT 3.695 0.54 3.835 1.16 ;
 END
 ANTENNADIFFAREA 0.574 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 4.59 1.585 4.73 2.8 ;
 RECT 3.225 2.05 3.365 2.8 ;
 RECT 4.165 2.05 4.305 2.8 ;
 RECT 0.115 2.21 0.255 2.8 ;
 RECT 1.055 2.21 1.195 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 2.16 1.365 2.26 2.62 ;
 RECT 1.54 0.335 1.64 0.8 ;
 RECT 1.54 1.085 1.64 1.265 ;
 RECT 1.54 1.265 2.26 1.365 ;
 RECT 1.43 0.8 1.66 1.085 ;
 RECT 0.68 0.335 0.78 1.53 ;
 RECT 0.84 1.795 0.94 2.62 ;
 RECT 0.68 1.53 0.91 1.695 ;
 RECT 0.68 1.695 0.94 1.795 ;
 RECT 3.29 1.17 3.58 1.28 ;
 RECT 3.29 1.28 4.05 1.38 ;
 RECT 3.95 1.38 4.05 2.76 ;
 RECT 3.48 1.38 3.58 2.76 ;
 RECT 3.48 0.35 3.58 1.17 ;
 RECT 3.95 0.35 4.05 1.28 ;
 RECT 1.15 0.335 1.25 1.485 ;
 RECT 1.69 1.645 1.79 2.62 ;
 RECT 1.15 1.485 1.4 1.545 ;
 RECT 1.15 1.645 1.4 1.695 ;
 RECT 1.15 1.545 1.79 1.645 ;
 RECT 0.37 0.335 0.47 1.5 ;
 RECT 0.37 1.71 0.47 2.62 ;
 RECT 0.21 1.5 0.47 1.71 ;
 RECT 3.01 0.64 3.11 1.9 ;
 RECT 2.875 1.9 3.11 2.11 ;
 LAYER CO ;
 RECT 3.23 2.11 3.36 2.24 ;
 RECT 3.7 1.74 3.83 1.87 ;
 RECT 4.17 2.11 4.3 2.24 ;
 RECT 3.7 2 3.83 2.13 ;
 RECT 4.17 0.595 4.3 0.725 ;
 RECT 4.17 2.37 4.3 2.5 ;
 RECT 1.47 0.86 1.6 0.99 ;
 RECT 3.7 0.595 3.83 0.725 ;
 RECT 0.12 2.26 0.25 2.39 ;
 RECT 0.12 0.555 0.25 0.685 ;
 RECT 1.22 1.525 1.35 1.655 ;
 RECT 3.34 1.21 3.47 1.34 ;
 RECT 3.23 2.37 3.36 2.5 ;
 RECT 4.595 0.6 4.725 0.73 ;
 RECT 3.23 0.595 3.36 0.725 ;
 RECT 0.26 1.54 0.39 1.67 ;
 RECT 4.595 0.34 4.725 0.47 ;
 RECT 4.595 1.895 4.725 2.025 ;
 RECT 0.73 1.57 0.86 1.7 ;
 RECT 2.76 0.78 2.89 0.91 ;
 RECT 1.06 2.26 1.19 2.39 ;
 RECT 0.9 0.555 1.03 0.685 ;
 RECT 1.44 2.2 1.57 2.33 ;
 RECT 4.595 2.155 4.725 2.285 ;
 RECT 3.7 2.26 3.83 2.39 ;
 RECT 2.925 1.94 3.055 2.07 ;
 RECT 2.38 2.2 2.51 2.33 ;
 RECT 4.595 1.635 4.725 1.765 ;
 RECT 1.91 2.2 2.04 2.33 ;
 RECT 0.59 2.26 0.72 2.39 ;
 RECT 1.76 0.555 1.89 0.685 ;
 RECT 2.76 1.555 2.89 1.685 ;
 LAYER M1 ;
 RECT 0.585 2.01 0.725 2.44 ;
 RECT 1.905 2.01 2.045 2.38 ;
 RECT 0.585 1.87 2.045 2.01 ;
 RECT 2.755 0.73 2.895 1.205 ;
 RECT 2.755 1.345 2.895 1.745 ;
 RECT 3.335 1.16 3.475 1.205 ;
 RECT 3.335 1.345 3.475 1.39 ;
 RECT 2.755 1.205 3.48 1.345 ;
 RECT 0.895 0.505 1.035 1.185 ;
 RECT 1.435 2.15 1.575 2.52 ;
 RECT 2.375 1.325 2.515 1.935 ;
 RECT 2.375 1.935 3.065 2.075 ;
 RECT 2.375 2.075 2.515 2.52 ;
 RECT 2.92 1.89 3.06 1.935 ;
 RECT 2.92 2.075 3.06 2.12 ;
 RECT 0.895 1.185 2.515 1.325 ;
 RECT 1.435 2.52 2.515 2.66 ;
 END
END AOI22X2

MACRO IBUFFX16
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.88 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 4.17 0.08 4.31 0.675 ;
 RECT 7.045 0.08 7.185 0.675 ;
 RECT 0.315 0.08 0.455 0.675 ;
 RECT 2.235 0.08 2.375 0.675 ;
 RECT 3.19 0.08 3.33 0.675 ;
 RECT 6.09 0.08 6.23 0.675 ;
 RECT 1.28 0.08 1.42 0.675 ;
 RECT 8.01 0.08 8.15 0.675 ;
 RECT 5.135 0.08 5.275 0.675 ;
 RECT 9.4 0.08 9.54 0.79 ;
 RECT 8.43 0.08 8.57 0.79 ;
 RECT 0 -0.08 10.88 0.08 ;
 RECT 10.28 0.08 10.42 0.795 ;
 END
 END VSS

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.53 0.515 7.67 0.84 ;
 RECT 6.575 0.84 7.67 0.865 ;
 RECT 6.575 0.515 6.715 0.84 ;
 RECT 7.53 1.085 7.67 2.36 ;
 RECT 6.575 1.085 6.715 2.36 ;
 RECT 6.575 1.005 7.67 1.085 ;
 RECT 5.62 1.005 5.76 2.36 ;
 RECT 5.62 0.515 5.76 0.865 ;
 RECT 4.655 1.005 4.795 2.36 ;
 RECT 4.655 0.515 4.795 0.865 ;
 RECT 3.675 1.005 3.815 2.36 ;
 RECT 3.675 0.515 3.815 0.865 ;
 RECT 1.765 1.005 1.905 2.36 ;
 RECT 1.765 0.515 1.905 0.865 ;
 RECT 0.8 1.005 0.94 2.36 ;
 RECT 0.8 0.865 7.67 1.005 ;
 RECT 0.8 0.515 0.94 0.865 ;
 RECT 2.72 1.005 2.86 2.36 ;
 RECT 2.72 0.515 2.86 0.865 ;
 END
 ANTENNADIFFAREA 4.784 ;
 END ZN

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.68 2.12 10.025 2.39 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END INP

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.88 2.96 ;
 RECT 9.4 1.84 9.54 2.8 ;
 RECT 8.43 1.84 8.57 2.8 ;
 RECT 10.295 1.535 10.435 2.8 ;
 RECT 8.035 1.91 8.175 2.8 ;
 RECT 4.17 1.91 4.31 2.8 ;
 RECT 6.09 1.91 6.23 2.8 ;
 RECT 7.045 1.91 7.185 2.8 ;
 RECT 3.19 1.91 3.33 2.8 ;
 RECT 1.28 1.91 1.42 2.8 ;
 RECT 0.315 1.91 0.455 2.8 ;
 RECT 2.235 1.91 2.375 2.8 ;
 RECT 5.135 1.91 5.275 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 4.425 0.23 4.525 1.23 ;
 RECT 4.425 1.33 4.525 2.74 ;
 RECT 0.57 1.23 7.885 1.33 ;
 RECT 2.49 0.23 2.59 1.23 ;
 RECT 2.49 1.33 2.59 2.74 ;
 RECT 1.535 0.23 1.635 1.23 ;
 RECT 1.535 1.33 1.635 2.74 ;
 RECT 3.445 0.23 3.545 1.23 ;
 RECT 3.445 1.33 3.545 2.74 ;
 RECT 1.055 0.23 1.155 1.23 ;
 RECT 1.055 1.33 1.155 2.74 ;
 RECT 7.785 1.18 7.885 1.23 ;
 RECT 7.785 1.33 7.885 2.74 ;
 RECT 0.57 0.23 0.67 1.23 ;
 RECT 2.975 0.23 3.075 1.23 ;
 RECT 2.02 0.23 2.12 1.23 ;
 RECT 3.93 0.23 4.03 1.23 ;
 RECT 6.345 0.23 6.445 1.23 ;
 RECT 5.39 0.23 5.49 1.23 ;
 RECT 4.91 0.23 5.01 1.23 ;
 RECT 6.83 0.23 6.93 1.23 ;
 RECT 5.875 0.23 5.975 1.23 ;
 RECT 7.3 0.23 7.4 1.23 ;
 RECT 0.57 1.33 0.67 2.74 ;
 RECT 2.975 1.33 3.075 2.74 ;
 RECT 2.02 1.33 2.12 2.74 ;
 RECT 3.93 1.33 4.03 2.74 ;
 RECT 6.345 1.33 6.445 2.74 ;
 RECT 5.39 1.33 5.49 2.74 ;
 RECT 4.91 1.33 5.01 2.74 ;
 RECT 6.83 1.33 6.93 2.74 ;
 RECT 5.875 1.33 5.975 2.74 ;
 RECT 7.3 1.33 7.4 2.74 ;
 RECT 7.785 0.23 7.885 0.95 ;
 RECT 7.785 0.95 8.04 1.18 ;
 RECT 8.69 0.255 8.79 1.2 ;
 RECT 8.69 1.2 9.285 1.3 ;
 RECT 8.69 1.3 8.79 2.76 ;
 RECT 9.185 0.255 9.285 1.12 ;
 RECT 9.055 1.12 9.285 1.2 ;
 RECT 9.055 1.3 9.285 1.35 ;
 RECT 9.185 1.35 9.285 2.755 ;
 RECT 9.655 0.385 9.755 2.16 ;
 RECT 9.655 2.16 9.885 2.39 ;
 LAYER CO ;
 RECT 10.285 0.615 10.415 0.745 ;
 RECT 7.535 1.95 7.665 2.08 ;
 RECT 6.095 0.495 6.225 0.625 ;
 RECT 4.175 0.495 4.305 0.625 ;
 RECT 4.66 1.95 4.79 2.08 ;
 RECT 6.58 1.95 6.71 2.08 ;
 RECT 10.3 1.845 10.43 1.975 ;
 RECT 5.14 0.495 5.27 0.625 ;
 RECT 4.66 1.645 4.79 1.775 ;
 RECT 2.24 0.495 2.37 0.625 ;
 RECT 1.77 0.565 1.9 0.695 ;
 RECT 6.095 1.96 6.225 2.09 ;
 RECT 10.285 0.355 10.415 0.485 ;
 RECT 9.405 0.605 9.535 0.735 ;
 RECT 2.725 0.565 2.855 0.695 ;
 RECT 3.68 1.645 3.81 1.775 ;
 RECT 2.24 1.96 2.37 2.09 ;
 RECT 5.625 1.645 5.755 1.775 ;
 RECT 1.285 0.495 1.415 0.625 ;
 RECT 10.3 2.105 10.43 2.235 ;
 RECT 3.68 1.645 3.81 1.775 ;
 RECT 1.285 1.96 1.415 2.09 ;
 RECT 5.625 1.95 5.755 2.08 ;
 RECT 7.535 1.645 7.665 1.775 ;
 RECT 0.805 1.95 0.935 2.08 ;
 RECT 0.805 1.645 0.935 1.775 ;
 RECT 0.805 0.565 0.935 0.695 ;
 RECT 6.58 1.645 6.71 1.775 ;
 RECT 7.535 1.645 7.665 1.775 ;
 RECT 3.68 1.95 3.81 2.08 ;
 RECT 9.875 0.605 10.005 0.735 ;
 RECT 10.3 1.585 10.43 1.715 ;
 RECT 2.725 1.645 2.855 1.775 ;
 RECT 9.875 1.75 10.005 1.88 ;
 RECT 1.77 1.645 1.9 1.775 ;
 RECT 2.725 1.645 2.855 1.775 ;
 RECT 9.705 2.21 9.835 2.34 ;
 RECT 4.66 1.645 4.79 1.775 ;
 RECT 7.05 0.495 7.18 0.625 ;
 RECT 9.405 1.9 9.535 2.03 ;
 RECT 8.435 0.605 8.565 0.735 ;
 RECT 8.435 1.9 8.565 2.03 ;
 RECT 3.68 0.565 3.81 0.695 ;
 RECT 1.77 1.95 1.9 2.08 ;
 RECT 4.66 0.565 4.79 0.695 ;
 RECT 7.86 1 7.99 1.13 ;
 RECT 4.175 1.96 4.305 2.09 ;
 RECT 0.32 0.495 0.45 0.625 ;
 RECT 7.535 0.565 7.665 0.695 ;
 RECT 9.105 1.17 9.235 1.3 ;
 RECT 8.04 1.96 8.17 2.09 ;
 RECT 5.625 1.645 5.755 1.775 ;
 RECT 6.58 0.565 6.71 0.695 ;
 RECT 2.725 1.95 2.855 2.08 ;
 RECT 8.915 1.705 9.045 1.835 ;
 RECT 6.58 1.645 6.71 1.775 ;
 RECT 3.195 0.495 3.325 0.625 ;
 RECT 0.32 1.96 0.45 2.09 ;
 RECT 0.805 1.645 0.935 1.775 ;
 RECT 8.915 1.705 9.045 1.835 ;
 RECT 5.14 1.96 5.27 2.09 ;
 RECT 1.77 1.645 1.9 1.775 ;
 RECT 8.915 0.605 9.045 0.735 ;
 RECT 7.05 1.96 7.18 2.09 ;
 RECT 3.195 1.96 3.325 2.09 ;
 RECT 8.015 0.495 8.145 0.625 ;
 RECT 5.625 0.565 5.755 0.695 ;
 LAYER M1 ;
 RECT 9.19 1.085 9.33 1.12 ;
 RECT 9.19 1.35 9.33 1.54 ;
 RECT 9.1 1.12 9.33 1.35 ;
 RECT 9.87 0.555 10.01 1.54 ;
 RECT 9.19 1.54 10.01 1.68 ;
 RECT 9.87 1.68 10.01 1.93 ;
 RECT 7.855 1.09 7.995 1.18 ;
 RECT 7.855 0.975 8.96 1.09 ;
 RECT 7.855 0.95 9.05 0.975 ;
 RECT 8.91 1.685 9.05 1.885 ;
 RECT 8.82 1.09 8.96 1.545 ;
 RECT 8.82 0.835 9.05 0.95 ;
 RECT 8.91 0.515 9.05 0.835 ;
 RECT 8.82 1.545 9.05 1.685 ;
 END
END IBUFFX16

MACRO IBUFFX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.395 2.095 2.795 2.39 ;
 END
 ANTENNAGATEAREA 0.076 ;
 END INP

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.41 0.835 0.875 1.085 ;
 RECT 0.735 0.515 0.875 0.835 ;
 RECT 0.735 1.085 0.875 2.36 ;
 END
 ANTENNADIFFAREA 0.606 ;
 END ZN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 2.115 0.08 2.255 0.79 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 1.215 0.08 1.355 0.675 ;
 RECT 0.25 0.08 0.39 0.675 ;
 RECT 2.995 0.08 3.135 0.795 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 2.115 1.84 2.255 2.8 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 1.24 1.91 1.38 2.8 ;
 RECT 0.25 1.91 0.39 2.8 ;
 RECT 3.01 1.535 3.15 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.99 1.18 1.09 1.23 ;
 RECT 0.99 1.33 1.09 2.74 ;
 RECT 0.505 1.23 1.09 1.33 ;
 RECT 0.505 0.23 0.605 1.23 ;
 RECT 0.99 0.215 1.09 0.95 ;
 RECT 0.505 1.33 0.605 2.74 ;
 RECT 0.99 0.95 1.245 1.18 ;
 RECT 2.37 0.385 2.47 2.16 ;
 RECT 2.37 2.16 2.6 2.39 ;
 RECT 1.9 0.38 2 1.12 ;
 RECT 1.9 1.35 2 2.305 ;
 RECT 1.77 1.12 2 1.35 ;
 LAYER CO ;
 RECT 3.015 2.105 3.145 2.235 ;
 RECT 3 0.355 3.13 0.485 ;
 RECT 3.015 1.845 3.145 1.975 ;
 RECT 3.015 1.585 3.145 1.715 ;
 RECT 3 0.615 3.13 0.745 ;
 RECT 2.12 0.605 2.25 0.735 ;
 RECT 0.255 0.495 0.385 0.625 ;
 RECT 0.255 1.96 0.385 2.09 ;
 RECT 1.065 1 1.195 1.13 ;
 RECT 0.74 1.95 0.87 2.08 ;
 RECT 0.74 1.645 0.87 1.775 ;
 RECT 0.74 0.565 0.87 0.695 ;
 RECT 0.74 1.645 0.87 1.775 ;
 RECT 1.245 1.96 1.375 2.09 ;
 RECT 1.63 0.605 1.76 0.735 ;
 RECT 2.12 1.9 2.25 2.03 ;
 RECT 2.42 2.21 2.55 2.34 ;
 RECT 1.82 1.17 1.95 1.3 ;
 RECT 1.63 1.705 1.76 1.835 ;
 RECT 1.22 0.495 1.35 0.625 ;
 RECT 2.59 1.75 2.72 1.88 ;
 RECT 1.63 1.705 1.76 1.835 ;
 RECT 2.59 0.605 2.72 0.735 ;
 LAYER M1 ;
 RECT 1.905 1.11 2.045 1.12 ;
 RECT 1.905 1.35 2.045 1.54 ;
 RECT 1.815 1.12 2.045 1.35 ;
 RECT 2.585 0.555 2.725 1.54 ;
 RECT 1.905 1.54 2.725 1.68 ;
 RECT 2.585 1.68 2.725 1.93 ;
 RECT 1.045 0.95 1.765 0.975 ;
 RECT 1.045 1.09 1.245 1.18 ;
 RECT 1.045 0.975 1.675 1.09 ;
 RECT 1.625 0.515 1.765 0.835 ;
 RECT 1.535 0.835 1.765 0.95 ;
 RECT 1.535 1.09 1.675 1.545 ;
 RECT 1.625 1.685 1.765 1.885 ;
 RECT 1.535 1.545 1.765 1.685 ;
 END
END IBUFFX2

MACRO IBUFFX32
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 19.52 BY 2.88 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.315 2.07 18.725 2.39 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END INP

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 15.215 1.08 15.355 2.36 ;
 RECT 13.305 1.005 13.445 2.36 ;
 RECT 14.26 1.005 14.4 2.36 ;
 RECT 12.34 1.005 12.48 2.36 ;
 RECT 14.745 1.005 15.355 1.08 ;
 RECT 11.36 1.005 11.5 2.36 ;
 RECT 10.405 1.005 10.545 2.36 ;
 RECT 8.485 1.005 8.625 2.36 ;
 RECT 9.45 1.005 9.59 2.36 ;
 RECT 7.51 1.005 7.65 2.36 ;
 RECT 3.655 1.005 3.795 2.36 ;
 RECT 4.635 1.005 4.775 2.36 ;
 RECT 6.555 1.005 6.695 2.36 ;
 RECT 5.6 1.005 5.74 2.36 ;
 RECT 1.745 1.005 1.885 2.36 ;
 RECT 2.7 1.005 2.84 2.36 ;
 RECT 0.78 1.005 0.92 2.36 ;
 RECT 0.78 0.865 15.355 1.005 ;
 RECT 14.745 0.84 15.355 0.865 ;
 RECT 13.305 0.515 13.445 0.865 ;
 RECT 15.215 0.515 15.355 0.84 ;
 RECT 14.26 0.515 14.4 0.865 ;
 RECT 12.34 0.515 12.48 0.865 ;
 RECT 11.36 0.515 11.5 0.865 ;
 RECT 10.405 0.515 10.545 0.865 ;
 RECT 8.485 0.515 8.625 0.865 ;
 RECT 9.45 0.515 9.59 0.865 ;
 RECT 7.51 0.515 7.65 0.865 ;
 RECT 3.655 0.515 3.795 0.865 ;
 RECT 4.635 0.515 4.775 0.865 ;
 RECT 6.555 0.515 6.695 0.865 ;
 RECT 5.6 0.515 5.74 0.865 ;
 RECT 1.745 0.515 1.885 0.865 ;
 RECT 2.7 0.515 2.84 0.865 ;
 RECT 0.78 0.515 0.92 0.865 ;
 END
 ANTENNADIFFAREA 9.568 ;
 END ZN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 10.875 0.08 11.015 0.675 ;
 RECT 12.82 0.08 12.96 0.675 ;
 RECT 5.115 0.08 5.255 0.675 ;
 RECT 6.07 0.08 6.21 0.675 ;
 RECT 7.025 0.08 7.165 0.675 ;
 RECT 3.17 0.08 3.31 0.675 ;
 RECT 1.26 0.08 1.4 0.675 ;
 RECT 2.215 0.08 2.355 0.675 ;
 RECT 11.855 0.08 11.995 0.675 ;
 RECT 8 0.08 8.14 0.675 ;
 RECT 15.695 0.08 15.835 0.675 ;
 RECT 9.92 0.08 10.06 0.675 ;
 RECT 8.965 0.08 9.105 0.675 ;
 RECT 4.15 0.08 4.29 0.675 ;
 RECT 0.295 0.08 0.435 0.675 ;
 RECT 14.73 0.08 14.87 0.675 ;
 RECT 13.775 0.08 13.915 0.675 ;
 RECT 18.035 0.08 18.175 0.79 ;
 RECT 0 -0.08 19.52 0.08 ;
 RECT 17.065 0.08 17.205 0.79 ;
 RECT 16.07 0.08 16.21 0.79 ;
 RECT 18.915 0.08 19.055 0.795 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 8 1.91 8.14 2.8 ;
 RECT 18.035 1.84 18.175 2.8 ;
 RECT 18.93 1.535 19.07 2.8 ;
 RECT 0 2.8 19.52 2.96 ;
 RECT 17.065 1.84 17.205 2.8 ;
 RECT 16.1 1.84 16.24 2.8 ;
 RECT 10.875 1.91 11.015 2.8 ;
 RECT 7.025 1.91 7.165 2.8 ;
 RECT 3.17 1.91 3.31 2.8 ;
 RECT 6.07 1.91 6.21 2.8 ;
 RECT 1.26 1.91 1.4 2.8 ;
 RECT 9.92 1.91 10.06 2.8 ;
 RECT 11.855 1.91 11.995 2.8 ;
 RECT 15.72 1.91 15.86 2.8 ;
 RECT 2.215 1.91 2.355 2.8 ;
 RECT 12.82 1.91 12.96 2.8 ;
 RECT 8.965 1.91 9.105 2.8 ;
 RECT 14.73 1.91 14.87 2.8 ;
 RECT 5.115 1.91 5.255 2.8 ;
 RECT 4.15 1.91 4.29 2.8 ;
 RECT 13.775 1.91 13.915 2.8 ;
 RECT 0.295 1.91 0.435 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 17.82 0.25 17.92 1.12 ;
 RECT 17.82 1.35 17.92 2.745 ;
 RECT 16.36 0.25 16.46 1.145 ;
 RECT 16.36 1.145 17.92 1.245 ;
 RECT 16.36 1.245 16.46 2.745 ;
 RECT 16.85 0.25 16.95 1.145 ;
 RECT 16.85 1.245 16.95 2.755 ;
 RECT 17.33 0.25 17.43 1.145 ;
 RECT 17.33 1.245 17.43 2.76 ;
 RECT 17.69 1.12 17.92 1.145 ;
 RECT 17.69 1.245 17.92 1.35 ;
 RECT 3.425 0.23 3.525 1.23 ;
 RECT 1.515 0.23 1.615 1.23 ;
 RECT 1.035 0.23 1.135 1.23 ;
 RECT 2.47 0.23 2.57 1.23 ;
 RECT 0.55 0.23 0.65 1.23 ;
 RECT 2.955 0.23 3.055 1.23 ;
 RECT 2 0.23 2.1 1.23 ;
 RECT 3.91 0.23 4.01 1.23 ;
 RECT 6.325 0.23 6.425 1.23 ;
 RECT 4.405 0.23 4.505 1.23 ;
 RECT 5.37 0.23 5.47 1.23 ;
 RECT 7.28 0.23 7.38 1.23 ;
 RECT 5.855 0.23 5.955 1.23 ;
 RECT 4.89 0.23 4.99 1.23 ;
 RECT 6.81 0.23 6.91 1.23 ;
 RECT 7.765 0.23 7.865 1.23 ;
 RECT 11.13 0.23 11.23 1.23 ;
 RECT 8.74 0.23 8.84 1.23 ;
 RECT 9.22 0.23 9.32 1.23 ;
 RECT 10.175 0.23 10.275 1.23 ;
 RECT 9.705 0.23 9.805 1.23 ;
 RECT 10.66 0.23 10.76 1.23 ;
 RECT 8.255 0.23 8.355 1.23 ;
 RECT 11.615 0.23 11.715 1.23 ;
 RECT 13.075 0.23 13.175 1.23 ;
 RECT 12.595 0.23 12.695 1.23 ;
 RECT 12.11 0.23 12.21 1.23 ;
 RECT 13.56 0.23 13.66 1.23 ;
 RECT 14.985 0.23 15.085 1.23 ;
 RECT 14.515 0.23 14.615 1.23 ;
 RECT 14.03 0.23 14.13 1.23 ;
 RECT 15.47 0.23 15.57 0.95 ;
 RECT 15.47 0.95 15.725 1.18 ;
 RECT 15.47 1.18 15.57 1.23 ;
 RECT 3.425 1.33 3.525 2.74 ;
 RECT 1.515 1.33 1.615 2.74 ;
 RECT 1.035 1.33 1.135 2.74 ;
 RECT 2.47 1.33 2.57 2.74 ;
 RECT 0.55 1.33 0.65 2.74 ;
 RECT 2.955 1.33 3.055 2.74 ;
 RECT 2 1.33 2.1 2.74 ;
 RECT 3.91 1.33 4.01 2.74 ;
 RECT 6.325 1.33 6.425 2.74 ;
 RECT 4.405 1.33 4.505 2.74 ;
 RECT 5.37 1.33 5.47 2.74 ;
 RECT 7.28 1.33 7.38 2.74 ;
 RECT 5.855 1.33 5.955 2.74 ;
 RECT 4.89 1.33 4.99 2.74 ;
 RECT 6.81 1.33 6.91 2.74 ;
 RECT 7.765 1.33 7.865 2.74 ;
 RECT 11.13 1.33 11.23 2.74 ;
 RECT 8.74 1.33 8.84 2.74 ;
 RECT 9.22 1.33 9.32 2.74 ;
 RECT 10.175 1.33 10.275 2.74 ;
 RECT 9.705 1.33 9.805 2.74 ;
 RECT 10.66 1.33 10.76 2.74 ;
 RECT 8.255 1.33 8.355 2.74 ;
 RECT 11.615 1.33 11.715 2.74 ;
 RECT 13.075 1.33 13.175 2.74 ;
 RECT 12.595 1.33 12.695 2.74 ;
 RECT 12.11 1.33 12.21 2.74 ;
 RECT 13.56 1.33 13.66 2.74 ;
 RECT 14.985 1.33 15.085 2.74 ;
 RECT 14.515 1.33 14.615 2.74 ;
 RECT 14.03 1.33 14.13 2.74 ;
 RECT 15.47 1.33 15.57 2.74 ;
 RECT 0.55 1.23 15.57 1.33 ;
 RECT 18.29 0.385 18.39 2.16 ;
 RECT 18.29 2.16 18.52 2.39 ;
 LAYER CO ;
 RECT 0.3 1.96 0.43 2.09 ;
 RECT 0.785 1.95 0.915 2.08 ;
 RECT 1.265 1.96 1.395 2.09 ;
 RECT 0.785 1.645 0.915 1.775 ;
 RECT 6.075 0.495 6.205 0.625 ;
 RECT 4.155 1.96 4.285 2.09 ;
 RECT 17.07 1.9 17.2 2.03 ;
 RECT 10.41 1.95 10.54 2.08 ;
 RECT 15.545 1 15.675 1.13 ;
 RECT 1.265 0.495 1.395 0.625 ;
 RECT 2.22 0.495 2.35 0.625 ;
 RECT 7.515 1.645 7.645 1.775 ;
 RECT 3.66 1.645 3.79 1.775 ;
 RECT 2.705 1.645 2.835 1.775 ;
 RECT 3.66 1.645 3.79 1.775 ;
 RECT 4.64 1.645 4.77 1.775 ;
 RECT 7.03 1.96 7.16 2.09 ;
 RECT 4.64 1.645 4.77 1.775 ;
 RECT 6.075 1.96 6.205 2.09 ;
 RECT 6.56 1.645 6.69 1.775 ;
 RECT 17.74 1.17 17.87 1.3 ;
 RECT 11.365 0.565 11.495 0.695 ;
 RECT 11.86 0.495 11.99 0.625 ;
 RECT 8.49 1.645 8.62 1.775 ;
 RECT 11.365 1.645 11.495 1.775 ;
 RECT 17.55 1.705 17.68 1.835 ;
 RECT 8.005 1.96 8.135 2.09 ;
 RECT 15.7 0.495 15.83 0.625 ;
 RECT 10.41 1.645 10.54 1.775 ;
 RECT 18.935 1.845 19.065 1.975 ;
 RECT 8.49 1.95 8.62 2.08 ;
 RECT 12.345 0.565 12.475 0.695 ;
 RECT 9.455 1.645 9.585 1.775 ;
 RECT 1.75 1.645 1.88 1.775 ;
 RECT 12.345 1.95 12.475 2.08 ;
 RECT 13.31 1.95 13.44 2.08 ;
 RECT 8.005 0.495 8.135 0.625 ;
 RECT 15.22 1.645 15.35 1.775 ;
 RECT 18.34 2.21 18.47 2.34 ;
 RECT 12.345 1.645 12.475 1.775 ;
 RECT 9.455 1.95 9.585 2.08 ;
 RECT 14.735 0.495 14.865 0.625 ;
 RECT 10.41 1.645 10.54 1.775 ;
 RECT 16.105 1.9 16.235 2.03 ;
 RECT 16.075 0.605 16.205 0.735 ;
 RECT 16.58 1.705 16.71 1.835 ;
 RECT 16.58 1.705 16.71 1.835 ;
 RECT 16.58 0.605 16.71 0.735 ;
 RECT 18.04 0.605 18.17 0.735 ;
 RECT 4.155 0.495 4.285 0.625 ;
 RECT 5.605 1.645 5.735 1.775 ;
 RECT 18.935 2.105 19.065 2.235 ;
 RECT 1.75 1.645 1.88 1.775 ;
 RECT 8.97 0.495 9.1 0.625 ;
 RECT 17.55 0.605 17.68 0.735 ;
 RECT 13.31 1.645 13.44 1.775 ;
 RECT 11.365 1.95 11.495 2.08 ;
 RECT 8.97 1.96 9.1 2.09 ;
 RECT 10.41 0.565 10.54 0.695 ;
 RECT 10.88 0.495 11.01 0.625 ;
 RECT 8.49 0.565 8.62 0.695 ;
 RECT 9.925 0.495 10.055 0.625 ;
 RECT 13.78 0.495 13.91 0.625 ;
 RECT 2.705 1.95 2.835 2.08 ;
 RECT 5.605 0.565 5.735 0.695 ;
 RECT 18.04 1.9 18.17 2.03 ;
 RECT 5.12 0.495 5.25 0.625 ;
 RECT 12.825 0.495 12.955 0.625 ;
 RECT 13.31 1.645 13.44 1.775 ;
 RECT 18.51 0.605 18.64 0.735 ;
 RECT 4.64 1.95 4.77 2.08 ;
 RECT 18.935 1.585 19.065 1.715 ;
 RECT 7.03 0.495 7.16 0.625 ;
 RECT 4.64 0.565 4.77 0.695 ;
 RECT 0.785 1.645 0.915 1.775 ;
 RECT 2.705 1.645 2.835 1.775 ;
 RECT 6.56 1.645 6.69 1.775 ;
 RECT 5.605 1.645 5.735 1.775 ;
 RECT 5.605 1.95 5.735 2.08 ;
 RECT 2.705 0.565 2.835 0.695 ;
 RECT 1.75 0.565 1.88 0.695 ;
 RECT 7.515 0.565 7.645 0.695 ;
 RECT 7.515 1.645 7.645 1.775 ;
 RECT 3.175 0.495 3.305 0.625 ;
 RECT 6.56 1.95 6.69 2.08 ;
 RECT 0.3 0.495 0.43 0.625 ;
 RECT 2.22 1.96 2.35 2.09 ;
 RECT 9.455 0.565 9.585 0.695 ;
 RECT 17.55 1.705 17.68 1.835 ;
 RECT 15.22 0.565 15.35 0.695 ;
 RECT 9.925 1.96 10.055 2.09 ;
 RECT 9.455 1.645 9.585 1.775 ;
 RECT 15.725 1.96 15.855 2.09 ;
 RECT 15.22 1.95 15.35 2.08 ;
 RECT 14.735 1.96 14.865 2.09 ;
 RECT 18.92 0.355 19.05 0.485 ;
 RECT 13.31 0.565 13.44 0.695 ;
 RECT 10.88 1.96 11.01 2.09 ;
 RECT 8.49 1.645 8.62 1.775 ;
 RECT 12.345 1.645 12.475 1.775 ;
 RECT 13.78 1.96 13.91 2.09 ;
 RECT 14.265 1.645 14.395 1.775 ;
 RECT 12.825 1.96 12.955 2.09 ;
 RECT 14.265 0.565 14.395 0.695 ;
 RECT 11.86 1.96 11.99 2.09 ;
 RECT 18.51 1.75 18.64 1.88 ;
 RECT 15.22 1.645 15.35 1.775 ;
 RECT 17.07 0.605 17.2 0.735 ;
 RECT 5.12 1.96 5.25 2.09 ;
 RECT 18.92 0.615 19.05 0.745 ;
 RECT 14.265 1.645 14.395 1.775 ;
 RECT 14.265 1.95 14.395 2.08 ;
 RECT 3.66 0.565 3.79 0.695 ;
 RECT 0.785 0.565 0.915 0.695 ;
 RECT 11.365 1.645 11.495 1.775 ;
 RECT 7.515 1.95 7.645 2.08 ;
 RECT 3.66 1.95 3.79 2.08 ;
 RECT 3.175 1.96 3.305 2.09 ;
 RECT 6.56 0.565 6.69 0.695 ;
 RECT 1.75 1.95 1.88 2.08 ;
 LAYER M1 ;
 RECT 16.575 1.09 16.715 1.885 ;
 RECT 16.575 0.515 16.715 0.95 ;
 RECT 15.54 1.09 15.68 1.18 ;
 RECT 17.545 1.685 17.685 1.885 ;
 RECT 17.455 1.09 17.595 1.545 ;
 RECT 15.54 0.975 17.595 1.09 ;
 RECT 15.54 0.95 17.685 0.975 ;
 RECT 17.455 0.835 17.685 0.95 ;
 RECT 17.545 0.515 17.685 0.835 ;
 RECT 17.455 1.545 17.685 1.685 ;
 RECT 17.825 1.085 17.965 1.12 ;
 RECT 17.735 1.12 17.965 1.35 ;
 RECT 17.825 1.35 17.965 1.54 ;
 RECT 18.505 1.68 18.645 1.93 ;
 RECT 18.505 0.555 18.645 1.54 ;
 RECT 17.825 1.54 18.645 1.68 ;
 END
END IBUFFX32

MACRO IBUFFX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.355 2.12 3.755 2.39 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END INP

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 3.075 1.84 3.215 2.8 ;
 RECT 3.97 1.535 4.11 2.8 ;
 RECT 1.21 1.91 1.35 2.8 ;
 RECT 2.2 1.91 2.34 2.8 ;
 RECT 0.255 1.91 0.395 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 2.175 0.08 2.315 0.675 ;
 RECT 1.21 0.08 1.35 0.675 ;
 RECT 0.255 0.08 0.395 0.675 ;
 RECT 3.075 0.08 3.215 0.79 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 3.955 0.08 4.095 0.795 ;
 END
 END VSS

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.74 0.965 1.835 1.105 ;
 RECT 1.695 0.515 1.835 0.965 ;
 RECT 0.74 0.515 0.88 0.835 ;
 RECT 0.74 0.835 1.155 0.965 ;
 RECT 0.74 1.105 0.88 2.36 ;
 RECT 1.695 1.105 1.835 2.36 ;
 END
 ANTENNADIFFAREA 1.196 ;
 END ZN

 OBS
 LAYER PO ;
 RECT 3.33 0.385 3.43 2.16 ;
 RECT 3.33 2.16 3.56 2.39 ;
 RECT 1.95 1.18 2.05 1.23 ;
 RECT 1.95 1.33 2.05 2.74 ;
 RECT 0.51 1.23 2.05 1.33 ;
 RECT 0.51 0.23 0.61 1.23 ;
 RECT 0.995 0.23 1.095 1.23 ;
 RECT 1.465 0.23 1.565 1.23 ;
 RECT 1.95 0.23 2.05 0.95 ;
 RECT 0.51 1.33 0.61 2.74 ;
 RECT 0.995 1.33 1.095 2.74 ;
 RECT 1.465 1.33 1.565 2.74 ;
 RECT 1.95 0.95 2.205 1.18 ;
 RECT 2.86 0.32 2.96 1.12 ;
 RECT 2.86 1.35 2.96 2.755 ;
 RECT 2.73 1.12 2.96 1.35 ;
 LAYER CO ;
 RECT 0.745 1.645 0.875 1.775 ;
 RECT 0.26 1.96 0.39 2.09 ;
 RECT 0.26 0.495 0.39 0.625 ;
 RECT 0.745 0.565 0.875 0.695 ;
 RECT 0.745 1.95 0.875 2.08 ;
 RECT 0.745 1.645 0.875 1.775 ;
 RECT 2.78 1.17 2.91 1.3 ;
 RECT 1.215 1.96 1.345 2.09 ;
 RECT 3.975 2.105 4.105 2.235 ;
 RECT 3.975 1.845 4.105 1.975 ;
 RECT 1.7 1.645 1.83 1.775 ;
 RECT 3.38 2.21 3.51 2.34 ;
 RECT 3.55 0.605 3.68 0.735 ;
 RECT 2.59 1.705 2.72 1.835 ;
 RECT 2.59 1.705 2.72 1.835 ;
 RECT 3.08 0.605 3.21 0.735 ;
 RECT 3.96 0.615 4.09 0.745 ;
 RECT 3.96 0.355 4.09 0.485 ;
 RECT 1.7 0.565 1.83 0.695 ;
 RECT 1.7 1.95 1.83 2.08 ;
 RECT 3.55 1.75 3.68 1.88 ;
 RECT 2.59 0.605 2.72 0.735 ;
 RECT 3.975 1.585 4.105 1.715 ;
 RECT 1.215 0.495 1.345 0.625 ;
 RECT 2.205 1.96 2.335 2.09 ;
 RECT 2.025 1 2.155 1.13 ;
 RECT 3.08 1.9 3.21 2.03 ;
 RECT 2.18 0.495 2.31 0.625 ;
 RECT 1.7 1.645 1.83 1.775 ;
 LAYER M1 ;
 RECT 2.865 1.085 3.005 1.12 ;
 RECT 2.775 1.12 3.005 1.35 ;
 RECT 2.865 1.35 3.005 1.54 ;
 RECT 3.545 1.68 3.685 1.93 ;
 RECT 3.545 0.555 3.685 1.54 ;
 RECT 2.865 1.54 3.685 1.68 ;
 RECT 2.02 1.09 2.16 1.18 ;
 RECT 2.585 0.515 2.725 0.835 ;
 RECT 2.585 1.685 2.725 1.885 ;
 RECT 2.495 0.835 2.725 0.95 ;
 RECT 2.01 0.95 2.725 0.975 ;
 RECT 2.01 0.975 2.635 1.09 ;
 RECT 2.495 1.09 2.635 1.545 ;
 RECT 2.495 1.545 2.725 1.685 ;
 END
END IBUFFX4

MACRO IBUFFX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.4 BY 2.88 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.205 2.07 5.61 2.39 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END INP

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 4.925 1.84 5.065 2.8 ;
 RECT 0 2.8 6.4 2.96 ;
 RECT 4.05 1.91 4.19 2.8 ;
 RECT 3.06 1.91 3.2 2.8 ;
 RECT 2.105 1.91 2.245 2.8 ;
 RECT 1.15 1.91 1.29 2.8 ;
 RECT 0.185 1.91 0.325 2.8 ;
 RECT 5.82 1.535 5.96 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 2.105 0.08 2.245 0.675 ;
 RECT 1.15 0.08 1.29 0.675 ;
 RECT 0.185 0.08 0.325 0.675 ;
 RECT 4.025 0.08 4.165 0.675 ;
 RECT 3.06 0.08 3.2 0.675 ;
 RECT 4.925 0.08 5.065 0.79 ;
 RECT 0 -0.08 6.4 0.08 ;
 RECT 5.805 0.08 5.945 0.795 ;
 END
 END VSS

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.59 0.515 2.73 0.865 ;
 RECT 1.635 0.515 1.775 0.865 ;
 RECT 0.67 0.515 0.81 0.865 ;
 RECT 3.545 1.29 3.685 2.36 ;
 RECT 3.105 1.005 3.685 1.29 ;
 RECT 2.59 1.005 2.73 2.36 ;
 RECT 1.635 1.005 1.775 2.36 ;
 RECT 0.67 1.005 0.81 2.36 ;
 RECT 3.545 0.515 3.685 0.865 ;
 RECT 0.67 0.865 3.685 1.005 ;
 END
 ANTENNADIFFAREA 2.392 ;
 END ZN

 OBS
 LAYER PO ;
 RECT 3.8 1.18 3.9 1.23 ;
 RECT 3.8 1.33 3.9 2.74 ;
 RECT 0.44 1.23 3.9 1.33 ;
 RECT 0.44 0.23 0.54 1.23 ;
 RECT 0.925 0.23 1.025 1.23 ;
 RECT 1.405 0.23 1.505 1.23 ;
 RECT 1.89 0.23 1.99 1.23 ;
 RECT 2.36 0.23 2.46 1.23 ;
 RECT 2.845 0.23 2.945 1.23 ;
 RECT 3.315 0.23 3.415 1.23 ;
 RECT 3.8 0.23 3.9 0.95 ;
 RECT 0.44 1.33 0.54 2.74 ;
 RECT 0.925 1.33 1.025 2.74 ;
 RECT 1.405 1.33 1.505 2.74 ;
 RECT 1.89 1.33 1.99 2.74 ;
 RECT 2.36 1.33 2.46 2.74 ;
 RECT 2.845 1.33 2.945 2.74 ;
 RECT 3.315 1.33 3.415 2.74 ;
 RECT 3.8 0.95 4.055 1.18 ;
 RECT 4.71 0.26 4.81 1.12 ;
 RECT 4.71 1.35 4.81 2.75 ;
 RECT 4.58 1.12 4.81 1.35 ;
 RECT 5.18 0.385 5.28 2.16 ;
 RECT 5.18 2.16 5.41 2.39 ;
 LAYER CO ;
 RECT 5.825 2.105 5.955 2.235 ;
 RECT 5.825 1.845 5.955 1.975 ;
 RECT 3.55 1.645 3.68 1.775 ;
 RECT 5.23 2.21 5.36 2.34 ;
 RECT 5.4 0.605 5.53 0.735 ;
 RECT 4.44 1.705 4.57 1.835 ;
 RECT 4.44 1.705 4.57 1.835 ;
 RECT 4.93 0.605 5.06 0.735 ;
 RECT 5.81 0.615 5.94 0.745 ;
 RECT 5.81 0.355 5.94 0.485 ;
 RECT 3.55 0.565 3.68 0.695 ;
 RECT 3.55 1.95 3.68 2.08 ;
 RECT 5.4 1.75 5.53 1.88 ;
 RECT 4.44 0.605 4.57 0.735 ;
 RECT 5.825 1.585 5.955 1.715 ;
 RECT 3.065 0.495 3.195 0.625 ;
 RECT 4.055 1.96 4.185 2.09 ;
 RECT 3.875 1 4.005 1.13 ;
 RECT 4.93 1.9 5.06 2.03 ;
 RECT 4.03 0.495 4.16 0.625 ;
 RECT 3.55 1.645 3.68 1.775 ;
 RECT 0.675 1.95 0.805 2.08 ;
 RECT 0.675 1.645 0.805 1.775 ;
 RECT 0.675 1.645 0.805 1.775 ;
 RECT 0.19 1.96 0.32 2.09 ;
 RECT 0.19 0.495 0.32 0.625 ;
 RECT 0.675 0.565 0.805 0.695 ;
 RECT 1.64 1.95 1.77 2.08 ;
 RECT 1.64 1.645 1.77 1.775 ;
 RECT 1.64 1.645 1.77 1.775 ;
 RECT 1.155 1.96 1.285 2.09 ;
 RECT 1.155 0.495 1.285 0.625 ;
 RECT 1.64 0.565 1.77 0.695 ;
 RECT 2.595 1.95 2.725 2.08 ;
 RECT 2.595 1.645 2.725 1.775 ;
 RECT 2.595 1.645 2.725 1.775 ;
 RECT 2.11 1.96 2.24 2.09 ;
 RECT 2.11 0.495 2.24 0.625 ;
 RECT 2.595 0.565 2.725 0.695 ;
 RECT 4.63 1.17 4.76 1.3 ;
 RECT 3.065 1.96 3.195 2.09 ;
 LAYER M1 ;
 RECT 4.715 1.085 4.855 1.12 ;
 RECT 4.625 1.12 4.855 1.35 ;
 RECT 4.715 1.35 4.855 1.54 ;
 RECT 5.395 1.68 5.535 1.93 ;
 RECT 5.395 0.555 5.535 1.54 ;
 RECT 4.715 1.54 5.535 1.68 ;
 RECT 3.87 1.09 4.01 1.18 ;
 RECT 3.87 0.95 4.575 0.975 ;
 RECT 3.87 0.975 4.485 1.09 ;
 RECT 4.435 0.515 4.575 0.835 ;
 RECT 4.345 0.835 4.575 0.95 ;
 RECT 4.345 1.09 4.485 1.545 ;
 RECT 4.435 1.685 4.575 1.885 ;
 RECT 4.345 1.545 4.575 1.685 ;
 END
END IBUFFX8

MACRO INVX0
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 1.92 BY 2.88 ;
 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.91 1.12 1.315 1.47 ;
 RECT 0.91 0.555 1.05 1.12 ;
 RECT 0.91 1.47 1.05 1.87 ;
 END
 ANTENNADIFFAREA 0.242 ;
 END ZN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 1.92 2.96 ;
 RECT 1.43 1.985 1.57 2.8 ;
 RECT 0.44 1.64 0.58 2.8 ;
 END
 END VDD

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.36 1.125 0.745 1.46 ;
 END
 ANTENNAGATEAREA 0.079 ;
 END INP

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 1.92 0.08 ;
 RECT 1.43 0.08 1.57 0.83 ;
 RECT 0.44 0.08 0.58 0.785 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.695 0.385 0.795 0.975 ;
 RECT 0.695 0.82 0.795 2.17 ;
 RECT 0.515 1.125 0.745 1.355 ;
 LAYER CO ;
 RECT 1.435 0.64 1.565 0.77 ;
 RECT 1.435 0.37 1.565 0.5 ;
 RECT 1.435 2.305 1.565 2.435 ;
 RECT 1.435 2.035 1.565 2.165 ;
 RECT 0.445 0.605 0.575 0.735 ;
 RECT 0.915 1.69 1.045 1.82 ;
 RECT 0.565 1.175 0.695 1.305 ;
 RECT 0.445 1.69 0.575 1.82 ;
 RECT 0.915 0.605 1.045 0.735 ;
 END
END INVX0

MACRO INVX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.24 BY 2.88 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.325 1.125 0.815 1.465 ;
 END
 ANTENNAGATEAREA 0.161 ;
 END INP

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.99 1.125 1.34 1.475 ;
 RECT 0.99 0.595 1.13 1.125 ;
 RECT 0.99 1.475 1.13 2.435 ;
 END
 ANTENNADIFFAREA 0.499 ;
 END ZN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.24 2.96 ;
 RECT 1.58 1.925 1.72 2.8 ;
 RECT 0.49 1.625 0.63 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.24 0.08 ;
 RECT 1.58 0.08 1.72 0.82 ;
 RECT 0.49 0.08 0.63 0.825 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 0.765 0.275 0.865 0.975 ;
 RECT 0.765 0.82 0.865 2.74 ;
 RECT 0.585 1.125 0.815 1.355 ;
 LAYER CO ;
 RECT 1.585 0.64 1.715 0.77 ;
 RECT 1.585 0.37 1.715 0.5 ;
 RECT 1.585 2.245 1.715 2.375 ;
 RECT 1.585 1.975 1.715 2.105 ;
 RECT 0.995 1.945 1.125 2.075 ;
 RECT 0.995 2.255 1.125 2.385 ;
 RECT 0.495 0.645 0.625 0.775 ;
 RECT 0.635 1.175 0.765 1.305 ;
 RECT 0.995 1.685 1.125 1.815 ;
 RECT 0.495 2.255 0.625 2.385 ;
 RECT 0.495 1.945 0.625 2.075 ;
 RECT 0.495 1.675 0.625 1.805 ;
 RECT 0.995 0.645 1.125 0.775 ;
 END
END INVX1

MACRO TNBUFFX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.32 BY 2.88 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.105 1.155 1.715 1.405 ;
 END
 ANTENNAGATEAREA 0.191 ;
 END ENB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.32 2.96 ;
 RECT 1.26 2.05 1.4 2.8 ;
 RECT 2.405 2.355 2.545 2.8 ;
 RECT 4.055 2.37 4.195 2.8 ;
 RECT 7.82 2.36 7.96 2.8 ;
 RECT 6.88 2.37 7.02 2.8 ;
 RECT 5.94 2.37 6.08 2.8 ;
 RECT 5 2.37 5.14 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.32 0.08 ;
 RECT 4.935 0.305 5.21 0.445 ;
 RECT 5.88 0.305 6.155 0.445 ;
 RECT 6.82 0.305 7.095 0.445 ;
 RECT 7.76 0.305 8.035 0.445 ;
 RECT 2.685 0.815 3.3 0.955 ;
 RECT 1.26 0.08 1.4 0.825 ;
 RECT 4.055 0.08 4.195 0.7 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 5 0.08 5.14 0.305 ;
 RECT 5.945 0.08 6.085 0.305 ;
 RECT 6.885 0.08 7.025 0.305 ;
 RECT 7.825 0.08 7.965 0.305 ;
 RECT 3.16 0.08 3.3 0.815 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.37 0.225 3.02 0.445 ;
 RECT 2.72 0.445 3.02 0.645 ;
 END
 ANTENNAGATEAREA 0.145 ;
 END INP

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.105 0.725 8.245 2.045 ;
 RECT 7.295 2.185 7.645 2.425 ;
 RECT 7.295 2.18 8.245 2.185 ;
 RECT 4.47 2.045 8.245 2.18 ;
 RECT 4.455 0.585 8.245 0.725 ;
 RECT 4.47 2.04 7.645 2.045 ;
 END
 ANTENNADIFFAREA 2.426 ;
 END Z

 OBS
 LAYER PO ;
 RECT 3.01 1.205 3.11 1.61 ;
 RECT 2.985 0.495 3.085 1.105 ;
 RECT 3.01 1.61 3.28 1.84 ;
 RECT 3.01 1.84 3.11 2.79 ;
 RECT 2.985 1.105 3.11 1.205 ;
 RECT 4.785 0.09 4.885 0.84 ;
 RECT 4.705 0.97 4.915 1.09 ;
 RECT 7.61 0.09 7.71 0.84 ;
 RECT 7.14 0.09 7.24 0.84 ;
 RECT 6.67 0.09 6.77 0.84 ;
 RECT 6.2 0.09 6.3 0.84 ;
 RECT 5.73 0.09 5.83 0.84 ;
 RECT 5.255 0.09 5.355 0.84 ;
 RECT 4.315 0.84 7.71 0.97 ;
 RECT 4.315 0.09 4.415 0.84 ;
 RECT 6.77 0.97 6.98 1.09 ;
 RECT 2.405 0.41 2.505 1.09 ;
 RECT 2.185 1.205 2.285 2.79 ;
 RECT 2.185 1.09 2.505 1.205 ;
 RECT 2.405 0.18 2.615 0.41 ;
 RECT 1.875 0.28 1.975 1.68 ;
 RECT 1.045 1.385 1.145 1.68 ;
 RECT 1.045 1.78 1.145 2.58 ;
 RECT 1.515 1.78 1.615 2.78 ;
 RECT 1.045 0.4 1.145 1.155 ;
 RECT 1.045 1.155 1.29 1.385 ;
 RECT 1.045 1.68 1.975 1.78 ;
 RECT 3.46 1.44 3.91 1.655 ;
 RECT 4.315 1.44 4.415 2.79 ;
 RECT 7.605 1.44 7.705 2.79 ;
 RECT 7.135 1.44 7.235 2.79 ;
 RECT 6.665 1.44 6.765 2.79 ;
 RECT 6.195 1.44 6.295 2.79 ;
 RECT 5.725 1.44 5.825 2.79 ;
 RECT 5.255 1.44 5.355 2.79 ;
 RECT 4.785 1.44 4.885 2.79 ;
 RECT 7.79 1.19 8 1.31 ;
 RECT 5.91 1.19 6.12 1.31 ;
 RECT 4.315 1.19 4.525 1.31 ;
 RECT 3.46 1.425 8 1.44 ;
 RECT 3.6 1.31 8 1.425 ;
 LAYER CO ;
 RECT 3.5 1.475 3.63 1.605 ;
 RECT 2.445 0.23 2.575 0.36 ;
 RECT 3.11 1.66 3.24 1.79 ;
 RECT 3.235 2.405 3.365 2.535 ;
 RECT 3.445 0.845 3.575 0.975 ;
 RECT 2.76 2.08 2.89 2.21 ;
 RECT 2.41 2.405 2.54 2.535 ;
 RECT 1.625 0.78 1.755 0.91 ;
 RECT 2.095 0.535 2.225 0.665 ;
 RECT 1.845 2.08 1.975 2.21 ;
 RECT 1.265 2.12 1.395 2.25 ;
 RECT 1.265 0.625 1.395 0.755 ;
 RECT 0.795 0.625 0.925 0.755 ;
 RECT 0.795 2.12 0.925 2.25 ;
 RECT 4.745 0.91 4.875 1.04 ;
 RECT 7.83 1.24 7.96 1.37 ;
 RECT 5.95 1.24 6.08 1.37 ;
 RECT 6.81 0.91 6.94 1.04 ;
 RECT 4.355 1.24 4.485 1.37 ;
 RECT 6.89 0.31 7.02 0.44 ;
 RECT 7.83 0.31 7.96 0.44 ;
 RECT 6.42 0.59 6.55 0.72 ;
 RECT 5.95 0.31 6.08 0.44 ;
 RECT 5.475 0.59 5.605 0.72 ;
 RECT 5.005 0.31 5.135 0.44 ;
 RECT 4.535 0.59 4.665 0.72 ;
 RECT 7.36 0.59 7.49 0.72 ;
 RECT 7.355 2.045 7.485 2.175 ;
 RECT 6.885 2.44 7.015 2.57 ;
 RECT 6.415 2.045 6.545 2.175 ;
 RECT 5.475 2.045 5.605 2.175 ;
 RECT 5.005 2.44 5.135 2.57 ;
 RECT 4.535 2.045 4.665 2.175 ;
 RECT 7.825 2.43 7.955 2.56 ;
 RECT 5.945 2.44 6.075 2.57 ;
 RECT 4.06 0.5 4.19 0.63 ;
 RECT 4.06 2.44 4.19 2.57 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 2.735 0.82 2.865 0.95 ;
 RECT 1.12 1.205 1.25 1.335 ;
 LAYER M1 ;
 RECT 5.945 1.18 6.085 1.645 ;
 RECT 7.825 1.18 7.965 1.645 ;
 RECT 4.35 1.19 4.49 1.645 ;
 RECT 4.35 1.645 7.965 1.785 ;
 RECT 0.79 1.555 1.835 1.655 ;
 RECT 0.79 0.555 0.93 1.555 ;
 RECT 0.79 1.695 0.93 2.32 ;
 RECT 1.695 1.695 3.31 1.795 ;
 RECT 0.79 1.655 3.31 1.695 ;
 RECT 2.09 1.015 2.23 1.375 ;
 RECT 1.62 0.71 1.76 0.875 ;
 RECT 1.62 0.875 2.23 1.015 ;
 RECT 3.495 1.515 3.635 2.075 ;
 RECT 2.09 1.375 3.635 1.515 ;
 RECT 1.665 2.075 3.635 2.215 ;
 RECT 3.44 0.775 3.58 0.865 ;
 RECT 3.44 1.005 3.915 1.095 ;
 RECT 2.37 1.095 3.915 1.235 ;
 RECT 3.775 1.235 3.915 2.4 ;
 RECT 3.165 2.4 3.915 2.54 ;
 RECT 2.09 0.595 2.545 0.735 ;
 RECT 2.405 0.735 2.545 1.095 ;
 RECT 2.09 0.46 2.23 0.595 ;
 RECT 4.695 1.005 4.925 1.045 ;
 RECT 3.44 0.865 6.99 1.005 ;
 RECT 6.76 1.005 6.99 1.045 ;
 END
END TNBUFFX8

MACRO XNOR2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 0.665 0.08 0.805 0.775 ;
 RECT 2.075 0.08 2.215 0.82 ;
 RECT 3.9 0.08 4.04 0.82 ;
 RECT 0.215 0.08 0.355 0.755 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.28 1.32 3.64 1.56 ;
 END
 ANTENNAGATEAREA 0.134 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.66 0.985 1 1.4 ;
 END
 ANTENNAGATEAREA 0.134 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.36 0.36 4.6 0.6 ;
 RECT 4.45 1.16 4.715 1.4 ;
 RECT 4.45 1.4 4.59 2.565 ;
 RECT 4.45 0.6 4.59 1.16 ;
 END
 ANTENNADIFFAREA 0.567 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 0.665 1.55 0.805 2.8 ;
 RECT 2.09 1.825 2.23 2.8 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 3.88 2.12 4.02 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 3.665 0.39 3.765 2.425 ;
 RECT 3.56 2.425 3.77 2.655 ;
 RECT 2.775 1.665 2.875 2.53 ;
 RECT 2.66 1.45 2.89 1.665 ;
 RECT 3.28 0.425 3.38 0.975 ;
 RECT 3.16 0.21 3.39 0.425 ;
 RECT 0.92 2.44 2.47 2.535 ;
 RECT 0.92 2.535 2.465 2.54 ;
 RECT 2.37 0.395 2.47 2.44 ;
 RECT 0.92 1.215 1.02 2.44 ;
 RECT 0.92 0.375 1.02 0.985 ;
 RECT 0.815 0.985 1.025 1.215 ;
 RECT 3.28 1.56 3.38 2.53 ;
 RECT 1.785 0.215 1.885 2.255 ;
 RECT 2.77 0.215 2.87 1.165 ;
 RECT 3.27 1.265 3.485 1.56 ;
 RECT 2.77 1.165 3.38 1.265 ;
 RECT 1.785 0.115 2.87 0.215 ;
 RECT 4.17 0.35 4.27 1.07 ;
 RECT 4.17 1.285 4.27 2.745 ;
 RECT 4.045 1.07 4.275 1.285 ;
 LAYER CO ;
 RECT 2.71 1.49 2.84 1.62 ;
 RECT 0.855 1.035 0.985 1.165 ;
 RECT 1.535 1.81 1.665 1.94 ;
 RECT 0.67 1.62 0.8 1.75 ;
 RECT 3.885 2.17 4.015 2.3 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 2.995 1.81 3.125 1.94 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 3.6 2.475 3.73 2.605 ;
 RECT 1.145 0.595 1.275 0.725 ;
 RECT 3.905 0.625 4.035 0.755 ;
 RECT 3.21 0.25 3.34 0.38 ;
 RECT 1.535 0.625 1.665 0.755 ;
 RECT 2.08 0.625 2.21 0.755 ;
 RECT 4.455 1.56 4.585 1.69 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 2.095 1.875 2.225 2.005 ;
 RECT 1.145 1.6 1.275 1.73 ;
 RECT 4.455 2.385 4.585 2.515 ;
 RECT 4.455 2.11 4.585 2.24 ;
 RECT 4.455 1.835 4.585 1.965 ;
 RECT 2.995 0.625 3.125 0.755 ;
 RECT 2.995 2.115 3.125 2.245 ;
 RECT 4.095 1.11 4.225 1.24 ;
 RECT 3.315 1.38 3.445 1.51 ;
 RECT 0.67 0.595 0.8 0.725 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 4.455 0.625 4.585 0.755 ;
 LAYER M1 ;
 RECT 1.14 0.48 1.28 2.235 ;
 RECT 1.14 2.235 1.95 2.375 ;
 RECT 1.81 1.645 1.95 2.235 ;
 RECT 1.81 1.505 2.52 1.645 ;
 RECT 2.38 1.645 2.52 2.475 ;
 RECT 3.59 2.425 3.74 2.475 ;
 RECT 3.59 2.615 3.74 2.655 ;
 RECT 2.38 2.475 3.74 2.615 ;
 RECT 1.53 0.3 1.67 0.97 ;
 RECT 1.53 1.11 1.67 1.99 ;
 RECT 2.705 0.385 2.845 0.97 ;
 RECT 2.705 1.11 2.845 1.44 ;
 RECT 1.53 0.97 2.845 1.11 ;
 RECT 2.7 1.44 2.85 1.675 ;
 RECT 2.705 0.245 3.39 0.385 ;
 RECT 2.99 0.535 3.13 0.625 ;
 RECT 2.99 0.765 3.13 2.295 ;
 RECT 2.99 0.625 3.745 0.765 ;
 RECT 3.605 0.765 3.745 1.02 ;
 RECT 4.085 1.16 4.235 1.295 ;
 RECT 3.605 1.02 4.27 1.16 ;
 END
END XNOR2X1

MACRO INVX32
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 16.32 BY 2.88 ;
 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 15.26 2 15.4 2.04 ;
 RECT 14.32 2 14.46 2.31 ;
 RECT 13.38 2 13.52 2.31 ;
 RECT 12.44 2 12.58 2.31 ;
 RECT 11.5 2 11.64 2.31 ;
 RECT 10.56 2 10.7 2.31 ;
 RECT 9.62 2 9.76 2.31 ;
 RECT 8.68 2 8.82 2.31 ;
 RECT 3.98 2 4.12 2.31 ;
 RECT 7.74 2 7.88 2.31 ;
 RECT 6.8 2 6.94 2.31 ;
 RECT 5.86 2 6 2.31 ;
 RECT 4.92 2 5.06 2.31 ;
 RECT 3.04 2 3.18 2.31 ;
 RECT 2.1 2 2.24 2.31 ;
 RECT 1.16 2 1.3 2.31 ;
 RECT 14.32 1.86 15.4 2 ;
 RECT 12.44 1.86 13.52 2 ;
 RECT 10.56 1.86 11.64 2 ;
 RECT 8.68 1.86 9.76 2 ;
 RECT 3.04 1.86 4.12 2 ;
 RECT 6.8 1.86 7.88 2 ;
 RECT 4.92 1.86 6 2 ;
 RECT 1.16 1.86 2.24 2 ;
 RECT 14.32 1.855 14.46 1.86 ;
 RECT 12.44 1.855 12.58 1.86 ;
 RECT 13.38 1.855 13.52 1.86 ;
 RECT 10.56 1.855 10.7 1.86 ;
 RECT 8.68 1.855 8.82 1.86 ;
 RECT 11.5 1.855 11.64 1.86 ;
 RECT 9.62 1.855 9.76 1.86 ;
 RECT 3.98 1.855 4.12 1.86 ;
 RECT 6.8 1.855 6.94 1.86 ;
 RECT 4.92 1.855 5.06 1.86 ;
 RECT 7.74 1.855 7.88 1.86 ;
 RECT 5.86 1.855 6 1.86 ;
 RECT 0.22 1.855 0.36 2.31 ;
 RECT 3.04 1.855 3.18 1.86 ;
 RECT 1.16 1.855 1.3 1.86 ;
 RECT 2.1 1.855 2.24 1.86 ;
 RECT 7.74 1.715 8.82 1.855 ;
 RECT 11.5 1.715 12.58 1.855 ;
 RECT 13.38 1.715 14.46 1.855 ;
 RECT 13.38 1.585 13.52 1.715 ;
 RECT 11.5 1.585 11.64 1.715 ;
 RECT 9.62 1.715 10.7 1.855 ;
 RECT 9.62 1.585 9.76 1.715 ;
 RECT 3.98 1.715 5.06 1.855 ;
 RECT 3.98 1.585 4.12 1.715 ;
 RECT 7.74 1.585 7.88 1.715 ;
 RECT 5.86 1.715 6.94 1.855 ;
 RECT 5.86 1.585 6 1.715 ;
 RECT 2.1 1.715 3.18 1.855 ;
 RECT 2.1 1.585 2.24 1.715 ;
 RECT 0.22 1.715 1.3 1.855 ;
 RECT 15.26 1.435 15.4 1.86 ;
 RECT 15.26 1.125 15.725 1.435 ;
 RECT 15.26 1.08 15.4 1.125 ;
 RECT 0.22 0.94 15.4 1.08 ;
 RECT 6.8 0.625 6.94 0.94 ;
 RECT 4.92 0.625 5.06 0.94 ;
 RECT 3.04 0.625 3.18 0.94 ;
 RECT 1.16 0.625 1.3 0.94 ;
 RECT 7.74 0.64 7.88 0.94 ;
 RECT 5.86 0.64 6 0.94 ;
 RECT 3.98 0.64 4.12 0.94 ;
 RECT 2.1 0.64 2.24 0.94 ;
 RECT 0.22 0.64 0.36 0.94 ;
 RECT 10.56 0.625 10.7 0.94 ;
 RECT 8.68 0.625 8.82 0.94 ;
 RECT 11.5 0.64 11.64 0.94 ;
 RECT 9.62 0.64 9.76 0.94 ;
 RECT 15.26 0.64 15.4 0.94 ;
 RECT 14.32 0.625 14.46 0.94 ;
 RECT 12.44 0.625 12.58 0.94 ;
 RECT 13.38 0.64 13.52 0.94 ;
 END
 ANTENNADIFFAREA 9.906 ;
 END ZN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 16.32 2.96 ;
 RECT 15.77 1.965 15.91 2.8 ;
 RECT 9.15 2.345 9.29 2.8 ;
 RECT 11.03 2.345 11.17 2.8 ;
 RECT 12.91 2.345 13.05 2.8 ;
 RECT 14.79 2.345 14.93 2.8 ;
 RECT 8.21 2.065 8.35 2.8 ;
 RECT 10.09 2.065 10.23 2.8 ;
 RECT 11.97 2.065 12.11 2.8 ;
 RECT 13.85 2.065 13.99 2.8 ;
 RECT 5.39 2.345 5.53 2.8 ;
 RECT 7.27 2.345 7.41 2.8 ;
 RECT 3.51 2.345 3.65 2.8 ;
 RECT 1.63 2.345 1.77 2.8 ;
 RECT 6.33 2.065 6.47 2.8 ;
 RECT 4.45 2.065 4.59 2.8 ;
 RECT 2.57 2.065 2.71 2.8 ;
 RECT 0.69 2.065 0.83 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 16.32 0.08 ;
 RECT 15.77 0.08 15.91 0.8 ;
 RECT 8.21 0.08 8.35 0.77 ;
 RECT 9.15 0.08 9.29 0.77 ;
 RECT 10.09 0.08 10.23 0.77 ;
 RECT 11.03 0.08 11.17 0.77 ;
 RECT 11.97 0.08 12.11 0.77 ;
 RECT 12.91 0.08 13.05 0.77 ;
 RECT 13.85 0.08 13.99 0.77 ;
 RECT 14.79 0.08 14.93 0.77 ;
 RECT 6.33 0.08 6.47 0.77 ;
 RECT 5.39 0.08 5.53 0.77 ;
 RECT 7.27 0.08 7.41 0.77 ;
 RECT 4.45 0.08 4.59 0.77 ;
 RECT 3.51 0.08 3.65 0.77 ;
 RECT 2.57 0.08 2.71 0.77 ;
 RECT 1.63 0.08 1.77 0.77 ;
 RECT 0.69 0.08 0.83 0.77 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.665 1.37 15.01 1.72 ;
 RECT 0.41 1.23 15.12 1.37 ;
 END
 ANTENNAGATEAREA 5.152 ;
 END INP

 OBS
 LAYER PO ;
 RECT 13.165 0.275 13.265 1.185 ;
 RECT 13.01 1.185 13.265 1.415 ;
 RECT 13.165 1.415 13.265 2.79 ;
 RECT 8.465 0.275 8.565 1.185 ;
 RECT 8.465 1.415 8.565 2.79 ;
 RECT 8.38 1.185 8.61 1.415 ;
 RECT 10.345 0.275 10.445 1.185 ;
 RECT 10.345 1.415 10.445 2.79 ;
 RECT 10.31 1.185 10.54 1.415 ;
 RECT 7.525 0.275 7.625 1.185 ;
 RECT 7.37 1.185 7.625 1.415 ;
 RECT 7.525 1.415 7.625 2.79 ;
 RECT 2.355 0.275 2.455 1.185 ;
 RECT 2.355 1.185 2.61 1.415 ;
 RECT 2.355 1.415 2.455 2.79 ;
 RECT 14.105 0.275 14.205 1.185 ;
 RECT 14.105 1.415 14.205 2.79 ;
 RECT 14.07 1.185 14.3 1.415 ;
 RECT 7.055 0.275 7.155 1.185 ;
 RECT 7.055 1.415 7.155 2.79 ;
 RECT 6.96 1.185 7.19 1.415 ;
 RECT 0.945 0.275 1.045 1.185 ;
 RECT 0.945 1.415 1.045 2.79 ;
 RECT 0.86 1.185 1.09 1.415 ;
 RECT 9.405 0.275 9.505 1.185 ;
 RECT 9.25 1.185 9.505 1.415 ;
 RECT 9.405 1.415 9.505 2.79 ;
 RECT 12.695 0.275 12.795 1.185 ;
 RECT 12.695 1.415 12.795 2.79 ;
 RECT 12.585 1.185 12.815 1.415 ;
 RECT 8.935 0.275 9.035 1.185 ;
 RECT 8.935 1.415 9.035 2.79 ;
 RECT 8.825 1.185 9.055 1.415 ;
 RECT 11.755 1.185 12.37 1.415 ;
 RECT 12.225 0.275 12.325 1.185 ;
 RECT 12.225 1.415 12.325 2.79 ;
 RECT 11.755 0.275 11.855 1.185 ;
 RECT 11.755 1.415 11.855 2.79 ;
 RECT 15.045 0.275 15.145 1.185 ;
 RECT 14.89 1.185 15.145 1.415 ;
 RECT 15.045 1.415 15.145 2.79 ;
 RECT 11.285 0.275 11.385 1.185 ;
 RECT 11.13 1.185 11.385 1.415 ;
 RECT 11.285 1.415 11.385 2.79 ;
 RECT 14.575 0.275 14.675 1.185 ;
 RECT 14.575 1.415 14.675 2.79 ;
 RECT 14.48 1.185 14.71 1.415 ;
 RECT 13.635 0.275 13.735 1.185 ;
 RECT 13.635 1.185 13.89 1.415 ;
 RECT 13.635 1.415 13.735 2.79 ;
 RECT 9.875 0.275 9.975 1.185 ;
 RECT 9.875 1.185 10.13 1.415 ;
 RECT 9.875 1.415 9.975 2.79 ;
 RECT 6.115 0.275 6.215 1.185 ;
 RECT 6.115 1.185 6.37 1.415 ;
 RECT 6.115 1.415 6.215 2.79 ;
 RECT 3.765 0.275 3.865 1.185 ;
 RECT 3.61 1.185 3.865 1.415 ;
 RECT 3.765 1.415 3.865 2.79 ;
 RECT 3.295 0.275 3.395 1.185 ;
 RECT 3.295 1.415 3.395 2.79 ;
 RECT 3.2 1.185 3.43 1.415 ;
 RECT 2.825 0.275 2.925 1.185 ;
 RECT 2.825 1.415 2.925 2.79 ;
 RECT 2.79 1.185 3.02 1.415 ;
 RECT 10.815 0.275 10.915 1.185 ;
 RECT 10.815 1.415 10.915 2.79 ;
 RECT 10.72 1.185 10.95 1.415 ;
 RECT 1.885 0.275 1.985 1.185 ;
 RECT 1.73 1.185 1.985 1.415 ;
 RECT 1.885 1.415 1.985 2.79 ;
 RECT 1.415 0.275 1.515 1.185 ;
 RECT 1.415 1.415 1.515 2.79 ;
 RECT 1.305 1.185 1.535 1.415 ;
 RECT 7.995 0.275 8.095 1.185 ;
 RECT 7.995 1.415 8.095 2.79 ;
 RECT 7.93 1.185 8.16 1.415 ;
 RECT 0.475 0.275 0.575 1.185 ;
 RECT 0.475 1.415 0.575 2.79 ;
 RECT 0.41 1.185 0.64 1.415 ;
 RECT 5.645 0.275 5.745 1.185 ;
 RECT 5.49 1.185 5.745 1.415 ;
 RECT 5.645 1.415 5.745 2.79 ;
 RECT 5.175 0.275 5.275 1.185 ;
 RECT 5.175 1.415 5.275 2.79 ;
 RECT 5.065 1.185 5.295 1.415 ;
 RECT 4.235 1.185 4.85 1.415 ;
 RECT 4.705 0.275 4.805 1.185 ;
 RECT 4.705 1.415 4.805 2.79 ;
 RECT 4.235 0.275 4.335 1.185 ;
 RECT 4.235 1.415 4.335 2.79 ;
 RECT 6.585 0.275 6.685 1.185 ;
 RECT 6.585 1.415 6.685 2.79 ;
 RECT 6.55 1.185 6.78 1.415 ;
 LAYER CO ;
 RECT 9.155 2.44 9.285 2.57 ;
 RECT 14.795 0.59 14.925 0.72 ;
 RECT 3.66 1.235 3.79 1.365 ;
 RECT 3.25 1.235 3.38 1.365 ;
 RECT 2.84 1.235 2.97 1.365 ;
 RECT 10.77 1.235 10.9 1.365 ;
 RECT 15.775 2.285 15.905 2.415 ;
 RECT 5.395 2.44 5.525 2.57 ;
 RECT 5.395 0.59 5.525 0.72 ;
 RECT 0.46 1.235 0.59 1.365 ;
 RECT 0.91 1.235 1.04 1.365 ;
 RECT 7.98 1.235 8.11 1.365 ;
 RECT 0.225 1.86 0.355 1.99 ;
 RECT 0.695 2.115 0.825 2.245 ;
 RECT 2.105 0.69 2.235 0.82 ;
 RECT 0.225 0.69 0.355 0.82 ;
 RECT 7.275 0.59 7.405 0.72 ;
 RECT 6.335 0.59 6.465 0.72 ;
 RECT 14.325 2.13 14.455 2.26 ;
 RECT 11.975 2.425 12.105 2.555 ;
 RECT 14.325 1.86 14.455 1.99 ;
 RECT 9.155 0.59 9.285 0.72 ;
 RECT 8.215 2.425 8.345 2.555 ;
 RECT 5.54 1.235 5.67 1.365 ;
 RECT 5.115 1.235 5.245 1.365 ;
 RECT 9.625 1.86 9.755 1.99 ;
 RECT 8.215 2.115 8.345 2.245 ;
 RECT 13.385 0.69 13.515 0.82 ;
 RECT 11.505 1.86 11.635 1.99 ;
 RECT 12.445 1.86 12.575 1.99 ;
 RECT 6.6 1.235 6.73 1.365 ;
 RECT 3.045 1.86 3.175 1.99 ;
 RECT 2.575 0.59 2.705 0.72 ;
 RECT 15.265 1.86 15.395 1.99 ;
 RECT 13.385 1.86 13.515 1.99 ;
 RECT 12.445 0.675 12.575 0.805 ;
 RECT 5.865 2.13 5.995 2.26 ;
 RECT 5.865 0.69 5.995 0.82 ;
 RECT 0.695 0.59 0.825 0.72 ;
 RECT 13.06 1.235 13.19 1.365 ;
 RECT 8.215 0.59 8.345 0.72 ;
 RECT 7.745 2.13 7.875 2.26 ;
 RECT 11.975 0.59 12.105 0.72 ;
 RECT 11.035 2.44 11.165 2.57 ;
 RECT 12.19 1.235 12.32 1.365 ;
 RECT 2.105 1.86 2.235 1.99 ;
 RECT 2.105 0.69 2.235 0.82 ;
 RECT 6.805 0.675 6.935 0.805 ;
 RECT 7.745 1.86 7.875 1.99 ;
 RECT 4.925 1.86 5.055 1.99 ;
 RECT 9.625 0.69 9.755 0.82 ;
 RECT 10.565 2.13 10.695 2.26 ;
 RECT 12.445 2.13 12.575 2.26 ;
 RECT 15.775 0.62 15.905 0.75 ;
 RECT 1.635 0.59 1.765 0.72 ;
 RECT 8.685 0.675 8.815 0.805 ;
 RECT 6.335 2.425 6.465 2.555 ;
 RECT 5.865 1.86 5.995 1.99 ;
 RECT 10.36 1.235 10.49 1.365 ;
 RECT 7.42 1.235 7.55 1.365 ;
 RECT 1.78 1.235 1.91 1.365 ;
 RECT 2.105 1.86 2.235 1.99 ;
 RECT 12.915 0.59 13.045 0.72 ;
 RECT 13.385 1.86 13.515 1.99 ;
 RECT 10.565 1.86 10.695 1.99 ;
 RECT 6.805 1.86 6.935 1.99 ;
 RECT 5.865 1.86 5.995 1.99 ;
 RECT 7.745 0.69 7.875 0.82 ;
 RECT 9.625 1.86 9.755 1.99 ;
 RECT 8.43 1.235 8.56 1.365 ;
 RECT 11.83 1.235 11.96 1.365 ;
 RECT 3.985 1.86 4.115 1.99 ;
 RECT 2.575 2.115 2.705 2.245 ;
 RECT 3.045 2.13 3.175 2.26 ;
 RECT 4.455 0.59 4.585 0.72 ;
 RECT 3.985 2.13 4.115 2.26 ;
 RECT 7.275 2.44 7.405 2.57 ;
 RECT 6.335 2.115 6.465 2.245 ;
 RECT 2.43 1.235 2.56 1.365 ;
 RECT 8.685 2.13 8.815 2.26 ;
 RECT 15.775 2.015 15.905 2.145 ;
 RECT 4.455 2.425 4.585 2.555 ;
 RECT 13.385 2.13 13.515 2.26 ;
 RECT 12.915 2.44 13.045 2.57 ;
 RECT 11.505 2.13 11.635 2.26 ;
 RECT 11.505 1.86 11.635 1.99 ;
 RECT 10.095 2.115 10.225 2.245 ;
 RECT 11.975 2.115 12.105 2.245 ;
 RECT 1.165 1.86 1.295 1.99 ;
 RECT 1.355 1.235 1.485 1.365 ;
 RECT 13.855 0.59 13.985 0.72 ;
 RECT 14.795 2.44 14.925 2.57 ;
 RECT 13.385 0.69 13.515 0.82 ;
 RECT 1.165 2.13 1.295 2.26 ;
 RECT 1.165 0.675 1.295 0.805 ;
 RECT 3.985 1.86 4.115 1.99 ;
 RECT 3.985 0.69 4.115 0.82 ;
 RECT 14.12 1.235 14.25 1.365 ;
 RECT 11.505 0.69 11.635 0.82 ;
 RECT 15.265 0.69 15.395 0.82 ;
 RECT 9.625 0.69 9.755 0.82 ;
 RECT 11.035 0.59 11.165 0.72 ;
 RECT 7.745 1.86 7.875 1.99 ;
 RECT 7.745 0.69 7.875 0.82 ;
 RECT 10.095 2.425 10.225 2.555 ;
 RECT 10.095 0.59 10.225 0.72 ;
 RECT 10.565 0.675 10.695 0.805 ;
 RECT 7.01 1.235 7.14 1.365 ;
 RECT 0.695 2.425 0.825 2.555 ;
 RECT 9.3 1.235 9.43 1.365 ;
 RECT 12.635 1.235 12.765 1.365 ;
 RECT 8.875 1.235 9.005 1.365 ;
 RECT 3.515 2.44 3.645 2.57 ;
 RECT 3.515 0.59 3.645 0.72 ;
 RECT 2.575 2.425 2.705 2.555 ;
 RECT 11.505 0.69 11.635 0.82 ;
 RECT 9.625 2.13 9.755 2.26 ;
 RECT 14.94 1.235 15.07 1.365 ;
 RECT 11.18 1.235 11.31 1.365 ;
 RECT 14.53 1.235 14.66 1.365 ;
 RECT 15.775 0.35 15.905 0.48 ;
 RECT 6.805 2.13 6.935 2.26 ;
 RECT 4.925 0.675 5.055 0.805 ;
 RECT 4.455 2.115 4.585 2.245 ;
 RECT 4.925 2.13 5.055 2.26 ;
 RECT 13.71 1.235 13.84 1.365 ;
 RECT 9.95 1.235 10.08 1.365 ;
 RECT 4.67 1.235 4.8 1.365 ;
 RECT 4.31 1.235 4.44 1.365 ;
 RECT 0.225 2.13 0.355 2.26 ;
 RECT 1.635 2.44 1.765 2.57 ;
 RECT 8.685 1.86 8.815 1.99 ;
 RECT 6.19 1.235 6.32 1.365 ;
 RECT 2.105 2.13 2.235 2.26 ;
 RECT 3.985 0.69 4.115 0.82 ;
 RECT 3.045 0.675 3.175 0.805 ;
 RECT 5.865 0.69 5.995 0.82 ;
 RECT 14.325 0.675 14.455 0.805 ;
 RECT 13.855 2.425 13.985 2.555 ;
 RECT 13.855 2.115 13.985 2.245 ;
 END
END INVX32

MACRO INVX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 2.605 0.08 2.745 0.805 ;
 RECT 1.525 0.08 1.665 0.77 ;
 RECT 0.585 0.08 0.725 0.77 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.275 1.655 1.575 1.72 ;
 RECT 0.3 1.37 1.575 1.655 ;
 RECT 0.305 1.23 1.855 1.3 ;
 RECT 0.3 1.3 1.855 1.37 ;
 END
 ANTENNAGATEAREA 0.644 ;
 END INP

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.995 1.1 2.62 1.48 ;
 RECT 0.115 0.94 2.135 1.08 ;
 RECT 1.995 1.48 2.135 1.86 ;
 RECT 1.055 0.625 1.195 0.94 ;
 RECT 1.995 1.08 2.135 1.1 ;
 RECT 1.995 0.64 2.135 0.94 ;
 RECT 1.995 2 2.135 2.11 ;
 RECT 0.115 1.86 2.135 2 ;
 RECT 0.115 0.64 0.255 0.94 ;
 RECT 1.055 2 1.195 2.38 ;
 RECT 0.115 2 0.255 2.38 ;
 END
 ANTENNADIFFAREA 1.562 ;
 END ZN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.525 2.345 1.665 2.8 ;
 RECT 2.605 1.975 2.745 2.8 ;
 RECT 0.585 2.305 0.725 2.8 ;
 RECT 0 2.8 3.2 2.96 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.84 0.275 0.94 1.185 ;
 RECT 0.84 1.415 0.94 2.79 ;
 RECT 0.755 1.185 0.985 1.415 ;
 RECT 1.78 0.275 1.88 1.185 ;
 RECT 1.625 1.185 1.88 1.415 ;
 RECT 1.78 1.415 1.88 2.79 ;
 RECT 1.31 0.275 1.41 1.185 ;
 RECT 1.31 1.415 1.41 2.79 ;
 RECT 1.2 1.185 1.43 1.415 ;
 RECT 0.37 0.275 0.47 1.185 ;
 RECT 0.37 1.415 0.47 2.79 ;
 RECT 0.305 1.185 0.535 1.415 ;
 LAYER CO ;
 RECT 2.61 0.625 2.74 0.755 ;
 RECT 2.61 2.025 2.74 2.155 ;
 RECT 2.61 2.295 2.74 2.425 ;
 RECT 2.61 0.355 2.74 0.485 ;
 RECT 0.59 0.59 0.72 0.72 ;
 RECT 0.59 2.425 0.72 2.555 ;
 RECT 0.355 1.235 0.485 1.365 ;
 RECT 0.805 1.235 0.935 1.365 ;
 RECT 0.12 2.2 0.25 2.33 ;
 RECT 1.53 2.44 1.66 2.57 ;
 RECT 1.675 1.235 1.805 1.365 ;
 RECT 2 1.93 2.13 2.06 ;
 RECT 1.06 1.93 1.19 2.06 ;
 RECT 1.25 1.235 1.38 1.365 ;
 RECT 0.12 1.93 0.25 2.06 ;
 RECT 2 0.69 2.13 0.82 ;
 RECT 0.12 0.69 0.25 0.82 ;
 RECT 1.06 2.2 1.19 2.33 ;
 RECT 1.06 0.675 1.19 0.805 ;
 RECT 1.53 0.59 1.66 0.72 ;
 END
END INVX4

MACRO INVX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 1.525 0.08 1.665 0.77 ;
 RECT 2.465 0.08 2.605 0.77 ;
 RECT 0.585 0.08 0.725 0.77 ;
 RECT 3.405 0.08 3.545 0.77 ;
 RECT 4.5 0.08 4.64 0.835 ;
 RECT 0 -0.08 5.12 0.08 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.195 1.37 3.535 1.76 ;
 RECT 0.305 1.23 3.735 1.37 ;
 END
 ANTENNAGATEAREA 1.288 ;
 END INP

 PIN ZN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.875 1.13 4.14 1.44 ;
 RECT 1.055 1.935 1.195 1.985 ;
 RECT 0.115 2.125 0.255 2.435 ;
 RECT 0.115 1.985 4.06 2.125 ;
 RECT 0.115 1.935 0.255 1.985 ;
 RECT 2.935 0.625 3.075 0.94 ;
 RECT 0.115 0.94 4.015 1.08 ;
 RECT 1.055 2.125 1.195 2.435 ;
 RECT 1.995 0.64 2.135 0.94 ;
 RECT 1.055 0.625 1.195 0.94 ;
 RECT 0.115 0.64 0.255 0.94 ;
 RECT 3.875 1.44 4.015 1.985 ;
 RECT 3.875 1.08 4.015 1.13 ;
 RECT 3.875 0.58 4.015 0.94 ;
 RECT 1.995 2.125 2.135 2.435 ;
 RECT 1.995 1.935 2.135 1.985 ;
 RECT 2.935 2.125 3.075 2.435 ;
 RECT 2.935 1.935 3.075 1.985 ;
 END
 ANTENNADIFFAREA 2.754 ;
 END ZN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.525 2.345 1.665 2.8 ;
 RECT 2.465 2.265 2.605 2.8 ;
 RECT 3.405 2.345 3.545 2.8 ;
 RECT 0.585 2.315 0.725 2.8 ;
 RECT 4.5 1.965 4.64 2.8 ;
 RECT 0 2.8 5.12 2.96 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 3.66 0.275 3.76 1.185 ;
 RECT 3.505 1.185 3.76 1.415 ;
 RECT 3.66 1.415 3.76 2.79 ;
 RECT 3.19 0.275 3.29 1.185 ;
 RECT 3.19 1.415 3.29 2.79 ;
 RECT 3.095 1.185 3.325 1.415 ;
 RECT 2.72 0.275 2.82 1.185 ;
 RECT 2.72 1.415 2.82 2.79 ;
 RECT 2.685 1.185 2.915 1.415 ;
 RECT 2.25 0.275 2.35 1.185 ;
 RECT 2.25 1.185 2.505 1.415 ;
 RECT 2.25 1.415 2.35 2.79 ;
 RECT 0.84 0.275 0.94 1.185 ;
 RECT 0.84 1.415 0.94 2.79 ;
 RECT 0.755 1.185 0.985 1.415 ;
 RECT 1.78 0.275 1.88 1.185 ;
 RECT 1.625 1.185 1.88 1.415 ;
 RECT 1.78 1.415 1.88 2.79 ;
 RECT 1.31 0.275 1.41 1.185 ;
 RECT 1.31 1.415 1.41 2.79 ;
 RECT 1.2 1.185 1.43 1.415 ;
 RECT 0.37 0.275 0.47 1.185 ;
 RECT 0.37 1.415 0.47 2.79 ;
 RECT 0.305 1.185 0.535 1.415 ;
 LAYER CO ;
 RECT 4.505 0.355 4.635 0.485 ;
 RECT 4.505 0.625 4.635 0.755 ;
 RECT 4.505 2.015 4.635 2.145 ;
 RECT 4.505 2.285 4.635 2.415 ;
 RECT 2.94 1.985 3.07 2.115 ;
 RECT 2.47 0.59 2.6 0.72 ;
 RECT 2 2.255 2.13 2.385 ;
 RECT 3.88 0.69 4.01 0.82 ;
 RECT 2.94 0.675 3.07 0.805 ;
 RECT 3.41 2.44 3.54 2.57 ;
 RECT 3.41 0.59 3.54 0.72 ;
 RECT 2.47 2.425 2.6 2.555 ;
 RECT 2 1.985 2.13 2.115 ;
 RECT 2 0.69 2.13 0.82 ;
 RECT 3.88 1.985 4.01 2.115 ;
 RECT 2.94 2.255 3.07 2.385 ;
 RECT 3.555 1.235 3.685 1.365 ;
 RECT 3.145 1.235 3.275 1.365 ;
 RECT 2.735 1.235 2.865 1.365 ;
 RECT 2.325 1.235 2.455 1.365 ;
 RECT 0.59 0.59 0.72 0.72 ;
 RECT 0.59 2.425 0.72 2.555 ;
 RECT 0.355 1.235 0.485 1.365 ;
 RECT 0.805 1.235 0.935 1.365 ;
 RECT 0.12 2.255 0.25 2.385 ;
 RECT 1.53 2.44 1.66 2.57 ;
 RECT 1.675 1.235 1.805 1.365 ;
 RECT 2 1.985 2.13 2.115 ;
 RECT 1.06 1.985 1.19 2.115 ;
 RECT 1.25 1.235 1.38 1.365 ;
 RECT 0.12 1.985 0.25 2.115 ;
 RECT 2 0.69 2.13 0.82 ;
 RECT 0.12 0.69 0.25 0.82 ;
 RECT 1.06 2.255 1.19 2.385 ;
 RECT 1.06 0.675 1.19 0.805 ;
 RECT 1.53 0.59 1.66 0.72 ;
 END
END INVX8

MACRO NAND2X0
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 1.92 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 1.92 2.96 ;
 RECT 0.585 1.575 0.725 2.8 ;
 RECT 1.47 1.735 1.61 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.865 2.075 1.24 2.36 ;
 END
 ANTENNAGATEAREA 0.065 ;
 END IN1

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 1.92 0.08 ;
 RECT 1.495 0.08 1.635 0.855 ;
 RECT 0.115 0.08 0.255 0.69 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 0.835 0.51 1.08 ;
 END
 ANTENNAGATEAREA 0.065 ;
 END IN2

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.115 1.25 1.4 1.4 ;
 RECT 1.055 1.51 1.195 1.76 ;
 RECT 0.115 1.415 0.255 1.76 ;
 RECT 1.05 1.415 1.195 1.51 ;
 RECT 0.115 1.4 1.195 1.415 ;
 RECT 1.045 0.43 1.195 1.15 ;
 RECT 1.045 1.15 1.4 1.25 ;
 END
 ANTENNADIFFAREA 0.315 ;
 END QN

 OBS
 LAYER PO ;
 RECT 0.37 1.08 0.47 2.055 ;
 RECT 0.37 0.26 0.47 0.85 ;
 RECT 0.24 0.85 0.47 1.08 ;
 RECT 0.84 0.26 0.94 2.085 ;
 RECT 0.84 2.085 1.095 2.315 ;
 LAYER CO ;
 RECT 1.475 1.795 1.605 1.925 ;
 RECT 1.5 0.675 1.63 0.805 ;
 RECT 1.06 1.565 1.19 1.695 ;
 RECT 1.5 0.415 1.63 0.545 ;
 RECT 0.29 0.9 0.42 1.03 ;
 RECT 1.475 2.055 1.605 2.185 ;
 RECT 0.12 0.48 0.25 0.61 ;
 RECT 0.915 2.135 1.045 2.265 ;
 RECT 0.59 1.65 0.72 1.78 ;
 RECT 1.06 1.565 1.19 1.695 ;
 RECT 1.06 0.48 1.19 0.61 ;
 RECT 0.12 1.565 0.25 1.695 ;
 END
END NAND2X0

MACRO NAND2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 1.92 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.2 0.81 0.49 1.08 ;
 END
 ANTENNAGATEAREA 0.13 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 1.92 0.08 ;
 RECT 0.135 0.08 0.275 0.58 ;
 RECT 1.515 0.08 1.655 0.855 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 1.92 2.96 ;
 RECT 0.605 1.93 0.745 2.8 ;
 RECT 1.49 1.485 1.63 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.635 0.765 0.92 1.085 ;
 END
 ANTENNAGATEAREA 0.13 ;
 END IN1

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.07 1.06 1.36 1.34 ;
 RECT 1.07 1.34 1.215 1.35 ;
 RECT 1.07 0.27 1.215 1.06 ;
 RECT 0.135 1.68 0.275 2.265 ;
 RECT 0.135 1.415 0.275 1.515 ;
 RECT 1.075 1.68 1.215 2.265 ;
 RECT 0.135 1.515 1.215 1.68 ;
 RECT 1.075 1.35 1.215 1.515 ;
 END
 ANTENNADIFFAREA 0.63 ;
 END QN

 OBS
 LAYER PO ;
 RECT 0.39 1.08 0.49 2.455 ;
 RECT 0.39 0.1 0.49 0.85 ;
 RECT 0.26 0.85 0.49 1.08 ;
 RECT 0.86 0.1 0.96 0.855 ;
 RECT 0.68 0.855 0.96 1.085 ;
 RECT 0.86 1.085 0.96 2.455 ;
 LAYER CO ;
 RECT 0.14 2.035 0.27 2.165 ;
 RECT 1.08 2.05 1.21 2.18 ;
 RECT 1.08 1.78 1.21 1.91 ;
 RECT 0.14 1.775 0.27 1.905 ;
 RECT 1.52 0.415 1.65 0.545 ;
 RECT 1.495 2.055 1.625 2.185 ;
 RECT 1.495 1.795 1.625 1.925 ;
 RECT 1.495 1.535 1.625 1.665 ;
 RECT 1.52 0.675 1.65 0.805 ;
 RECT 0.14 0.32 0.27 0.45 ;
 RECT 0.14 1.505 0.27 1.635 ;
 RECT 1.08 0.32 1.21 0.45 ;
 RECT 0.61 2.03 0.74 2.16 ;
 RECT 0.31 0.9 0.44 1.03 ;
 RECT 0.73 0.905 0.86 1.035 ;
 RECT 1.08 1.51 1.21 1.64 ;
 END
END NAND2X1

MACRO NAND2X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.11 1.56 1.405 ;
 END
 ANTENNAGATEAREA 0.26 ;
 END IN1

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.725 1.76 2.035 2.075 ;
 RECT 1.725 0.71 1.87 1.26 ;
 RECT 0.79 1.76 0.93 2.3 ;
 RECT 0.79 1.54 0.93 1.595 ;
 RECT 0.79 1.595 1.87 1.76 ;
 RECT 1.73 1.26 1.87 1.595 ;
 END
 ANTENNADIFFAREA 0.778 ;
 END QN

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.84 1.11 1.145 1.4 ;
 END
 ANTENNAGATEAREA 0.26 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 2.66 0.08 2.8 0.855 ;
 RECT 0.79 0.08 0.93 0.655 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 2.635 1.485 2.775 2.8 ;
 RECT 1.26 1.96 1.4 2.8 ;
 RECT 2.205 1.55 2.345 2.8 ;
 RECT 0.315 1.55 0.455 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 1.045 0.255 1.145 1.12 ;
 RECT 0.575 0.255 0.675 1.19 ;
 RECT 0.575 1.29 0.675 2.495 ;
 RECT 1.045 1.35 1.145 2.485 ;
 RECT 0.915 1.12 1.145 1.19 ;
 RECT 0.915 1.29 1.145 1.35 ;
 RECT 0.575 1.19 1.145 1.29 ;
 RECT 1.34 1.17 1.615 1.4 ;
 RECT 1.515 1.4 1.615 2.5 ;
 RECT 1.985 0.255 2.085 1.07 ;
 RECT 1.985 1.17 2.085 2.505 ;
 RECT 1.515 0.255 1.615 1.07 ;
 RECT 1.515 1.07 2.085 1.17 ;
 LAYER CO ;
 RECT 0.795 1.59 0.925 1.72 ;
 RECT 2.21 0.745 2.34 0.875 ;
 RECT 1.265 0.735 1.395 0.865 ;
 RECT 0.325 0.745 0.455 0.875 ;
 RECT 0.32 2.12 0.45 2.25 ;
 RECT 0.32 1.86 0.45 1.99 ;
 RECT 2.21 2.125 2.34 2.255 ;
 RECT 2.21 1.865 2.34 1.995 ;
 RECT 0.795 2.12 0.925 2.25 ;
 RECT 0.795 1.86 0.925 1.99 ;
 RECT 0.325 0.475 0.455 0.605 ;
 RECT 2.21 0.475 2.34 0.605 ;
 RECT 1.265 0.475 1.395 0.605 ;
 RECT 0.32 1.6 0.45 1.73 ;
 RECT 0.32 1.6 0.45 1.73 ;
 RECT 2.21 1.6 2.34 1.73 ;
 RECT 2.21 1.6 2.34 1.73 ;
 RECT 0.965 1.17 1.095 1.3 ;
 RECT 1.265 2.06 1.395 2.19 ;
 RECT 1.735 1.815 1.865 1.945 ;
 RECT 2.64 1.535 2.77 1.665 ;
 RECT 2.64 1.795 2.77 1.925 ;
 RECT 2.64 2.055 2.77 2.185 ;
 RECT 2.665 0.415 2.795 0.545 ;
 RECT 1.735 0.765 1.865 0.895 ;
 RECT 2.665 0.675 2.795 0.805 ;
 RECT 1.735 1.545 1.865 1.675 ;
 RECT 1.39 1.22 1.52 1.35 ;
 RECT 0.795 0.475 0.925 0.605 ;
 LAYER M1 ;
 RECT 0.32 0.405 0.46 0.83 ;
 RECT 1.26 0.515 1.4 0.83 ;
 RECT 0.32 0.83 1.4 0.97 ;
 RECT 2.205 0.515 2.345 0.945 ;
 RECT 1.26 0.375 2.345 0.515 ;
 END
END NAND2X2

MACRO NAND2X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.73 0.64 3.875 1.35 ;
 RECT 2.775 0.64 2.92 1.35 ;
 RECT 3.735 1.71 3.875 2.32 ;
 RECT 3.735 1.63 3.98 1.71 ;
 RECT 3.735 1.47 3.98 1.49 ;
 RECT 3.735 1.35 3.875 1.47 ;
 RECT 0.88 1.81 1.02 2.26 ;
 RECT 0.88 1.495 1.02 1.645 ;
 RECT 1.84 1.81 1.98 2.26 ;
 RECT 2.78 1.81 2.92 2.31 ;
 RECT 0.875 1.645 2.92 1.81 ;
 RECT 2.78 1.63 2.92 1.645 ;
 RECT 2.78 1.49 3.98 1.63 ;
 RECT 2.78 1.35 2.92 1.49 ;
 END
 ANTENNADIFFAREA 1.57 ;
 END QN

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.605 1.125 2.06 1.435 ;
 END
 ANTENNAGATEAREA 0.52 ;
 END IN2

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 1.365 2.025 1.505 2.8 ;
 RECT 2.31 1.96 2.45 2.8 ;
 RECT 4.215 1.55 4.355 2.8 ;
 RECT 0.405 1.505 0.545 2.8 ;
 RECT 3.255 1.78 3.395 2.8 ;
 RECT 4.645 1.485 4.785 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 1.775 0.445 2.045 0.585 ;
 RECT 0.815 0.445 1.085 0.585 ;
 RECT 4.67 0.08 4.81 0.855 ;
 RECT 1.84 0.08 1.98 0.445 ;
 RECT 0.88 0.08 1.02 0.445 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.035 0.84 4.375 1.245 ;
 END
 ANTENNAGATEAREA 0.52 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 1.625 1.195 1.915 1.24 ;
 RECT 1.625 0.23 1.725 1.195 ;
 RECT 1.625 1.34 1.915 1.425 ;
 RECT 1.625 1.425 1.725 2.495 ;
 RECT 0.66 0.23 0.76 1.24 ;
 RECT 1.14 0.23 1.24 1.24 ;
 RECT 2.095 0.23 2.195 1.24 ;
 RECT 0.66 1.34 0.76 2.495 ;
 RECT 1.14 1.34 1.24 2.495 ;
 RECT 2.095 1.34 2.195 2.485 ;
 RECT 0.66 1.24 2.195 1.34 ;
 RECT 3.995 1.005 4.375 1.045 ;
 RECT 3.52 0.23 3.62 1.045 ;
 RECT 3.52 1.145 3.62 2.505 ;
 RECT 2.565 0.23 2.665 1.045 ;
 RECT 2.565 1.145 2.665 2.5 ;
 RECT 3.995 1.145 4.375 1.235 ;
 RECT 3.995 1.235 4.095 2.505 ;
 RECT 3.995 0.23 4.095 1.005 ;
 RECT 2.565 1.045 4.375 1.145 ;
 RECT 3.035 0.23 3.135 1.045 ;
 RECT 3.035 1.145 3.135 2.505 ;
 LAYER CO ;
 RECT 4.65 1.795 4.78 1.925 ;
 RECT 1.72 1.245 1.85 1.375 ;
 RECT 2.785 1.815 2.915 1.945 ;
 RECT 4.675 0.675 4.805 0.805 ;
 RECT 1.845 2.07 1.975 2.2 ;
 RECT 4.65 2.055 4.78 2.185 ;
 RECT 2.315 0.45 2.445 0.58 ;
 RECT 1.845 0.45 1.975 0.58 ;
 RECT 4.675 0.415 4.805 0.545 ;
 RECT 2.785 0.74 2.915 0.87 ;
 RECT 4.65 1.535 4.78 1.665 ;
 RECT 1.375 0.45 1.505 0.58 ;
 RECT 4.195 1.055 4.325 1.185 ;
 RECT 2.785 1.545 2.915 1.675 ;
 RECT 0.41 1.58 0.54 1.71 ;
 RECT 0.41 1.86 0.54 1.99 ;
 RECT 2.785 2.08 2.915 2.21 ;
 RECT 3.26 2.12 3.39 2.25 ;
 RECT 3.26 1.86 3.39 1.99 ;
 RECT 3.74 2.075 3.87 2.205 ;
 RECT 4.22 2.125 4.35 2.255 ;
 RECT 4.22 1.86 4.35 1.99 ;
 RECT 0.41 0.45 0.54 0.58 ;
 RECT 0.41 2.12 0.54 2.25 ;
 RECT 0.885 0.45 1.015 0.58 ;
 RECT 0.885 1.545 1.015 1.675 ;
 RECT 0.885 2.07 1.015 2.2 ;
 RECT 0.885 1.805 1.015 1.935 ;
 RECT 0.885 1.545 1.015 1.675 ;
 RECT 4.215 0.45 4.345 0.58 ;
 RECT 4.22 1.6 4.35 1.73 ;
 RECT 4.22 1.6 4.35 1.73 ;
 RECT 3.74 1.545 3.87 1.675 ;
 RECT 3.74 0.74 3.87 0.87 ;
 RECT 3.74 1.815 3.87 1.945 ;
 RECT 2.315 2.06 2.445 2.19 ;
 RECT 1.845 1.805 1.975 1.935 ;
 RECT 3.26 0.45 3.39 0.58 ;
 RECT 1.37 2.12 1.5 2.25 ;
 LAYER M1 ;
 RECT 3.255 0.49 3.395 0.67 ;
 RECT 2.31 0.35 3.395 0.49 ;
 RECT 0.405 0.725 1.535 0.865 ;
 RECT 1.37 0.38 1.51 0.73 ;
 RECT 0.405 0.35 0.545 0.865 ;
 RECT 2.31 0.49 2.45 0.73 ;
 RECT 1.37 0.73 2.45 0.87 ;
 RECT 4.21 0.49 4.35 0.69 ;
 RECT 3.275 0.35 4.35 0.49 ;
 END
END NAND2X4

MACRO NAND3X0
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 RECT 1.585 1.805 1.725 2.8 ;
 RECT 0.645 1.45 0.785 2.8 ;
 RECT 0.23 1.51 0.37 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 RECT 0.645 0.08 0.785 0.805 ;
 RECT 0.23 0.08 0.37 0.845 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.745 1 2.04 1.24 ;
 RECT 1.115 1.525 2.2 1.665 ;
 RECT 1.695 0.31 2.245 0.455 ;
 RECT 2.06 1.665 2.2 1.915 ;
 RECT 1.115 1.665 1.255 1.89 ;
 RECT 1.745 1.24 1.885 1.525 ;
 RECT 2.06 0.455 2.2 0.8 ;
 RECT 2.06 0.245 2.2 0.31 ;
 RECT 1.745 0.455 1.885 1 ;
 END
 ANTENNADIFFAREA 0.55 ;
 END QN

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.925 2.1 1.24 2.36 ;
 END
 ANTENNAGATEAREA 0.11 ;
 END IN3

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 0.84 1.56 1.105 ;
 END
 ANTENNAGATEAREA 0.11 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.87 2.38 2.2 2.655 ;
 END
 ANTENNAGATEAREA 0.11 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 1.84 0.1 1.94 2.41 ;
 RECT 1.84 2.64 1.94 2.655 ;
 RECT 1.84 2.41 2.07 2.64 ;
 RECT 0.9 0.1 1 2.125 ;
 RECT 0.9 2.125 1.13 2.355 ;
 RECT 1.37 1.105 1.47 2.23 ;
 RECT 1.37 0.1 1.47 0.875 ;
 RECT 1.315 0.875 1.545 1.105 ;
 LAYER CO ;
 RECT 2.065 0.585 2.195 0.715 ;
 RECT 0.65 0.585 0.78 0.715 ;
 RECT 0.65 1.855 0.78 1.985 ;
 RECT 1.59 1.855 1.72 1.985 ;
 RECT 2.065 1.69 2.195 1.82 ;
 RECT 1.89 2.46 2.02 2.59 ;
 RECT 0.235 0.405 0.365 0.535 ;
 RECT 0.235 2.08 0.365 2.21 ;
 RECT 0.65 1.595 0.78 1.725 ;
 RECT 0.235 0.665 0.365 0.795 ;
 RECT 1.12 1.675 1.25 1.805 ;
 RECT 0.95 2.175 1.08 2.305 ;
 RECT 0.235 1.56 0.365 1.69 ;
 RECT 0.235 1.82 0.365 1.95 ;
 RECT 1.365 0.925 1.495 1.055 ;
 RECT 0.65 0.32 0.78 0.45 ;
 RECT 2.065 0.32 2.195 0.45 ;
 END
END NAND3X0

MACRO NAND3X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 3.17 1.395 3.31 2.8 ;
 RECT 0.23 1.51 0.37 2.8 ;
 RECT 0.645 1.55 0.785 2.8 ;
 RECT 1.585 1.545 1.725 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.12 1.95 1.435 2.295 ;
 END
 ANTENNAGATEAREA 0.058 ;
 END IN2

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.575 1.15 0.92 1.405 ;
 END
 ANTENNAGATEAREA 0.058 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 0.645 0.08 0.785 0.55 ;
 RECT 0.23 0.08 0.37 0.75 ;
 RECT 3.02 0.08 3.16 0.875 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.93 0.84 2.28 1.08 ;
 END
 ANTENNAGATEAREA 0.058 ;
 END IN1

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.56 1.16 3.8 1.465 ;
 RECT 3.66 1.465 3.8 2.595 ;
 RECT 3.66 0.29 3.8 1.16 ;
 END
 ANTENNADIFFAREA 0.502 ;
 END QN

 OBS
 LAYER PO ;
 RECT 0.9 1.395 1 2.01 ;
 RECT 0.9 0.1 1 1.165 ;
 RECT 0.705 1.165 1 1.395 ;
 RECT 1.84 0.1 1.94 0.865 ;
 RECT 1.84 0.865 2.16 1.095 ;
 RECT 1.84 1.095 1.94 2.005 ;
 RECT 2.795 0.395 2.895 1.95 ;
 RECT 2.735 1.95 2.965 2.18 ;
 RECT 1.37 0.1 1.47 1.95 ;
 RECT 1.24 1.95 1.47 2.18 ;
 RECT 3.435 0.11 3.535 1 ;
 RECT 3.435 1.23 3.535 2.765 ;
 RECT 3.185 1 3.535 1.23 ;
 LAYER CO ;
 RECT 3.175 1.59 3.305 1.72 ;
 RECT 3.665 1.59 3.795 1.72 ;
 RECT 1.59 1.645 1.72 1.775 ;
 RECT 0.65 1.645 0.78 1.775 ;
 RECT 2.065 1.645 2.195 1.775 ;
 RECT 1.12 1.57 1.25 1.7 ;
 RECT 0.235 2.08 0.365 2.21 ;
 RECT 0.235 1.56 0.365 1.69 ;
 RECT 0.235 1.82 0.365 1.95 ;
 RECT 0.65 0.32 0.78 0.45 ;
 RECT 0.755 1.215 0.885 1.345 ;
 RECT 1.98 0.915 2.11 1.045 ;
 RECT 2.065 0.32 2.195 0.45 ;
 RECT 1.29 2 1.42 2.13 ;
 RECT 0.235 0.31 0.365 0.44 ;
 RECT 0.235 0.57 0.365 0.7 ;
 RECT 3.665 2.11 3.795 2.24 ;
 RECT 2.505 0.63 2.635 0.76 ;
 RECT 2.785 2 2.915 2.13 ;
 RECT 3.175 1.85 3.305 1.98 ;
 RECT 3.235 1.05 3.365 1.18 ;
 RECT 3.665 0.36 3.795 0.49 ;
 RECT 3.665 0.62 3.795 0.75 ;
 RECT 3.025 0.63 3.155 0.76 ;
 RECT 3.665 1.85 3.795 1.98 ;
 RECT 3.665 2.375 3.795 2.505 ;
 RECT 2.505 1.59 2.635 1.72 ;
 RECT 3.175 2.11 3.305 2.24 ;
 LAYER M1 ;
 RECT 2.5 0.58 2.64 1.04 ;
 RECT 2.5 1.19 2.64 1.82 ;
 RECT 2.5 1.04 3.415 1.19 ;
 RECT 1.115 1.39 1.255 1.79 ;
 RECT 1.65 0.455 1.79 1.25 ;
 RECT 2.06 1.39 2.2 2.025 ;
 RECT 1.115 1.25 2.2 1.39 ;
 RECT 2.735 1.95 2.965 2.025 ;
 RECT 2.735 2.165 2.965 2.18 ;
 RECT 2.06 2.025 2.965 2.165 ;
 RECT 1.63 0.31 2.245 0.455 ;
 END
END NAND3X1

MACRO NAND3X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.59 1.16 0.92 1.4 ;
 END
 ANTENNAGATEAREA 0.058 ;
 END IN3

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 1.91 1.445 2.36 ;
 END
 ANTENNAGATEAREA 0.058 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 0.23 0.08 0.37 0.77 ;
 RECT 0.645 0.08 0.785 0.55 ;
 RECT 3.02 0.08 3.16 0.865 ;
 RECT 4.145 0.08 4.285 0.865 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.93 0.84 2.215 1.105 ;
 END
 ANTENNAGATEAREA 0.058 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 0.23 1.51 0.37 2.8 ;
 RECT 3.17 1.415 3.31 2.8 ;
 RECT 4.145 1.37 4.285 2.8 ;
 RECT 0.645 1.55 0.785 2.8 ;
 RECT 1.585 1.56 1.725 2.8 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.56 1.15 3.8 1.405 ;
 RECT 3.66 1.405 3.8 2.63 ;
 RECT 3.66 0.32 3.8 1.15 ;
 END
 ANTENNADIFFAREA 0.616 ;
 END QN

 OBS
 LAYER PO ;
 RECT 2.795 0.43 2.895 1.945 ;
 RECT 2.795 2.175 2.895 2.22 ;
 RECT 2.735 1.945 2.965 2.175 ;
 RECT 3.435 1.25 3.535 2.77 ;
 RECT 3.915 0.145 4.015 1.115 ;
 RECT 3.915 1.215 4.015 2.77 ;
 RECT 3.195 1.02 3.535 1.115 ;
 RECT 3.195 1.215 3.535 1.25 ;
 RECT 3.195 1.115 4.015 1.215 ;
 RECT 3.435 0.145 3.535 1.02 ;
 RECT 1.37 0.1 1.47 1.91 ;
 RECT 1.24 1.91 1.47 2.14 ;
 RECT 0.9 0.1 1 1.165 ;
 RECT 0.9 1.395 1 2.01 ;
 RECT 0.705 1.165 1 1.395 ;
 RECT 1.84 0.1 1.94 0.865 ;
 RECT 1.84 1.095 1.94 2.005 ;
 RECT 1.84 0.865 2.16 1.095 ;
 LAYER CO ;
 RECT 1.12 1.575 1.25 1.705 ;
 RECT 0.755 1.215 0.885 1.345 ;
 RECT 3.665 1.845 3.795 1.975 ;
 RECT 3.235 1.07 3.365 1.2 ;
 RECT 3.025 0.66 3.155 0.79 ;
 RECT 2.505 1.585 2.635 1.715 ;
 RECT 0.235 2.08 0.365 2.21 ;
 RECT 0.235 1.56 0.365 1.69 ;
 RECT 3.175 1.585 3.305 1.715 ;
 RECT 0.235 1.82 0.365 1.95 ;
 RECT 1.29 1.96 1.42 2.09 ;
 RECT 3.665 0.65 3.795 0.78 ;
 RECT 4.15 0.66 4.28 0.79 ;
 RECT 4.15 2.105 4.28 2.235 ;
 RECT 4.15 1.585 4.28 1.715 ;
 RECT 4.15 1.845 4.28 1.975 ;
 RECT 3.175 2.105 3.305 2.235 ;
 RECT 3.665 1.585 3.795 1.715 ;
 RECT 1.59 1.645 1.72 1.775 ;
 RECT 2.785 1.995 2.915 2.125 ;
 RECT 2.065 1.645 2.195 1.775 ;
 RECT 0.65 0.32 0.78 0.45 ;
 RECT 3.665 2.105 3.795 2.235 ;
 RECT 3.175 1.845 3.305 1.975 ;
 RECT 1.98 0.915 2.11 1.045 ;
 RECT 3.665 0.39 3.795 0.52 ;
 RECT 2.065 0.32 2.195 0.45 ;
 RECT 0.235 0.33 0.365 0.46 ;
 RECT 3.665 2.37 3.795 2.5 ;
 RECT 2.505 0.66 2.635 0.79 ;
 RECT 0.65 1.645 0.78 1.775 ;
 RECT 0.235 0.59 0.365 0.72 ;
 LAYER M1 ;
 RECT 2.5 0.61 2.64 1.08 ;
 RECT 2.5 1.23 2.64 1.875 ;
 RECT 3.23 1.015 3.37 1.08 ;
 RECT 3.23 1.23 3.37 1.25 ;
 RECT 2.5 1.08 3.42 1.23 ;
 RECT 1.115 1.41 1.255 1.765 ;
 RECT 1.65 0.455 1.79 1.27 ;
 RECT 2.06 1.41 2.2 2.105 ;
 RECT 2.06 1.25 2.2 1.27 ;
 RECT 1.115 1.275 2.2 1.41 ;
 RECT 1.165 1.27 2.2 1.275 ;
 RECT 2.78 1.945 2.92 2.105 ;
 RECT 2.06 2.105 2.92 2.245 ;
 RECT 1.63 0.31 2.245 0.455 ;
 END
END NAND3X2

MACRO NAND3X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 4.145 1.37 4.285 2.8 ;
 RECT 3.17 1.425 3.31 2.8 ;
 RECT 5.13 1.37 5.27 2.8 ;
 RECT 0.23 1.51 0.37 2.8 ;
 RECT 1.585 1.56 1.725 2.8 ;
 RECT 0.645 1.55 0.785 2.8 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.56 1.16 3.885 1.415 ;
 RECT 3.66 1.415 3.8 2.64 ;
 RECT 3.66 0.87 4.76 1.01 ;
 RECT 4.62 1.01 4.76 2.645 ;
 RECT 4.62 0.32 4.76 0.87 ;
 RECT 3.66 1.01 3.8 1.16 ;
 RECT 3.66 0.32 3.8 0.87 ;
 END
 ANTENNADIFFAREA 1.264 ;
 END QN

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.515 1.16 0.925 1.4 ;
 END
 ANTENNAGATEAREA 0.058 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 0.23 0.08 0.37 0.77 ;
 RECT 0.645 0.08 0.785 0.55 ;
 RECT 4.145 0.08 4.285 0.63 ;
 RECT 3.02 0.08 3.16 0.865 ;
 RECT 5.125 0.08 5.265 0.79 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.11 1.94 1.445 2.285 ;
 END
 ANTENNAGATEAREA 0.058 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.93 0.84 2.225 1.125 ;
 END
 ANTENNAGATEAREA 0.058 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 0.9 0.1 1 1.165 ;
 RECT 0.705 1.165 1 1.395 ;
 RECT 0.9 1.395 1 2.01 ;
 RECT 3.14 1.02 3.535 1.115 ;
 RECT 3.435 0.145 3.535 1.02 ;
 RECT 3.14 1.215 3.535 1.25 ;
 RECT 3.435 1.25 3.535 2.765 ;
 RECT 3.915 0.145 4.015 1.115 ;
 RECT 3.915 1.215 4.015 2.765 ;
 RECT 4.4 0.145 4.5 1.115 ;
 RECT 4.4 1.215 4.5 2.765 ;
 RECT 4.9 0.145 5 1.115 ;
 RECT 4.9 1.215 5 2.765 ;
 RECT 3.14 1.115 5 1.215 ;
 RECT 1.84 0.1 1.94 0.865 ;
 RECT 1.84 0.865 2.16 1.095 ;
 RECT 1.84 1.095 1.94 2.005 ;
 RECT 2.795 0.43 2.895 1.94 ;
 RECT 2.735 1.94 2.965 2.17 ;
 RECT 1.37 0.1 1.47 1.96 ;
 RECT 1.24 1.96 1.47 2.19 ;
 LAYER CO ;
 RECT 5.13 0.44 5.26 0.57 ;
 RECT 5.135 1.58 5.265 1.71 ;
 RECT 5.135 2.1 5.265 2.23 ;
 RECT 5.135 1.84 5.265 1.97 ;
 RECT 4.625 1.84 4.755 1.97 ;
 RECT 4.625 2.1 4.755 2.23 ;
 RECT 4.625 2.365 4.755 2.495 ;
 RECT 4.625 0.65 4.755 0.78 ;
 RECT 4.625 0.39 4.755 0.52 ;
 RECT 4.625 1.58 4.755 1.71 ;
 RECT 3.665 0.39 3.795 0.52 ;
 RECT 3.025 0.66 3.155 0.79 ;
 RECT 3.665 1.58 3.795 1.71 ;
 RECT 2.065 1.645 2.195 1.775 ;
 RECT 3.665 2.1 3.795 2.23 ;
 RECT 3.665 1.84 3.795 1.97 ;
 RECT 0.235 1.56 0.365 1.69 ;
 RECT 3.665 2.365 3.795 2.495 ;
 RECT 2.505 1.58 2.635 1.71 ;
 RECT 0.755 1.215 0.885 1.345 ;
 RECT 3.175 2.1 3.305 2.23 ;
 RECT 0.65 0.32 0.78 0.45 ;
 RECT 0.235 1.82 0.365 1.95 ;
 RECT 0.235 0.59 0.365 0.72 ;
 RECT 3.175 1.58 3.305 1.71 ;
 RECT 2.065 0.32 2.195 0.45 ;
 RECT 3.18 1.07 3.31 1.2 ;
 RECT 0.235 2.08 0.365 2.21 ;
 RECT 2.785 1.99 2.915 2.12 ;
 RECT 0.65 1.645 0.78 1.775 ;
 RECT 1.29 2.01 1.42 2.14 ;
 RECT 1.12 1.585 1.25 1.715 ;
 RECT 1.59 1.645 1.72 1.775 ;
 RECT 0.235 0.33 0.365 0.46 ;
 RECT 1.98 0.915 2.11 1.045 ;
 RECT 4.15 1.58 4.28 1.71 ;
 RECT 3.175 1.84 3.305 1.97 ;
 RECT 4.15 1.84 4.28 1.97 ;
 RECT 4.15 0.44 4.28 0.57 ;
 RECT 4.15 2.1 4.28 2.23 ;
 RECT 3.665 0.65 3.795 0.78 ;
 RECT 2.505 0.66 2.635 0.79 ;
 LAYER M1 ;
 RECT 2.5 0.61 2.64 1.135 ;
 RECT 2.5 1.285 2.64 1.89 ;
 RECT 3.175 1.015 3.315 1.135 ;
 RECT 2.5 1.135 3.42 1.285 ;
 RECT 1.115 1.41 1.255 1.8 ;
 RECT 1.65 0.455 1.79 1.27 ;
 RECT 2.06 1.41 2.2 2.1 ;
 RECT 1.115 1.275 2.2 1.41 ;
 RECT 1.165 1.27 2.2 1.275 ;
 RECT 2.78 1.94 2.92 2.1 ;
 RECT 2.06 2.1 2.92 2.24 ;
 RECT 1.63 0.31 2.245 0.455 ;
 END
END NAND3X4

MACRO NAND4X0
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.88 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.655 1.155 1.005 1.395 ;
 END
 ANTENNAGATEAREA 0.101 ;
 END IN1

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.2 1.28 2.28 1.42 ;
 RECT 1.62 1.16 1.86 1.28 ;
 RECT 1.2 1.42 1.34 1.79 ;
 RECT 2.14 1.42 2.28 1.79 ;
 RECT 0.73 0.475 1.805 0.615 ;
 RECT 0.73 0.275 0.87 0.475 ;
 RECT 1.665 0.615 1.805 1.16 ;
 END
 ANTENNADIFFAREA 0.517 ;
 END QN

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.27 2.055 1.53 2.365 ;
 END
 ANTENNAGATEAREA 0.101 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.88 0.08 ;
 RECT 0.315 0.08 0.455 0.91 ;
 RECT 2.615 0.08 2.755 0.505 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.88 2.96 ;
 RECT 1.67 1.64 1.81 2.8 ;
 RECT 0.73 1.555 0.87 2.8 ;
 RECT 2.62 1.54 2.76 2.8 ;
 RECT 0.32 1.495 0.46 2.8 ;
 END
 END VDD

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.96 2.065 2.255 2.365 ;
 END
 ANTENNAGATEAREA 0.101 ;
 END IN3

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.42 1.155 2.795 1.4 ;
 END
 ANTENNAGATEAREA 0.101 ;
 END IN4

 OBS
 LAYER PO ;
 RECT 1.925 0.105 2.025 2.065 ;
 RECT 1.915 2.065 2.145 2.295 ;
 RECT 2.4 0.1 2.5 1.165 ;
 RECT 2.4 1.165 2.655 1.395 ;
 RECT 2.4 1.395 2.5 2.425 ;
 RECT 0.985 0.105 1.085 1.165 ;
 RECT 0.775 1.165 1.085 1.395 ;
 RECT 0.985 1.395 1.085 2.18 ;
 RECT 1.455 0.105 1.555 2.055 ;
 RECT 1.3 2.055 1.555 2.175 ;
 RECT 1.3 2.175 1.53 2.285 ;
 LAYER CO ;
 RECT 1.965 2.115 2.095 2.245 ;
 RECT 1.675 1.74 1.805 1.87 ;
 RECT 1.205 1.61 1.335 1.74 ;
 RECT 2.475 1.215 2.605 1.345 ;
 RECT 0.325 1.805 0.455 1.935 ;
 RECT 2.62 0.325 2.75 0.455 ;
 RECT 0.32 0.73 0.45 0.86 ;
 RECT 0.735 0.325 0.865 0.455 ;
 RECT 1.35 2.105 1.48 2.235 ;
 RECT 2.145 1.61 2.275 1.74 ;
 RECT 2.625 1.72 2.755 1.85 ;
 RECT 0.825 1.215 0.955 1.345 ;
 RECT 0.325 2.065 0.455 2.195 ;
 RECT 0.325 1.545 0.455 1.675 ;
 RECT 2.145 1.61 2.275 1.74 ;
 RECT 0.735 1.61 0.865 1.74 ;
 RECT 0.32 0.47 0.45 0.6 ;
 END
END NAND4X0

MACRO NAND4X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.48 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.48 2.96 ;
 RECT 0.78 1.695 0.92 2.8 ;
 RECT 2.67 1.855 2.81 2.8 ;
 RECT 1.72 1.89 1.86 2.8 ;
 RECT 0.37 1.495 0.51 2.8 ;
 RECT 3.6 1.515 3.74 2.8 ;
 END
 END VDD

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.425 1 2.68 1.4 ;
 END
 ANTENNAGATEAREA 0.1 ;
 END IN4

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.77 1.16 1.08 1.4 ;
 END
 ANTENNAGATEAREA 0.1 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.22 0.84 1.56 1.11 ;
 END
 ANTENNAGATEAREA 0.1 ;
 END IN2

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2 2.18 2.36 2.555 ;
 END
 ANTENNAGATEAREA 0.1 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.48 0.08 ;
 RECT 3.595 0.08 3.735 0.655 ;
 RECT 2.67 0.08 2.81 0.505 ;
 RECT 0.365 0.08 0.505 0.91 ;
 END
 END VSS

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.04 0.825 4.28 1.085 ;
 RECT 4.085 1.085 4.225 2.555 ;
 RECT 4.085 0.375 4.225 0.825 ;
 END
 ANTENNADIFFAREA 0.52 ;
 END QN

 OBS
 LAYER PO ;
 RECT 3.855 0.175 3.955 1.135 ;
 RECT 3.67 1.135 3.955 1.365 ;
 RECT 3.855 1.365 3.955 2.76 ;
 RECT 1.505 0.105 1.605 0.87 ;
 RECT 1.505 1.1 1.605 2.455 ;
 RECT 1.315 0.87 1.605 1.1 ;
 RECT 2.45 0.1 2.55 1.165 ;
 RECT 2.45 1.395 2.55 2.455 ;
 RECT 2.425 1.165 2.655 1.395 ;
 RECT 1.975 0.105 2.075 2.325 ;
 RECT 1.975 2.325 2.195 2.555 ;
 RECT 3 0.395 3.1 1.45 ;
 RECT 3 1.68 3.1 2.585 ;
 RECT 2.845 1.45 3.1 1.68 ;
 RECT 1.035 1.395 1.135 2.445 ;
 RECT 1.035 0.105 1.135 1.165 ;
 RECT 0.825 1.165 1.135 1.395 ;
 LAYER CO ;
 RECT 3.225 0.615 3.355 0.745 ;
 RECT 0.37 0.47 0.5 0.6 ;
 RECT 1.365 0.92 1.495 1.05 ;
 RECT 2.895 1.5 3.025 1.63 ;
 RECT 2.195 1.8 2.325 1.93 ;
 RECT 0.375 2.065 0.505 2.195 ;
 RECT 0.875 1.215 1.005 1.345 ;
 RECT 2.015 2.375 2.145 2.505 ;
 RECT 1.725 1.99 1.855 2.12 ;
 RECT 3.225 2.135 3.355 2.265 ;
 RECT 1.255 2.07 1.385 2.2 ;
 RECT 0.785 2.06 0.915 2.19 ;
 RECT 4.09 2.345 4.22 2.475 ;
 RECT 4.09 2.08 4.22 2.21 ;
 RECT 4.09 1.82 4.22 1.95 ;
 RECT 3.605 2.36 3.735 2.49 ;
 RECT 3.605 2.095 3.735 2.225 ;
 RECT 3.605 1.835 3.735 1.965 ;
 RECT 0.785 0.59 0.915 0.72 ;
 RECT 3.6 0.45 3.73 0.58 ;
 RECT 3.605 1.565 3.735 1.695 ;
 RECT 4.09 1.56 4.22 1.69 ;
 RECT 4.09 0.475 4.22 0.605 ;
 RECT 2.675 1.97 2.805 2.1 ;
 RECT 3.72 1.185 3.85 1.315 ;
 RECT 0.785 1.8 0.915 1.93 ;
 RECT 2.475 1.215 2.605 1.345 ;
 RECT 0.375 1.545 0.505 1.675 ;
 RECT 3.225 1.86 3.355 1.99 ;
 RECT 0.785 0.325 0.915 0.455 ;
 RECT 0.37 0.73 0.5 0.86 ;
 RECT 2.675 0.325 2.805 0.455 ;
 RECT 1.255 1.795 1.385 1.925 ;
 RECT 0.375 1.805 0.505 1.935 ;
 LAYER M1 ;
 RECT 3.22 0.27 3.36 0.965 ;
 RECT 3.22 1.105 3.36 2.385 ;
 RECT 3.22 0.965 3.9 1.105 ;
 RECT 3.675 1.105 3.9 1.375 ;
 RECT 0.78 0.275 0.92 0.475 ;
 RECT 0.78 0.615 0.92 0.795 ;
 RECT 1.7 0.615 1.84 1.57 ;
 RECT 0.78 0.475 1.84 0.615 ;
 RECT 1.25 1.71 1.39 2.255 ;
 RECT 2.19 1.715 2.33 2.04 ;
 RECT 1.25 1.57 2.33 1.575 ;
 RECT 2.845 1.49 3.075 1.575 ;
 RECT 2.19 1.71 3.075 1.715 ;
 RECT 1.25 1.575 3.075 1.71 ;
 END
END NAND4X1

MACRO NBUFFX16
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.28 BY 2.88 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.36 1.35 0.89 1.395 ;
 RECT 0.35 1.21 0.89 1.35 ;
 RECT 0.36 1.165 0.89 1.21 ;
 RECT 0.36 1.395 0.84 1.4 ;
 RECT 0.36 1.16 0.84 1.165 ;
 END
 ANTENNAGATEAREA 0.298 ;
 END INP

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.28 0.08 ;
 RECT 8.475 0.755 8.845 0.895 ;
 RECT 8.475 0.08 8.615 0.755 ;
 RECT 8.93 0.08 9.07 0.4 ;
 RECT 4.9 0.08 5.04 0.755 ;
 RECT 6.78 0.08 6.92 0.77 ;
 RECT 2.08 0.08 2.22 0.77 ;
 RECT 3.02 0.08 3.16 0.77 ;
 RECT 3.96 0.08 4.1 0.77 ;
 RECT 1.14 0.08 1.28 0.735 ;
 RECT 5.84 0.08 5.98 0.77 ;
 RECT 7.72 0.08 7.86 0.77 ;
 RECT 0.2 0.08 0.34 0.81 ;
 END
 END VSS

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.61 1.645 8.33 1.78 ;
 RECT 8.185 1.395 8.33 1.645 ;
 RECT 8.185 1.155 8.615 1.395 ;
 RECT 8.185 1.08 8.33 1.155 ;
 RECT 4.43 1.585 4.57 1.645 ;
 RECT 8.19 0.625 8.33 0.94 ;
 RECT 2.55 1.585 2.69 1.64 ;
 RECT 1.61 1.585 1.75 1.64 ;
 RECT 1.61 1.64 3.63 1.645 ;
 RECT 3.49 1.78 5.59 1.785 ;
 RECT 7.25 1.78 8.33 1.785 ;
 RECT 5.37 1.585 5.51 1.64 ;
 RECT 6.31 1.585 6.45 1.64 ;
 RECT 5.37 1.64 7.39 1.645 ;
 RECT 7.25 0.64 7.39 0.94 ;
 RECT 3.49 1.785 3.63 2.075 ;
 RECT 7.25 1.785 7.39 2.075 ;
 RECT 6.31 0.625 6.45 0.94 ;
 RECT 5.37 0.64 5.51 0.94 ;
 RECT 4.43 0.625 4.57 0.94 ;
 RECT 3.49 0.64 3.63 0.94 ;
 RECT 2.55 0.625 2.69 0.94 ;
 RECT 1.61 0.64 1.8 0.87 ;
 RECT 1.66 0.87 1.8 0.94 ;
 RECT 3.49 1.535 3.63 1.64 ;
 RECT 7.25 1.535 7.39 1.64 ;
 RECT 1.66 0.94 8.33 1.08 ;
 RECT 2.55 1.78 2.69 2.335 ;
 RECT 6.31 1.78 6.45 2.335 ;
 RECT 1.61 1.78 1.75 2.335 ;
 RECT 5.37 1.785 5.51 2.335 ;
 RECT 4.43 1.785 4.57 2.335 ;
 RECT 8.19 1.785 8.33 2.335 ;
 END
 ANTENNADIFFAREA 4.592 ;
 END Z

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.28 2.96 ;
 RECT 8.595 2.135 8.8 2.275 ;
 RECT 3.02 2.23 3.16 2.8 ;
 RECT 6.78 2.23 6.92 2.8 ;
 RECT 8.595 2.275 8.735 2.8 ;
 RECT 4.9 2.3 5.04 2.8 ;
 RECT 1.14 1.95 1.28 2.8 ;
 RECT 8.93 2.415 9.07 2.8 ;
 RECT 0.2 2 0.34 2.8 ;
 RECT 8.66 1.89 8.8 2.135 ;
 RECT 3.96 2.04 4.1 2.8 ;
 RECT 7.72 2.04 7.86 2.8 ;
 RECT 2.08 2.06 2.22 2.8 ;
 RECT 5.84 2.06 5.98 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 7.035 0.335 7.135 1.185 ;
 RECT 6.885 1.185 7.135 1.415 ;
 RECT 7.035 1.415 7.135 2.79 ;
 RECT 4.685 0.335 4.785 1.185 ;
 RECT 4.53 1.185 4.785 1.415 ;
 RECT 4.685 1.415 4.785 2.79 ;
 RECT 4.215 0.335 4.315 1.185 ;
 RECT 4.215 1.415 4.315 2.79 ;
 RECT 4.12 1.185 4.35 1.415 ;
 RECT 1.865 0.335 1.965 1.185 ;
 RECT 1.865 1.415 1.965 2.79 ;
 RECT 1.78 1.185 2.01 1.415 ;
 RECT 2.805 0.335 2.905 1.185 ;
 RECT 2.65 1.185 2.905 1.415 ;
 RECT 2.805 1.415 2.905 2.79 ;
 RECT 6.565 0.335 6.665 1.185 ;
 RECT 6.41 1.185 6.665 1.415 ;
 RECT 6.565 1.415 6.665 2.79 ;
 RECT 0.35 1.165 1.025 1.395 ;
 RECT 0.455 0.395 0.555 1.165 ;
 RECT 0.455 1.395 0.555 2.79 ;
 RECT 0.925 0.395 1.025 1.165 ;
 RECT 0.925 1.395 1.025 2.79 ;
 RECT 2.335 0.335 2.435 1.185 ;
 RECT 2.335 1.415 2.435 2.79 ;
 RECT 2.225 1.185 2.455 1.415 ;
 RECT 5.625 0.335 5.725 1.185 ;
 RECT 5.625 1.415 5.725 2.79 ;
 RECT 5.54 1.185 5.77 1.415 ;
 RECT 5.155 0.335 5.255 1.185 ;
 RECT 5.155 1.415 5.255 2.79 ;
 RECT 5.09 1.185 5.32 1.415 ;
 RECT 7.81 1.185 8.075 1.265 ;
 RECT 7.975 0.335 8.075 1.185 ;
 RECT 7.81 1.365 8.075 1.415 ;
 RECT 7.975 1.415 8.075 2.79 ;
 RECT 8.445 0.335 8.545 1.265 ;
 RECT 8.445 1.365 8.545 2.79 ;
 RECT 7.81 1.265 8.545 1.365 ;
 RECT 1.395 0.335 1.495 1.19 ;
 RECT 1.395 1.42 1.495 2.79 ;
 RECT 1.335 1.19 1.565 1.42 ;
 RECT 6.095 0.335 6.195 1.185 ;
 RECT 6.095 1.415 6.195 2.79 ;
 RECT 5.985 1.185 6.215 1.415 ;
 RECT 7.505 0.335 7.605 1.185 ;
 RECT 7.37 1.185 7.605 1.415 ;
 RECT 7.505 1.415 7.605 2.79 ;
 RECT 3.745 0.335 3.845 1.185 ;
 RECT 3.745 1.415 3.845 2.79 ;
 RECT 3.71 1.185 3.94 1.415 ;
 RECT 3.275 0.335 3.375 1.185 ;
 RECT 3.275 1.185 3.53 1.415 ;
 RECT 3.275 1.415 3.375 2.79 ;
 LAYER CO ;
 RECT 5.14 1.235 5.27 1.365 ;
 RECT 2.085 2.11 2.215 2.24 ;
 RECT 2.275 1.235 2.405 1.365 ;
 RECT 0.755 1.215 0.885 1.345 ;
 RECT 4.435 2.155 4.565 2.285 ;
 RECT 4.435 1.895 4.565 2.025 ;
 RECT 0.205 2.315 0.335 2.445 ;
 RECT 1.145 2.31 1.275 2.44 ;
 RECT 0.4 1.215 0.53 1.345 ;
 RECT 5.59 1.235 5.72 1.365 ;
 RECT 6.315 2.155 6.445 2.285 ;
 RECT 5.845 2.11 5.975 2.24 ;
 RECT 8.935 0.2 9.065 0.33 ;
 RECT 7.86 1.235 7.99 1.365 ;
 RECT 3.495 0.69 3.625 0.82 ;
 RECT 1.615 0.69 1.745 0.82 ;
 RECT 2.085 2.38 2.215 2.51 ;
 RECT 2.555 0.675 2.685 0.805 ;
 RECT 2.085 0.59 2.215 0.72 ;
 RECT 6.785 2.355 6.915 2.485 ;
 RECT 8.935 2.465 9.065 2.595 ;
 RECT 0.205 0.63 0.335 0.76 ;
 RECT 0.205 2.05 0.335 2.18 ;
 RECT 6.035 1.235 6.165 1.365 ;
 RECT 5.845 2.38 5.975 2.51 ;
 RECT 7.255 1.895 7.385 2.025 ;
 RECT 1.145 2 1.275 2.13 ;
 RECT 4.905 2.4 5.035 2.53 ;
 RECT 8.665 1.94 8.795 2.07 ;
 RECT 8.665 0.76 8.795 0.89 ;
 RECT 4.435 0.675 4.565 0.805 ;
 RECT 4.435 1.635 4.565 1.765 ;
 RECT 3.965 0.59 4.095 0.72 ;
 RECT 3.495 1.895 3.625 2.025 ;
 RECT 3.495 1.585 3.625 1.715 ;
 RECT 8.195 0.675 8.325 0.805 ;
 RECT 7.725 2.36 7.855 2.49 ;
 RECT 4.905 0.565 5.035 0.695 ;
 RECT 6.315 1.635 6.445 1.765 ;
 RECT 8.195 1.895 8.325 2.025 ;
 RECT 3.76 1.235 3.89 1.365 ;
 RECT 3.35 1.235 3.48 1.365 ;
 RECT 7.255 0.69 7.385 0.82 ;
 RECT 5.375 1.635 5.505 1.765 ;
 RECT 6.46 1.235 6.59 1.365 ;
 RECT 3.965 2.09 4.095 2.22 ;
 RECT 1.615 2.155 1.745 2.285 ;
 RECT 1.615 1.635 1.745 1.765 ;
 RECT 1.615 1.895 1.745 2.025 ;
 RECT 2.7 1.235 2.83 1.365 ;
 RECT 7.42 1.235 7.55 1.365 ;
 RECT 6.935 1.235 7.065 1.365 ;
 RECT 5.845 0.59 5.975 0.72 ;
 RECT 7.255 1.585 7.385 1.715 ;
 RECT 6.785 0.59 6.915 0.72 ;
 RECT 5.375 0.69 5.505 0.82 ;
 RECT 7.725 0.59 7.855 0.72 ;
 RECT 8.195 1.635 8.325 1.765 ;
 RECT 5.375 2.155 5.505 2.285 ;
 RECT 6.315 1.895 6.445 2.025 ;
 RECT 0.675 0.63 0.805 0.76 ;
 RECT 0.675 2.05 0.805 2.18 ;
 RECT 6.315 0.675 6.445 0.805 ;
 RECT 7.725 2.09 7.855 2.22 ;
 RECT 3.025 0.59 3.155 0.72 ;
 RECT 3.025 2.355 3.155 2.485 ;
 RECT 2.555 2.155 2.685 2.285 ;
 RECT 2.555 1.635 2.685 1.765 ;
 RECT 2.555 1.895 2.685 2.025 ;
 RECT 3.965 2.36 4.095 2.49 ;
 RECT 4.58 1.235 4.71 1.365 ;
 RECT 4.17 1.235 4.3 1.365 ;
 RECT 1.145 0.555 1.275 0.685 ;
 RECT 5.375 1.895 5.505 2.025 ;
 RECT 1.385 1.24 1.515 1.37 ;
 RECT 1.83 1.235 1.96 1.365 ;
 RECT 8.195 2.155 8.325 2.285 ;
 LAYER M1 ;
 RECT 6.885 1.23 7.115 1.37 ;
 RECT 7.37 1.23 7.6 1.37 ;
 RECT 6.41 1.23 6.64 1.37 ;
 RECT 5.985 1.23 6.215 1.37 ;
 RECT 5.54 1.23 5.77 1.37 ;
 RECT 5.09 1.23 5.32 1.37 ;
 RECT 4.53 1.23 4.76 1.37 ;
 RECT 4.12 1.23 4.35 1.37 ;
 RECT 3.71 1.23 3.94 1.37 ;
 RECT 3.3 1.23 3.53 1.37 ;
 RECT 2.65 1.23 2.88 1.37 ;
 RECT 2.225 1.23 2.455 1.37 ;
 RECT 1.78 1.23 2.01 1.37 ;
 RECT 0.67 0.88 1.435 1.02 ;
 RECT 0.67 1.54 1.435 1.68 ;
 RECT 1.295 1.02 1.435 1.365 ;
 RECT 1.295 1.19 1.435 1.54 ;
 RECT 1.38 1.19 1.52 1.42 ;
 RECT 0.67 2 0.81 2.23 ;
 RECT 0.67 0.58 0.81 1.02 ;
 RECT 0.67 1.68 0.81 2.07 ;
 RECT 7.81 1.23 8.04 1.37 ;
 RECT 1.44 1.23 8.02 1.37 ;
 END
END NBUFFX16

MACRO NBUFFX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 1.92 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 1.92 2.96 ;
 RECT 1.555 2.48 1.695 2.8 ;
 RECT 1.095 1.91 1.235 2.8 ;
 RECT 0.115 1.91 0.255 2.8 ;
 END
 END VDD

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 1.48 1.34 1.72 ;
 RECT 1.17 1.17 1.4 1.31 ;
 RECT 1.2 1.31 1.34 1.48 ;
 END
 ANTENNAGATEAREA 0.083 ;
 END INP

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 1.92 0.08 ;
 RECT 1.565 0.08 1.705 0.465 ;
 RECT 1.095 0.08 1.235 0.715 ;
 RECT 0.115 0.08 0.255 0.73 ;
 END
 END VSS

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.395 1.545 0.745 1.685 ;
 RECT 0.395 0.975 0.535 1.545 ;
 RECT 0.395 0.835 0.745 0.975 ;
 RECT 0.605 2.105 0.92 2.36 ;
 RECT 0.605 0.57 0.745 0.835 ;
 RECT 0.605 1.685 0.745 2.105 ;
 END
 ANTENNADIFFAREA 0.636 ;
 END Z

 OBS
 LAYER PO ;
 RECT 0.66 1.12 0.98 1.125 ;
 RECT 0.88 0.315 0.98 1.12 ;
 RECT 0.66 1.225 0.98 1.35 ;
 RECT 0.88 1.35 0.98 2.74 ;
 RECT 0.37 0.315 0.47 1.125 ;
 RECT 0.37 1.225 0.47 2.74 ;
 RECT 0.37 1.125 0.98 1.225 ;
 RECT 1.35 0.44 1.45 1.125 ;
 RECT 1.17 1.125 1.45 1.355 ;
 RECT 1.35 1.355 1.45 2.24 ;
 LAYER CO ;
 RECT 0.71 1.17 0.84 1.3 ;
 RECT 1.1 1.96 1.23 2.09 ;
 RECT 0.61 1.645 0.74 1.775 ;
 RECT 0.61 1.95 0.74 2.08 ;
 RECT 1.1 0.535 1.23 0.665 ;
 RECT 0.61 1.645 0.74 1.775 ;
 RECT 0.12 0.55 0.25 0.68 ;
 RECT 0.61 0.62 0.74 0.75 ;
 RECT 0.12 1.96 0.25 2.09 ;
 RECT 1.56 2.55 1.69 2.68 ;
 RECT 1.57 0.235 1.7 0.365 ;
 RECT 1.57 0.755 1.7 0.885 ;
 RECT 1.22 1.175 1.35 1.305 ;
 RECT 1.57 1.69 1.7 1.82 ;
 LAYER M1 ;
 RECT 0.71 1.12 1.025 1.26 ;
 RECT 0.885 0.995 1.025 1.12 ;
 RECT 0.705 1.12 0.845 1.35 ;
 RECT 0.885 0.855 1.705 0.995 ;
 RECT 1.565 0.7 1.705 1.725 ;
 RECT 1.565 1.64 1.705 1.87 ;
 END
END NBUFFX2

MACRO NBUFFX32
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 19.2 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 19.2 0.08 ;
 RECT 18.26 0.66 18.585 0.8 ;
 RECT 8.09 0.08 8.23 0.75 ;
 RECT 14.685 0.08 14.825 0.75 ;
 RECT 18.715 0.08 18.855 0.4 ;
 RECT 18.26 0.08 18.4 0.66 ;
 RECT 9.03 0.08 9.17 0.77 ;
 RECT 1.5 0.08 1.64 0.77 ;
 RECT 2.44 0.08 2.58 0.77 ;
 RECT 0.655 0.08 0.795 0.735 ;
 RECT 3.38 0.08 3.52 0.77 ;
 RECT 4.32 0.08 4.46 0.77 ;
 RECT 5.27 0.08 5.41 0.77 ;
 RECT 6.21 0.08 6.35 0.77 ;
 RECT 7.15 0.08 7.29 0.77 ;
 RECT 10.91 0.08 11.05 0.77 ;
 RECT 9.97 0.08 10.11 0.77 ;
 RECT 12.805 0.08 12.945 0.77 ;
 RECT 13.745 0.08 13.885 0.77 ;
 RECT 11.865 0.08 12.005 0.77 ;
 RECT 15.625 0.08 15.765 0.77 ;
 RECT 16.565 0.08 16.705 0.77 ;
 RECT 17.505 0.08 17.645 0.77 ;
 RECT 18.445 0.8 18.585 0.92 ;
 END
 END VSS

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 17.035 1.785 17.175 2.075 ;
 RECT 17.975 1.785 18.115 2.335 ;
 RECT 15.155 1.785 15.295 2.335 ;
 RECT 13.275 1.785 13.415 2.075 ;
 RECT 14.215 1.785 14.355 2.335 ;
 RECT 7.62 1.785 7.76 2.335 ;
 RECT 8.56 1.785 8.7 2.335 ;
 RECT 6.68 1.785 6.82 2.075 ;
 RECT 13.275 1.78 15.375 1.785 ;
 RECT 16.095 1.78 16.235 2.335 ;
 RECT 17.035 1.78 18.175 1.785 ;
 RECT 12.335 1.78 12.475 2.335 ;
 RECT 11.395 1.78 11.535 2.335 ;
 RECT 6.68 1.78 8.78 1.785 ;
 RECT 10.44 1.78 10.58 2.075 ;
 RECT 9.5 1.78 9.64 2.335 ;
 RECT 3.85 1.78 3.99 2.075 ;
 RECT 5.74 1.78 5.88 2.335 ;
 RECT 4.8 1.78 4.94 2.335 ;
 RECT 3.85 1.645 18.175 1.78 ;
 RECT 8.56 1.64 13.415 1.645 ;
 RECT 17.975 1.585 18.175 1.645 ;
 RECT 15.155 1.585 15.295 1.64 ;
 RECT 16.095 1.585 16.235 1.64 ;
 RECT 17.035 1.535 17.175 1.64 ;
 RECT 15.155 1.64 17.175 1.645 ;
 RECT 14.215 1.585 14.355 1.645 ;
 RECT 12.335 1.585 12.475 1.64 ;
 RECT 11.395 1.585 11.535 1.64 ;
 RECT 13.275 1.535 13.415 1.64 ;
 RECT 7.62 1.585 7.76 1.645 ;
 RECT 8.56 1.585 8.7 1.64 ;
 RECT 9.5 1.585 9.64 1.64 ;
 RECT 10.44 1.535 10.58 1.64 ;
 RECT 5.74 1.585 5.88 1.64 ;
 RECT 4.8 1.585 4.94 1.64 ;
 RECT 3.85 1.535 3.99 1.64 ;
 RECT 6.68 1.535 6.82 1.64 ;
 RECT 3.85 1.64 6.82 1.645 ;
 RECT 18.035 1.4 18.175 1.585 ;
 RECT 18.035 1.16 18.53 1.4 ;
 RECT 18.035 1.08 18.175 1.16 ;
 RECT 3.85 0.94 18.175 1.08 ;
 RECT 9.5 0.625 9.64 0.94 ;
 RECT 7.62 0.625 7.76 0.94 ;
 RECT 5.74 0.625 5.88 0.94 ;
 RECT 4.8 0.64 4.99 0.94 ;
 RECT 10.44 0.64 10.58 0.94 ;
 RECT 8.56 0.64 8.7 0.94 ;
 RECT 6.68 0.64 6.82 0.94 ;
 RECT 3.85 0.64 3.99 0.94 ;
 RECT 14.215 0.625 14.355 0.94 ;
 RECT 12.335 0.625 12.475 0.94 ;
 RECT 11.395 0.64 11.585 0.94 ;
 RECT 13.275 0.64 13.415 0.94 ;
 RECT 17.975 0.625 18.115 0.94 ;
 RECT 16.095 0.625 16.235 0.94 ;
 RECT 17.035 0.64 17.175 0.94 ;
 RECT 15.155 0.64 15.295 0.94 ;
 END
 ANTENNADIFFAREA 9.184 ;
 END Z

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.305 1.16 0.61 1.4 ;
 END
 ANTENNAGATEAREA 0.081 ;
 END INP

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 19.2 2.96 ;
 RECT 18.38 2.135 18.585 2.275 ;
 RECT 1.5 2.23 1.64 2.8 ;
 RECT 0.655 1.82 0.795 2.8 ;
 RECT 3.38 2.23 3.52 2.8 ;
 RECT 6.21 2.23 6.35 2.8 ;
 RECT 8.09 2.3 8.23 2.8 ;
 RECT 9.97 2.23 10.11 2.8 ;
 RECT 12.805 2.23 12.945 2.8 ;
 RECT 14.685 2.3 14.825 2.8 ;
 RECT 16.565 2.23 16.705 2.8 ;
 RECT 18.38 2.275 18.52 2.8 ;
 RECT 18.715 2.415 18.855 2.8 ;
 RECT 18.445 1.865 18.585 2.135 ;
 RECT 2.44 2.06 2.58 2.8 ;
 RECT 4.32 2.04 4.46 2.8 ;
 RECT 5.27 2.06 5.41 2.8 ;
 RECT 7.15 2.04 7.29 2.8 ;
 RECT 10.91 2.04 11.05 2.8 ;
 RECT 9.03 2.06 9.17 2.8 ;
 RECT 11.865 2.06 12.005 2.8 ;
 RECT 13.745 2.04 13.885 2.8 ;
 RECT 15.625 2.06 15.765 2.8 ;
 RECT 17.505 2.04 17.645 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 13.495 1.185 13.725 1.415 ;
 RECT 11.18 0.335 11.28 1.19 ;
 RECT 11.18 1.42 11.28 2.79 ;
 RECT 11.12 1.19 11.35 1.42 ;
 RECT 14 0.335 14.1 1.185 ;
 RECT 14 1.415 14.1 2.79 ;
 RECT 13.905 1.185 14.135 1.415 ;
 RECT 16.35 0.335 16.45 1.185 ;
 RECT 16.195 1.185 16.45 1.415 ;
 RECT 16.35 1.415 16.45 2.79 ;
 RECT 17.76 0.335 17.86 1.185 ;
 RECT 17.76 1.415 17.86 2.79 ;
 RECT 18.23 0.335 18.33 1.265 ;
 RECT 18.23 1.365 18.33 2.79 ;
 RECT 17.665 1.185 17.895 1.265 ;
 RECT 17.665 1.365 17.895 1.415 ;
 RECT 17.665 1.265 18.33 1.365 ;
 RECT 9.755 0.335 9.855 1.185 ;
 RECT 9.6 1.185 9.855 1.415 ;
 RECT 9.755 1.415 9.855 2.79 ;
 RECT 12.59 0.335 12.69 1.185 ;
 RECT 12.435 1.185 12.69 1.415 ;
 RECT 12.59 1.415 12.69 2.79 ;
 RECT 9.285 0.335 9.385 1.185 ;
 RECT 9.285 1.415 9.385 2.79 ;
 RECT 9.175 1.185 9.405 1.415 ;
 RECT 6.465 0.335 6.565 1.185 ;
 RECT 6.465 1.185 6.72 1.415 ;
 RECT 6.465 1.415 6.565 2.79 ;
 RECT 4.585 0.335 4.685 1.19 ;
 RECT 4.585 1.42 4.685 2.79 ;
 RECT 4.525 1.19 4.755 1.42 ;
 RECT 5.055 0.335 5.155 1.185 ;
 RECT 5.055 1.415 5.155 2.79 ;
 RECT 4.97 1.185 5.2 1.415 ;
 RECT 16.82 0.335 16.92 1.185 ;
 RECT 16.82 1.185 17.075 1.415 ;
 RECT 16.82 1.415 16.92 2.79 ;
 RECT 10.225 0.335 10.325 1.185 ;
 RECT 10.225 1.185 10.48 1.415 ;
 RECT 10.225 1.415 10.325 2.79 ;
 RECT 6.935 0.335 7.035 1.185 ;
 RECT 6.935 1.415 7.035 2.79 ;
 RECT 6.9 1.185 7.13 1.415 ;
 RECT 8.815 0.335 8.915 1.185 ;
 RECT 8.815 1.415 8.915 2.79 ;
 RECT 8.73 1.185 8.96 1.415 ;
 RECT 15.88 0.335 15.98 1.185 ;
 RECT 15.88 1.415 15.98 2.79 ;
 RECT 15.77 1.185 16 1.415 ;
 RECT 0.44 0.335 0.54 1.165 ;
 RECT 0.305 1.165 0.54 1.395 ;
 RECT 0.44 1.395 0.54 2.32 ;
 RECT 13.06 0.335 13.16 1.185 ;
 RECT 13.06 1.185 13.315 1.415 ;
 RECT 13.06 1.415 13.16 2.79 ;
 RECT 14.47 0.335 14.57 1.185 ;
 RECT 14.315 1.185 14.57 1.415 ;
 RECT 14.47 1.415 14.57 2.79 ;
 RECT 5.995 0.335 6.095 1.185 ;
 RECT 5.84 1.185 6.095 1.415 ;
 RECT 5.995 1.415 6.095 2.79 ;
 RECT 8.345 0.335 8.445 1.185 ;
 RECT 8.345 1.415 8.445 2.79 ;
 RECT 8.28 1.185 8.51 1.415 ;
 RECT 5.525 0.335 5.625 1.185 ;
 RECT 5.525 1.415 5.625 2.79 ;
 RECT 5.415 1.185 5.645 1.415 ;
 RECT 10.695 0.335 10.795 1.185 ;
 RECT 10.695 1.415 10.795 2.79 ;
 RECT 10.66 1.185 10.89 1.415 ;
 RECT 1.755 0.335 1.855 1.185 ;
 RECT 1.755 1.415 1.855 2.79 ;
 RECT 1.68 1.185 1.91 1.415 ;
 RECT 7.875 0.335 7.975 1.185 ;
 RECT 7.72 1.185 7.975 1.415 ;
 RECT 7.875 1.415 7.975 2.79 ;
 RECT 0.91 0.335 1.01 1.165 ;
 RECT 0.735 1.165 1.01 1.395 ;
 RECT 0.91 1.395 1.01 2.79 ;
 RECT 2.695 0.335 2.795 1.185 ;
 RECT 2.695 1.415 2.795 2.79 ;
 RECT 2.585 1.185 2.815 1.415 ;
 RECT 3.165 0.335 3.265 1.185 ;
 RECT 3.01 1.185 3.265 1.415 ;
 RECT 3.165 1.415 3.265 2.79 ;
 RECT 7.405 0.335 7.505 1.185 ;
 RECT 7.405 1.415 7.505 2.79 ;
 RECT 7.31 1.185 7.54 1.415 ;
 RECT 4.105 0.335 4.205 1.185 ;
 RECT 4.105 1.415 4.205 2.79 ;
 RECT 4.07 1.185 4.3 1.415 ;
 RECT 17.29 0.335 17.39 1.185 ;
 RECT 17.29 1.415 17.39 2.79 ;
 RECT 17.255 1.185 17.485 1.415 ;
 RECT 15.41 0.335 15.51 1.185 ;
 RECT 15.41 1.415 15.51 2.79 ;
 RECT 15.325 1.185 15.555 1.415 ;
 RECT 2.225 0.335 2.325 1.185 ;
 RECT 2.225 1.415 2.325 2.79 ;
 RECT 2.14 1.185 2.37 1.415 ;
 RECT 3.635 0.335 3.735 1.185 ;
 RECT 3.635 1.185 3.89 1.415 ;
 RECT 3.635 1.415 3.735 2.79 ;
 RECT 11.65 0.335 11.75 1.185 ;
 RECT 11.65 1.415 11.75 2.79 ;
 RECT 11.565 1.185 11.795 1.415 ;
 RECT 14.94 0.335 15.04 1.185 ;
 RECT 14.94 1.415 15.04 2.79 ;
 RECT 14.875 1.185 15.105 1.415 ;
 RECT 12.12 0.335 12.22 1.185 ;
 RECT 12.12 1.415 12.22 2.79 ;
 RECT 12.01 1.185 12.24 1.415 ;
 RECT 13.53 0.335 13.63 1.185 ;
 RECT 13.53 1.415 13.63 2.79 ;
 LAYER CO ;
 RECT 7.36 1.235 7.49 1.365 ;
 RECT 5.465 1.235 5.595 1.365 ;
 RECT 7.625 2.155 7.755 2.285 ;
 RECT 4.805 2.155 4.935 2.285 ;
 RECT 9.035 0.59 9.165 0.72 ;
 RECT 6.215 2.355 6.345 2.485 ;
 RECT 7.625 0.675 7.755 0.805 ;
 RECT 9.035 2.11 9.165 2.24 ;
 RECT 10.71 1.235 10.84 1.365 ;
 RECT 7.625 1.635 7.755 1.765 ;
 RECT 8.095 0.565 8.225 0.695 ;
 RECT 10.915 2.09 11.045 2.22 ;
 RECT 5.275 2.38 5.405 2.51 ;
 RECT 7.625 1.895 7.755 2.025 ;
 RECT 9.975 0.59 10.105 0.72 ;
 RECT 18.72 0.2 18.85 0.33 ;
 RECT 18.72 2.465 18.85 2.595 ;
 RECT 14.69 2.4 14.82 2.53 ;
 RECT 9.505 1.895 9.635 2.025 ;
 RECT 15.63 2.11 15.76 2.24 ;
 RECT 11.87 2.38 12 2.51 ;
 RECT 9.225 1.235 9.355 1.365 ;
 RECT 10.445 0.69 10.575 0.82 ;
 RECT 4.805 1.895 4.935 2.025 ;
 RECT 9.65 1.235 9.78 1.365 ;
 RECT 6.215 0.59 6.345 0.72 ;
 RECT 8.095 2.4 8.225 2.53 ;
 RECT 15.16 2.155 15.29 2.285 ;
 RECT 5.745 1.895 5.875 2.025 ;
 RECT 0.19 0.555 0.32 0.685 ;
 RECT 0.66 1.87 0.79 2 ;
 RECT 11.87 0.59 12 0.72 ;
 RECT 13.28 0.69 13.41 0.82 ;
 RECT 17.305 1.235 17.435 1.365 ;
 RECT 12.06 1.235 12.19 1.365 ;
 RECT 15.82 1.235 15.95 1.365 ;
 RECT 0.19 1.87 0.32 2 ;
 RECT 0.355 1.215 0.485 1.345 ;
 RECT 2.915 1.895 3.045 2.025 ;
 RECT 2.445 0.59 2.575 0.72 ;
 RECT 2.635 1.235 2.765 1.365 ;
 RECT 11.615 1.235 11.745 1.365 ;
 RECT 2.915 2.155 3.045 2.285 ;
 RECT 1.975 0.69 2.105 0.82 ;
 RECT 13.75 2.09 13.88 2.22 ;
 RECT 17.98 0.675 18.11 0.805 ;
 RECT 16.895 1.235 17.025 1.365 ;
 RECT 12.485 1.235 12.615 1.365 ;
 RECT 13.955 1.235 14.085 1.365 ;
 RECT 17.04 1.895 17.17 2.025 ;
 RECT 16.1 1.635 16.23 1.765 ;
 RECT 17.715 1.235 17.845 1.365 ;
 RECT 17.98 1.635 18.11 1.765 ;
 RECT 12.34 1.895 12.47 2.025 ;
 RECT 6.95 1.235 7.08 1.365 ;
 RECT 9.505 1.635 9.635 1.765 ;
 RECT 8.78 1.235 8.91 1.365 ;
 RECT 7.155 2.09 7.285 2.22 ;
 RECT 5.275 2.11 5.405 2.24 ;
 RECT 5.89 1.235 6.02 1.365 ;
 RECT 5.275 0.59 5.405 0.72 ;
 RECT 8.33 1.235 8.46 1.365 ;
 RECT 10.445 1.585 10.575 1.715 ;
 RECT 9.505 0.675 9.635 0.805 ;
 RECT 7.155 2.36 7.285 2.49 ;
 RECT 7.155 0.59 7.285 0.72 ;
 RECT 6.685 0.69 6.815 0.82 ;
 RECT 5.02 1.235 5.15 1.365 ;
 RECT 10.915 0.59 11.045 0.72 ;
 RECT 4.575 1.235 4.705 1.365 ;
 RECT 0.66 2.355 0.79 2.485 ;
 RECT 1.505 2.355 1.635 2.485 ;
 RECT 5.745 1.635 5.875 1.765 ;
 RECT 8.565 1.895 8.695 2.025 ;
 RECT 4.325 0.59 4.455 0.72 ;
 RECT 10.915 2.36 11.045 2.49 ;
 RECT 8.565 2.155 8.695 2.285 ;
 RECT 10.445 1.895 10.575 2.025 ;
 RECT 6.685 1.585 6.815 1.715 ;
 RECT 3.385 2.355 3.515 2.485 ;
 RECT 3.385 0.59 3.515 0.72 ;
 RECT 4.805 0.69 4.935 0.82 ;
 RECT 6.54 1.235 6.67 1.365 ;
 RECT 1.975 2.155 2.105 2.285 ;
 RECT 3.855 1.895 3.985 2.025 ;
 RECT 1.73 1.235 1.86 1.365 ;
 RECT 3.06 1.235 3.19 1.365 ;
 RECT 9.035 2.38 9.165 2.51 ;
 RECT 8.565 1.635 8.695 1.765 ;
 RECT 1.13 0.69 1.26 0.82 ;
 RECT 5.745 2.155 5.875 2.285 ;
 RECT 8.565 0.69 8.695 0.82 ;
 RECT 1.975 1.635 2.105 1.765 ;
 RECT 2.445 2.11 2.575 2.24 ;
 RECT 4.805 1.635 4.935 1.765 ;
 RECT 2.915 1.635 3.045 1.765 ;
 RECT 3.855 1.585 3.985 1.715 ;
 RECT 2.19 1.235 2.32 1.365 ;
 RECT 2.915 0.675 3.045 0.805 ;
 RECT 11.17 1.235 11.3 1.365 ;
 RECT 0.785 1.215 0.915 1.345 ;
 RECT 12.34 0.675 12.47 0.805 ;
 RECT 7.77 1.235 7.9 1.365 ;
 RECT 9.505 2.155 9.635 2.285 ;
 RECT 1.13 1.635 1.26 1.765 ;
 RECT 1.13 2.155 1.26 2.285 ;
 RECT 1.13 1.895 1.26 2.025 ;
 RECT 1.505 0.59 1.635 0.72 ;
 RECT 3.71 1.235 3.84 1.365 ;
 RECT 4.325 2.09 4.455 2.22 ;
 RECT 1.975 1.895 2.105 2.025 ;
 RECT 2.445 2.38 2.575 2.51 ;
 RECT 4.12 1.235 4.25 1.365 ;
 RECT 6.685 1.895 6.815 2.025 ;
 RECT 4.325 2.36 4.455 2.49 ;
 RECT 3.855 0.69 3.985 0.82 ;
 RECT 15.63 2.38 15.76 2.51 ;
 RECT 13.75 2.36 13.88 2.49 ;
 RECT 16.57 2.355 16.7 2.485 ;
 RECT 13.135 1.235 13.265 1.365 ;
 RECT 12.34 2.155 12.47 2.285 ;
 RECT 16.57 0.59 16.7 0.72 ;
 RECT 14.22 1.635 14.35 1.765 ;
 RECT 15.375 1.235 15.505 1.365 ;
 RECT 11.4 2.155 11.53 2.285 ;
 RECT 14.69 0.565 14.82 0.695 ;
 RECT 13.28 1.585 13.41 1.715 ;
 RECT 12.81 0.59 12.94 0.72 ;
 RECT 13.28 1.895 13.41 2.025 ;
 RECT 14.925 1.235 15.055 1.365 ;
 RECT 11.4 1.895 11.53 2.025 ;
 RECT 14.365 1.235 14.495 1.365 ;
 RECT 16.1 1.895 16.23 2.025 ;
 RECT 11.87 2.11 12 2.24 ;
 RECT 17.04 1.585 17.17 1.715 ;
 RECT 14.22 2.155 14.35 2.285 ;
 RECT 13.545 1.235 13.675 1.365 ;
 RECT 17.51 2.09 17.64 2.22 ;
 RECT 15.63 0.59 15.76 0.72 ;
 RECT 14.22 0.675 14.35 0.805 ;
 RECT 14.22 1.895 14.35 2.025 ;
 RECT 17.51 2.36 17.64 2.49 ;
 RECT 10.3 1.235 10.43 1.365 ;
 RECT 5.745 0.675 5.875 0.805 ;
 RECT 15.16 0.69 15.29 0.82 ;
 RECT 13.75 0.59 13.88 0.72 ;
 RECT 17.98 2.155 18.11 2.285 ;
 RECT 9.975 2.355 10.105 2.485 ;
 RECT 17.98 1.895 18.11 2.025 ;
 RECT 12.34 1.635 12.47 1.765 ;
 RECT 17.04 0.69 17.17 0.82 ;
 RECT 16.245 1.235 16.375 1.365 ;
 RECT 18.45 0.74 18.58 0.87 ;
 RECT 12.81 2.355 12.94 2.485 ;
 RECT 15.16 1.895 15.29 2.025 ;
 RECT 16.1 2.155 16.23 2.285 ;
 RECT 18.45 1.915 18.58 2.045 ;
 RECT 16.1 0.675 16.23 0.805 ;
 RECT 17.51 0.59 17.64 0.72 ;
 RECT 0.66 0.555 0.79 0.685 ;
 RECT 11.4 0.69 11.53 0.82 ;
 RECT 15.16 1.635 15.29 1.765 ;
 RECT 11.4 1.635 11.53 1.765 ;
 LAYER M1 ;
 RECT 1.125 1.37 1.265 2.335 ;
 RECT 1.125 0.64 1.265 1.23 ;
 RECT 1.125 1.23 3.24 1.37 ;
 RECT 0.185 0.505 0.325 0.88 ;
 RECT 0.185 1.68 0.325 2.05 ;
 RECT 0.78 1.165 0.925 1.395 ;
 RECT 0.785 1.395 0.925 1.54 ;
 RECT 0.785 1.02 0.925 1.165 ;
 RECT 0.185 0.88 0.925 1.02 ;
 RECT 0.185 1.54 0.925 1.68 ;
 RECT 1.97 1.64 3.71 1.78 ;
 RECT 1.97 0.94 3.71 1.075 ;
 RECT 2.91 0.935 3.71 0.94 ;
 RECT 3.57 1.075 3.71 1.23 ;
 RECT 3.57 1.37 3.71 1.64 ;
 RECT 2.91 1.78 3.05 2.335 ;
 RECT 2.91 1.585 3.05 1.64 ;
 RECT 1.97 1.075 3.05 1.08 ;
 RECT 2.91 0.625 3.05 0.935 ;
 RECT 1.97 1.78 2.11 2.335 ;
 RECT 1.97 1.585 2.11 1.64 ;
 RECT 1.97 0.64 2.11 0.94 ;
 RECT 3.57 1.23 17.895 1.37 ;
 END
END NBUFFX32

MACRO NBUFFX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 3.165 0.08 3.305 0.4 ;
 RECT 1.485 0.08 1.625 0.77 ;
 RECT 2.425 0.08 2.565 0.77 ;
 RECT 0.175 0.08 0.315 0.785 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.18 1.15 0.535 1.405 ;
 END
 ANTENNAGATEAREA 0.083 ;
 END INP

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.205 0.94 3.035 1.08 ;
 RECT 1.015 0.745 1.345 0.885 ;
 RECT 1.015 1.715 2.095 1.855 ;
 RECT 2.895 1.115 3.355 1.45 ;
 RECT 1.955 0.625 2.095 0.94 ;
 RECT 2.895 1.08 3.035 1.115 ;
 RECT 2.895 0.695 3.035 0.94 ;
 RECT 1.955 1.86 3.035 2 ;
 RECT 1.205 0.885 1.345 0.94 ;
 RECT 1.015 0.64 1.155 0.745 ;
 RECT 1.955 1.855 2.095 1.86 ;
 RECT 1.015 1.855 1.155 2.31 ;
 RECT 1.955 2 2.095 2.31 ;
 RECT 2.895 2 3.035 2.04 ;
 RECT 2.895 1.45 3.035 1.86 ;
 END
 ANTENNADIFFAREA 1.408 ;
 END Z

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 2.425 2.345 2.565 2.8 ;
 RECT 1.485 2.065 1.625 2.8 ;
 RECT 3.165 2.415 3.305 2.8 ;
 RECT 0.175 1.835 0.315 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 0.43 0.385 0.53 1.185 ;
 RECT 0.265 1.185 0.53 1.415 ;
 RECT 0.43 1.415 0.53 2.425 ;
 RECT 1.74 0.335 1.84 1.185 ;
 RECT 1.74 1.415 1.84 2.79 ;
 RECT 1.655 1.185 1.885 1.415 ;
 RECT 2.68 0.335 2.78 1.185 ;
 RECT 2.525 1.185 2.78 1.415 ;
 RECT 2.68 1.415 2.78 2.79 ;
 RECT 2.21 0.335 2.31 1.185 ;
 RECT 2.21 1.415 2.31 2.79 ;
 RECT 2.1 1.185 2.33 1.415 ;
 RECT 1.27 0.335 1.37 1.185 ;
 RECT 1.27 1.415 1.37 2.79 ;
 RECT 1.205 1.185 1.435 1.415 ;
 LAYER CO ;
 RECT 0.315 1.235 0.445 1.365 ;
 RECT 0.65 0.605 0.78 0.735 ;
 RECT 0.18 1.885 0.31 2.015 ;
 RECT 0.18 0.605 0.31 0.735 ;
 RECT 0.65 1.875 0.78 2.005 ;
 RECT 1.49 0.59 1.62 0.72 ;
 RECT 1.49 2.425 1.62 2.555 ;
 RECT 1.255 1.235 1.385 1.365 ;
 RECT 1.705 1.235 1.835 1.365 ;
 RECT 1.02 2.13 1.15 2.26 ;
 RECT 3.17 0.2 3.3 0.33 ;
 RECT 2.43 2.44 2.56 2.57 ;
 RECT 2.575 1.235 2.705 1.365 ;
 RECT 2.9 1.86 3.03 1.99 ;
 RECT 1.96 1.86 2.09 1.99 ;
 RECT 2.15 1.235 2.28 1.365 ;
 RECT 1.02 1.86 1.15 1.99 ;
 RECT 1.49 2.115 1.62 2.245 ;
 RECT 2.9 0.76 3.03 0.89 ;
 RECT 3.17 2.465 3.3 2.595 ;
 RECT 1.02 0.69 1.15 0.82 ;
 RECT 1.96 2.13 2.09 2.26 ;
 RECT 1.96 0.675 2.09 0.805 ;
 RECT 2.43 0.59 2.56 0.72 ;
 LAYER M1 ;
 RECT 1.655 1.23 1.885 1.37 ;
 RECT 0.72 1.23 1.325 1.37 ;
 RECT 1.205 1.23 1.435 1.37 ;
 RECT 0.645 1.825 0.785 2.055 ;
 RECT 0.645 0.555 0.785 0.785 ;
 RECT 0.645 1.695 0.785 2 ;
 RECT 0.645 0.715 0.785 0.87 ;
 RECT 0.645 1.555 0.855 1.695 ;
 RECT 0.645 0.87 0.86 1.01 ;
 RECT 0.715 1 0.855 1.555 ;
 RECT 0.72 1.01 0.86 1.23 ;
 RECT 2.1 1.23 2.33 1.37 ;
 RECT 2.525 1.23 2.755 1.37 ;
 RECT 1.315 1.23 2.69 1.37 ;
 END
END NBUFFX4

MACRO NBUFFX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 4.315 0.64 4.64 0.78 ;
 RECT 4.315 0.08 4.455 0.64 ;
 RECT 0.74 0.08 0.88 0.755 ;
 RECT 4.77 0.08 4.91 0.4 ;
 RECT 3.56 0.08 3.7 0.77 ;
 RECT 4.5 0.78 4.64 0.94 ;
 RECT 1.68 0.08 1.82 0.745 ;
 RECT 2.62 0.08 2.76 0.735 ;
 END
 END VSS

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.09 1.08 4.23 1.27 ;
 RECT 4.03 0.625 4.17 0.94 ;
 RECT 3.09 0.64 3.23 0.94 ;
 RECT 1.21 0.89 2.76 0.94 ;
 RECT 1.21 1.585 1.35 1.64 ;
 RECT 2.15 0.625 2.29 0.89 ;
 RECT 1.21 0.64 1.35 0.89 ;
 RECT 4.025 1.63 4.59 1.645 ;
 RECT 4.03 1.585 4.59 1.63 ;
 RECT 4.09 1.27 4.59 1.585 ;
 RECT 3.09 1.535 3.23 1.64 ;
 RECT 2.62 1.03 4.23 1.08 ;
 RECT 2.15 1.585 2.29 1.64 ;
 RECT 1.21 1.77 4.17 1.78 ;
 RECT 2.15 1.03 2.29 1.035 ;
 RECT 1.21 0.94 4.23 1.03 ;
 RECT 3.09 1.78 4.17 1.785 ;
 RECT 3.09 1.785 3.23 2.075 ;
 RECT 1.21 1.645 4.59 1.725 ;
 RECT 1.21 1.64 3.23 1.645 ;
 RECT 2.15 1.78 2.29 2.335 ;
 RECT 4.03 1.785 4.17 2.335 ;
 RECT 1.21 1.78 1.35 2.335 ;
 RECT 1.21 1.725 4.23 1.77 ;
 END
 ANTENNADIFFAREA 2.296 ;
 END Z

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 4.435 2.135 4.64 2.275 ;
 RECT 4.435 2.275 4.575 2.8 ;
 RECT 2.62 2.23 2.76 2.8 ;
 RECT 0.74 2.3 0.88 2.8 ;
 RECT 4.77 2.415 4.91 2.8 ;
 RECT 4.5 1.865 4.64 2.135 ;
 RECT 1.68 2.06 1.82 2.8 ;
 RECT 3.56 2.04 3.7 2.8 ;
 END
 END VDD

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.325 1.18 0.625 1.6 ;
 RECT 0.36 1.175 0.59 1.18 ;
 END
 ANTENNAGATEAREA 0.155 ;
 END INP

 OBS
 LAYER PO ;
 RECT 3.815 0.335 3.915 1.185 ;
 RECT 3.815 1.415 3.915 2.79 ;
 RECT 4.285 0.335 4.385 1.265 ;
 RECT 4.285 1.365 4.385 2.79 ;
 RECT 3.72 1.185 3.95 1.265 ;
 RECT 3.72 1.365 3.95 1.415 ;
 RECT 3.72 1.265 4.385 1.365 ;
 RECT 3.345 0.335 3.445 1.185 ;
 RECT 3.345 1.415 3.445 2.79 ;
 RECT 3.31 1.185 3.54 1.415 ;
 RECT 2.875 0.335 2.975 1.185 ;
 RECT 2.875 1.185 3.13 1.415 ;
 RECT 2.875 1.415 2.975 2.79 ;
 RECT 1.465 0.335 1.565 1.17 ;
 RECT 1.465 1.4 1.565 2.79 ;
 RECT 1.38 1.17 1.61 1.4 ;
 RECT 2.405 0.335 2.505 1.185 ;
 RECT 2.25 1.185 2.505 1.415 ;
 RECT 2.405 1.415 2.505 2.79 ;
 RECT 1.935 0.335 2.035 1.185 ;
 RECT 1.935 1.415 2.035 2.79 ;
 RECT 1.825 1.185 2.055 1.415 ;
 RECT 0.995 0.335 1.095 1.14 ;
 RECT 0.995 1.37 1.095 2.79 ;
 RECT 0.91 1.14 1.14 1.37 ;
 RECT 0.525 0.335 0.625 1.13 ;
 RECT 0.36 1.13 0.625 1.36 ;
 RECT 0.525 1.36 0.625 2.79 ;
 LAYER CO ;
 RECT 3.095 1.895 3.225 2.025 ;
 RECT 4.505 1.915 4.635 2.045 ;
 RECT 3.095 1.585 3.225 1.715 ;
 RECT 3.565 2.36 3.695 2.49 ;
 RECT 3.77 1.235 3.9 1.365 ;
 RECT 3.36 1.235 3.49 1.365 ;
 RECT 2.95 1.235 3.08 1.365 ;
 RECT 0.745 0.565 0.875 0.695 ;
 RECT 0.96 1.19 1.09 1.32 ;
 RECT 1.43 1.22 1.56 1.35 ;
 RECT 2.3 1.235 2.43 1.365 ;
 RECT 1.685 2.11 1.815 2.24 ;
 RECT 1.875 1.235 2.005 1.365 ;
 RECT 3.095 0.69 3.225 0.82 ;
 RECT 1.215 0.69 1.345 0.82 ;
 RECT 1.685 2.38 1.815 2.51 ;
 RECT 2.155 0.675 2.285 0.805 ;
 RECT 1.685 0.555 1.815 0.685 ;
 RECT 1.215 2.155 1.345 2.285 ;
 RECT 1.215 1.635 1.345 1.765 ;
 RECT 1.215 1.895 1.345 2.025 ;
 RECT 2.155 2.155 2.285 2.285 ;
 RECT 2.155 1.635 2.285 1.765 ;
 RECT 2.155 1.895 2.285 2.025 ;
 RECT 0.41 1.18 0.54 1.31 ;
 RECT 4.035 2.155 4.165 2.285 ;
 RECT 4.035 1.895 4.165 2.025 ;
 RECT 0.745 2.4 0.875 2.53 ;
 RECT 0.275 0.725 0.405 0.855 ;
 RECT 0.275 2.05 0.405 2.18 ;
 RECT 3.565 2.09 3.695 2.22 ;
 RECT 2.625 0.555 2.755 0.685 ;
 RECT 2.625 2.355 2.755 2.485 ;
 RECT 4.775 0.2 4.905 0.33 ;
 RECT 4.505 0.76 4.635 0.89 ;
 RECT 4.035 0.675 4.165 0.805 ;
 RECT 4.035 1.635 4.165 1.765 ;
 RECT 4.775 2.465 4.905 2.595 ;
 RECT 3.565 0.59 3.695 0.72 ;
 LAYER M1 ;
 RECT 2.25 1.23 2.48 1.37 ;
 RECT 1.825 1.23 2.055 1.37 ;
 RECT 1.38 1.215 1.61 1.355 ;
 RECT 0.27 0.895 1.07 1.035 ;
 RECT 0.91 1.185 1.14 1.325 ;
 RECT 0.93 1.035 1.07 2.02 ;
 RECT 0.27 2.02 1.07 2.16 ;
 RECT 0.27 0.675 0.41 0.94 ;
 RECT 0.27 2 0.41 2.23 ;
 RECT 3.31 1.23 3.54 1.37 ;
 RECT 2.9 1.23 3.13 1.37 ;
 RECT 3.72 1.23 3.95 1.37 ;
 RECT 1.04 1.23 3.875 1.37 ;
 END
END NBUFFX8

MACRO NOR2X0
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 1.92 BY 2.88 ;
 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.185 1.08 1.43 1.21 ;
 RECT 0.715 1.21 1.43 1.36 ;
 RECT 1.185 0.255 1.325 1.08 ;
 RECT 0.715 1.36 0.855 2.28 ;
 END
 ANTENNADIFFAREA 0.318 ;
 END QN

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.535 0.68 1.04 1.065 ;
 END
 ANTENNAGATEAREA 0.101 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 1.92 2.96 ;
 RECT 1.655 1.42 1.795 2.8 ;
 RECT 0.3 1.495 0.44 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 1.92 0.08 ;
 RECT 0.715 0.08 0.855 0.505 ;
 RECT 1.655 0.08 1.795 0.555 ;
 RECT 0.255 0.08 0.395 0.755 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.11 2.28 1.515 2.66 ;
 END
 ANTENNAGATEAREA 0.101 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 0.97 0.915 1.07 2.435 ;
 RECT 0.97 0.105 1.07 0.685 ;
 RECT 0.81 0.685 1.07 0.915 ;
 RECT 1.44 0.105 1.54 2.35 ;
 RECT 1.31 2.35 1.54 2.58 ;
 LAYER CO ;
 RECT 1.66 1.805 1.79 1.935 ;
 RECT 0.72 2.07 0.85 2.2 ;
 RECT 0.72 1.81 0.85 1.94 ;
 RECT 1.36 2.4 1.49 2.53 ;
 RECT 1.66 1.54 1.79 1.67 ;
 RECT 0.305 2.065 0.435 2.195 ;
 RECT 1.66 0.325 1.79 0.455 ;
 RECT 0.72 0.325 0.85 0.455 ;
 RECT 1.19 0.325 1.32 0.455 ;
 RECT 0.26 0.315 0.39 0.445 ;
 RECT 0.305 1.805 0.435 1.935 ;
 RECT 0.86 0.735 0.99 0.865 ;
 RECT 0.305 1.545 0.435 1.675 ;
 RECT 0.72 1.545 0.85 1.675 ;
 RECT 0.26 0.575 0.39 0.705 ;
 END
END NOR2X0

MACRO NOR2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.24 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 0.8 1.1 1.08 ;
 END
 ANTENNAGATEAREA 0.14 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.24 2.96 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 1.71 1.495 1.85 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.24 0.08 ;
 RECT 0.77 0.08 0.91 0.62 ;
 RECT 1.71 0.08 1.85 0.6 ;
 RECT 0.31 0.08 0.45 0.755 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.535 0.745 1.88 1.08 ;
 END
 ANTENNAGATEAREA 0.14 ;
 END IN2

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.77 1.56 0.91 2.605 ;
 RECT 1.24 0.345 1.38 1.32 ;
 RECT 0.77 1.32 1.38 1.56 ;
 END
 ANTENNADIFFAREA 0.44 ;
 END QN

 OBS
 LAYER PO ;
 RECT 1.025 1.07 1.125 2.74 ;
 RECT 1.025 0.165 1.125 0.84 ;
 RECT 0.865 0.84 1.125 1.07 ;
 RECT 1.495 0.165 1.595 0.745 ;
 RECT 1.495 0.975 1.595 2.74 ;
 RECT 1.495 0.745 1.725 0.975 ;
 LAYER CO ;
 RECT 1.715 2.38 1.845 2.51 ;
 RECT 1.715 2.105 1.845 2.235 ;
 RECT 1.715 1.83 1.845 1.96 ;
 RECT 0.775 2.375 0.905 2.505 ;
 RECT 0.775 2.1 0.905 2.23 ;
 RECT 0.775 1.825 0.905 1.955 ;
 RECT 1.545 0.795 1.675 0.925 ;
 RECT 1.715 1.545 1.845 1.675 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 1.715 0.415 1.845 0.545 ;
 RECT 0.775 0.405 0.905 0.535 ;
 RECT 1.245 0.4 1.375 0.53 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 0.915 0.89 1.045 1.02 ;
 RECT 1.715 1.545 1.845 1.675 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 0.775 1.545 0.905 1.675 ;
 RECT 0.315 0.575 0.445 0.705 ;
 END
END NOR2X1

MACRO NOR2X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.28 0.675 2.52 0.99 ;
 END
 ANTENNAGATEAREA 0.28 ;
 END IN2

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 2.21 2.245 2.35 2.8 ;
 RECT 0.355 1.495 0.495 2.8 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.69 0.27 2.83 1.205 ;
 RECT 1.73 0.275 1.89 0.505 ;
 RECT 0.785 0.25 0.925 1.21 ;
 RECT 1.7 1.205 2.83 1.21 ;
 RECT 1.735 0.505 1.875 1.16 ;
 RECT 0.785 1.21 2.83 1.345 ;
 RECT 1.735 1.16 2.04 1.205 ;
 RECT 1.27 1.36 1.41 1.725 ;
 RECT 0.785 1.345 2.04 1.35 ;
 RECT 1.735 1.36 2.04 1.4 ;
 RECT 1.27 1.35 2.04 1.36 ;
 END
 ANTENNADIFFAREA 0.706 ;
 END QN

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 0.83 1.545 1.07 ;
 END
 ANTENNAGATEAREA 0.28 ;
 END IN1

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 1.27 0.08 1.41 0.505 ;
 RECT 2.21 0.08 2.35 0.535 ;
 RECT 0.31 0.08 0.45 0.755 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 1.32 0.83 1.625 0.895 ;
 RECT 1.32 0.995 1.625 1.07 ;
 RECT 1.04 0.895 1.625 0.995 ;
 RECT 1.04 0.105 1.14 0.895 ;
 RECT 1.04 0.995 1.14 2.74 ;
 RECT 1.525 0.105 1.625 0.83 ;
 RECT 1.525 1.07 1.625 2.74 ;
 RECT 2.315 0.745 2.575 0.805 ;
 RECT 2.475 0.105 2.575 0.745 ;
 RECT 2.315 0.905 2.575 0.975 ;
 RECT 2.475 0.975 2.575 2.74 ;
 RECT 1.995 0.105 2.095 0.805 ;
 RECT 1.995 0.805 2.585 0.905 ;
 RECT 1.995 0.905 2.095 2.74 ;
 LAYER CO ;
 RECT 2.695 0.335 2.825 0.465 ;
 RECT 2.695 1.915 2.825 2.045 ;
 RECT 0.79 0.325 0.92 0.455 ;
 RECT 1.745 1.915 1.875 2.045 ;
 RECT 0.79 1.915 0.92 2.045 ;
 RECT 1.275 1.545 1.405 1.675 ;
 RECT 1.745 0.325 1.875 0.455 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 1.275 0.325 1.405 0.455 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 1.375 0.89 1.505 1.02 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 2.215 0.325 2.345 0.455 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 2.365 0.795 2.495 0.925 ;
 RECT 2.215 2.37 2.345 2.5 ;
 RECT 0.315 0.315 0.445 0.445 ;
 LAYER M1 ;
 RECT 0.715 1.91 2.945 2.05 ;
 END
END NOR2X2

MACRO NOR2X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 2.32 0.08 2.46 0.505 ;
 RECT 1.345 0.08 1.485 0.505 ;
 RECT 3.26 0.08 3.4 0.555 ;
 RECT 0.31 0.08 0.45 0.755 ;
 RECT 4.22 0.08 4.36 0.555 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.28 0.68 2.645 1.06 ;
 END
 ANTENNAGATEAREA 0.56 ;
 END IN1

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.92 1.61 4.84 1.75 ;
 RECT 2.78 0.275 2.94 0.505 ;
 RECT 2.32 1.35 2.46 1.725 ;
 RECT 1.835 0.25 1.975 1.205 ;
 RECT 1.355 1.35 1.495 1.725 ;
 RECT 0.83 1.345 1.52 1.35 ;
 RECT 0.83 0.25 0.97 1.205 ;
 RECT 3.74 0.27 3.88 0.71 ;
 RECT 4.7 0.85 4.84 1.61 ;
 RECT 3.74 0.71 4.84 0.85 ;
 RECT 4.7 0.265 4.84 0.71 ;
 RECT 2.785 0.505 2.925 1.205 ;
 RECT 2.92 1.35 3.175 1.61 ;
 RECT 1.835 1.345 3.175 1.35 ;
 RECT 0.83 1.205 3.175 1.345 ;
 END
 ANTENNADIFFAREA 1.394 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 3.26 2.245 3.4 2.8 ;
 RECT 4.22 2.245 4.36 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.365 1.015 3.98 1.155 ;
 RECT 3.695 1.155 3.98 1.415 ;
 RECT 3.365 0.745 3.6 1.015 ;
 END
 ANTENNAGATEAREA 0.56 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 1.085 0.995 1.185 2.745 ;
 RECT 1.085 0.105 1.185 0.895 ;
 RECT 1.61 0.995 1.71 2.74 ;
 RECT 1.61 0.105 1.71 0.895 ;
 RECT 2.09 0.995 2.19 2.74 ;
 RECT 2.09 0.105 2.19 0.895 ;
 RECT 2.575 0.105 2.675 0.83 ;
 RECT 2.575 1.06 2.675 2.74 ;
 RECT 2.37 0.83 2.675 0.895 ;
 RECT 1.085 0.895 2.675 0.995 ;
 RECT 2.37 0.995 2.675 1.06 ;
 RECT 3.365 0.745 3.625 0.805 ;
 RECT 3.525 0.105 3.625 0.745 ;
 RECT 3.365 0.905 3.625 0.975 ;
 RECT 3.525 0.975 3.625 2.74 ;
 RECT 3.045 0.105 3.145 0.805 ;
 RECT 3.045 0.905 3.145 2.74 ;
 RECT 4.475 0.105 4.575 0.805 ;
 RECT 4.475 0.905 4.575 2.74 ;
 RECT 4 0.105 4.1 0.805 ;
 RECT 4 0.905 4.1 2.74 ;
 RECT 3.045 0.805 4.575 0.905 ;
 LAYER CO ;
 RECT 4.705 0.335 4.835 0.465 ;
 RECT 4.695 1.915 4.825 2.045 ;
 RECT 4.225 2.37 4.355 2.5 ;
 RECT 4.225 0.325 4.355 0.455 ;
 RECT 0.835 0.325 0.965 0.455 ;
 RECT 0.83 1.915 0.96 2.045 ;
 RECT 1.36 1.545 1.49 1.675 ;
 RECT 1.35 0.325 1.48 0.455 ;
 RECT 3.745 0.335 3.875 0.465 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 3.745 1.915 3.875 2.045 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 3.265 0.325 3.395 0.455 ;
 RECT 1.84 0.325 1.97 0.455 ;
 RECT 3.265 2.37 3.395 2.5 ;
 RECT 2.325 0.325 2.455 0.455 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 1.84 1.915 1.97 2.045 ;
 RECT 2.795 1.915 2.925 2.045 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 2.795 0.325 2.925 0.455 ;
 RECT 2.325 1.545 2.455 1.675 ;
 RECT 3.415 0.795 3.545 0.925 ;
 RECT 2.42 0.88 2.55 1.01 ;
 LAYER M1 ;
 RECT 0.78 1.91 4.9 2.05 ;
 END
END NOR2X4

MACRO NOR3X0
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.88 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.04 1.625 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN2

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.815 0.275 1.975 0.505 ;
 RECT 0.86 0.26 1 0.685 ;
 RECT 1.82 1.32 2.205 1.54 ;
 RECT 0.865 1.68 1.005 2.65 ;
 RECT 0.725 1.56 1.96 1.68 ;
 RECT 0.725 1.54 2.205 1.56 ;
 RECT 1.82 0.825 1.96 1.32 ;
 RECT 0.86 0.685 1.96 0.825 ;
 RECT 1.82 0.505 1.96 0.685 ;
 END
 ANTENNADIFFAREA 0.605 ;
 END QN

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.88 0.08 ;
 RECT 1.34 0.08 1.48 0.505 ;
 RECT 0.31 0.08 0.45 0.755 ;
 RECT 2.3 0.08 2.44 0.555 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.88 2.96 ;
 RECT 2.39 1.52 2.53 2.8 ;
 RECT 0.355 1.495 0.495 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.11 1.125 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.125 0.745 2.535 1.045 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN3

 OBS
 LAYER PO ;
 RECT 1.4 1.14 1.705 1.37 ;
 RECT 1.605 0.105 1.705 1.14 ;
 RECT 1.605 1.37 1.705 2.755 ;
 RECT 0.9 1.14 1.22 1.37 ;
 RECT 1.12 0.105 1.22 1.14 ;
 RECT 1.12 1.37 1.22 2.76 ;
 RECT 2.085 0.105 2.185 0.745 ;
 RECT 2.085 0.975 2.185 2.765 ;
 RECT 2.085 0.745 2.315 0.975 ;
 LAYER CO ;
 RECT 0.87 2.36 1 2.49 ;
 RECT 0.87 2.09 1 2.22 ;
 RECT 0.87 1.815 1 1.945 ;
 RECT 2.395 1.675 2.525 1.805 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 2.395 2.225 2.525 2.355 ;
 RECT 0.95 1.19 1.08 1.32 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 1.345 0.325 1.475 0.455 ;
 RECT 1.83 0.325 1.96 0.455 ;
 RECT 0.87 1.545 1 1.675 ;
 RECT 0.865 0.325 0.995 0.455 ;
 RECT 2.135 0.795 2.265 0.925 ;
 RECT 1.45 1.19 1.58 1.32 ;
 RECT 2.305 0.325 2.435 0.455 ;
 END
END NOR3X0

MACRO NOR3X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.12 1.68 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 2.3 0.08 2.44 0.555 ;
 RECT 3.4 0.08 3.54 0.875 ;
 RECT 1.34 0.08 1.48 0.505 ;
 RECT 0.31 0.08 0.45 0.755 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 3.39 2.13 3.53 2.8 ;
 RECT 2.39 1.64 2.53 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.11 1.135 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.12 0.745 2.485 1.08 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN3

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.72 0.68 4.01 0.92 ;
 RECT 3.87 0.92 4.01 2.245 ;
 RECT 3.87 0.31 4.01 0.68 ;
 END
 ANTENNADIFFAREA 0.498 ;
 END QN

 OBS
 LAYER PO ;
 RECT 0.9 1.14 1.22 1.37 ;
 RECT 1.12 0.105 1.22 1.14 ;
 RECT 1.12 1.37 1.22 2.745 ;
 RECT 3.655 0.155 3.755 1.12 ;
 RECT 3.655 1.35 3.755 2.785 ;
 RECT 3.495 1.12 3.755 1.35 ;
 RECT 2.085 0.105 2.185 0.745 ;
 RECT 2.085 0.975 2.185 2.745 ;
 RECT 2.085 0.745 2.315 0.975 ;
 RECT 1.445 1.14 1.705 1.37 ;
 RECT 1.605 0.105 1.705 1.14 ;
 RECT 1.605 1.37 1.705 2.745 ;
 RECT 2.715 0.105 2.815 1.12 ;
 RECT 2.715 1.35 2.815 2.185 ;
 RECT 2.61 1.12 2.84 1.35 ;
 LAYER CO ;
 RECT 2.66 1.17 2.79 1.3 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 1.345 0.325 1.475 0.455 ;
 RECT 1.83 0.325 1.96 0.455 ;
 RECT 0.87 1.545 1 1.675 ;
 RECT 2.95 1.805 3.08 1.935 ;
 RECT 0.865 0.325 0.995 0.455 ;
 RECT 2.135 0.795 2.265 0.925 ;
 RECT 1.495 1.19 1.625 1.32 ;
 RECT 2.95 0.325 3.08 0.455 ;
 RECT 2.305 0.325 2.435 0.455 ;
 RECT 3.545 1.17 3.675 1.3 ;
 RECT 3.875 1.505 4.005 1.635 ;
 RECT 3.875 0.46 4.005 0.59 ;
 RECT 3.875 2.025 4.005 2.155 ;
 RECT 3.875 1.765 4.005 1.895 ;
 RECT 3.405 0.68 3.535 0.81 ;
 RECT 3.405 0.405 3.535 0.535 ;
 RECT 3.395 2.185 3.525 2.315 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 2.395 1.735 2.525 1.865 ;
 RECT 2.95 1.545 3.08 1.675 ;
 RECT 0.95 1.19 1.08 1.32 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 0.315 0.575 0.445 0.705 ;
 LAYER M1 ;
 RECT 0.86 0.26 1 0.685 ;
 RECT 1.82 0.825 1.96 1.255 ;
 RECT 1.82 0.505 1.96 0.685 ;
 RECT 0.86 0.685 1.96 0.825 ;
 RECT 1.82 1.395 1.96 1.54 ;
 RECT 0.725 1.54 1.96 1.68 ;
 RECT 1.815 0.275 1.975 0.505 ;
 RECT 2.645 1.12 2.8 1.255 ;
 RECT 1.82 1.255 2.8 1.395 ;
 RECT 2.945 0.275 3.085 1.185 ;
 RECT 2.945 1.325 3.085 2.03 ;
 RECT 3.53 1.12 3.685 1.185 ;
 RECT 3.53 1.325 3.685 1.35 ;
 RECT 2.945 1.185 3.685 1.325 ;
 END
END NOR3X1

MACRO LSDNSSX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 RECT 1.97 0.08 2.11 0.765 ;
 RECT 0.62 0.08 0.76 0.53 ;
 RECT 1.565 0.08 1.705 0.59 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.36 0.8 0.66 1.155 ;
 END
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 RECT 0.615 1.66 0.755 2.8 ;
 RECT 1.56 1.725 1.7 2.8 ;
 RECT 1.97 1.935 2.11 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.965 1.705 1.285 2.08 ;
 RECT 1.09 0.505 1.23 1.705 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 1.345 0.1 1.445 1.175 ;
 RECT 1.345 1.275 1.445 2.785 ;
 RECT 0.755 1.175 1.445 1.275 ;
 RECT 0.755 1.275 0.985 1.405 ;
 RECT 0.875 0.1 0.975 1.175 ;
 RECT 0.875 1.405 0.975 2.785 ;
 RECT 0.4 0.1 0.5 0.92 ;
 RECT 0.4 1.15 0.5 2.235 ;
 RECT 0.33 0.92 0.56 1.15 ;
 LAYER CO ;
 RECT 0.145 1.815 0.275 1.945 ;
 RECT 0.805 1.225 0.935 1.355 ;
 RECT 1.975 2.265 2.105 2.395 ;
 RECT 1.975 2.005 2.105 2.135 ;
 RECT 1.565 1.795 1.695 1.925 ;
 RECT 1.565 2.31 1.695 2.44 ;
 RECT 1.095 0.57 1.225 0.7 ;
 RECT 0.62 2.31 0.75 2.44 ;
 RECT 1.095 1.915 1.225 2.045 ;
 RECT 1.57 0.39 1.7 0.52 ;
 RECT 1.095 1.615 1.225 1.745 ;
 RECT 0.625 0.33 0.755 0.46 ;
 RECT 0.62 1.735 0.75 1.865 ;
 RECT 0.38 0.97 0.51 1.1 ;
 RECT 0.145 1.545 0.275 1.675 ;
 RECT 0.15 0.33 0.28 0.46 ;
 RECT 1.975 0.305 2.105 0.435 ;
 RECT 1.975 0.565 2.105 0.695 ;
 LAYER M1 ;
 RECT 0.145 0.26 0.285 0.52 ;
 RECT 0.08 0.52 0.285 0.66 ;
 RECT 0.08 0.66 0.22 1.295 ;
 RECT 0.08 1.295 0.28 1.435 ;
 RECT 0.14 1.435 0.28 2.015 ;
 RECT 0.8 1.105 0.94 1.425 ;
 RECT 0.145 1.295 0.94 1.435 ;
 END
END LSDNSSX2

MACRO LSDNSSX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 0.615 0.08 0.755 0.54 ;
 RECT 1.56 0.08 1.7 0.59 ;
 RECT 2.515 0.08 2.655 0.59 ;
 RECT 2.925 0.08 3.065 0.89 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.36 0.84 0.66 1.14 ;
 END
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 0.615 1.625 0.755 2.8 ;
 RECT 1.56 1.725 1.7 2.8 ;
 RECT 2.925 1.935 3.065 2.8 ;
 RECT 2.51 1.725 2.65 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.965 1.705 1.285 2.08 ;
 RECT 1.09 1.27 2.18 1.41 ;
 RECT 1.09 1.41 1.23 1.705 ;
 RECT 1.09 0.505 1.23 1.27 ;
 RECT 2.04 1.41 2.18 2.13 ;
 RECT 2.04 0.505 2.18 1.27 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 0.87 0.89 1.445 0.96 ;
 RECT 0.87 0.96 2.395 0.99 ;
 RECT 1.345 0.99 2.395 1.06 ;
 RECT 1.345 1.06 1.445 2.785 ;
 RECT 0.87 0.1 0.97 0.89 ;
 RECT 0.87 0.99 0.97 1.17 ;
 RECT 1.815 0.1 1.915 0.96 ;
 RECT 1.815 1.06 1.915 2.785 ;
 RECT 2.295 0.1 2.395 0.96 ;
 RECT 2.295 1.06 2.395 2.785 ;
 RECT 1.345 0.1 1.445 0.89 ;
 RECT 0.87 1.4 0.97 2.785 ;
 RECT 0.755 1.17 0.985 1.4 ;
 RECT 0.4 0.1 0.5 0.91 ;
 RECT 0.4 1.14 0.5 2.335 ;
 RECT 0.345 0.91 0.575 1.14 ;
 LAYER CO ;
 RECT 2.93 0.43 3.06 0.56 ;
 RECT 2.93 0.69 3.06 0.82 ;
 RECT 2.045 1.915 2.175 2.045 ;
 RECT 2.515 1.795 2.645 1.925 ;
 RECT 2.52 0.39 2.65 0.52 ;
 RECT 2.045 1.615 2.175 1.745 ;
 RECT 2.515 2.31 2.645 2.44 ;
 RECT 2.045 0.57 2.175 0.7 ;
 RECT 0.805 1.22 0.935 1.35 ;
 RECT 2.93 2.265 3.06 2.395 ;
 RECT 2.93 2.005 3.06 2.135 ;
 RECT 1.565 1.795 1.695 1.925 ;
 RECT 1.565 2.31 1.695 2.44 ;
 RECT 1.095 0.57 1.225 0.7 ;
 RECT 0.62 2.31 0.75 2.44 ;
 RECT 1.095 1.915 1.225 2.045 ;
 RECT 1.565 0.39 1.695 0.52 ;
 RECT 1.095 1.615 1.225 1.745 ;
 RECT 0.62 0.34 0.75 0.47 ;
 RECT 0.62 1.735 0.75 1.865 ;
 RECT 0.395 0.96 0.525 1.09 ;
 RECT 0.15 1.545 0.28 1.675 ;
 RECT 0.15 0.33 0.28 0.46 ;
 LAYER M1 ;
 RECT 0.145 0.26 0.285 0.52 ;
 RECT 0.08 0.52 0.285 0.66 ;
 RECT 0.08 0.66 0.22 1.295 ;
 RECT 0.08 1.295 0.285 1.435 ;
 RECT 0.145 1.435 0.285 1.74 ;
 RECT 0.8 1.15 0.94 1.425 ;
 RECT 0.145 1.285 0.94 1.425 ;
 END
END LSDNSSX4

MACRO NOR4X0
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 0.625 0.08 0.765 0.505 ;
 RECT 1.575 0.08 1.735 0.505 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 2.65 0.08 2.79 0.505 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.16 1.14 1.455 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.52 1.14 0.905 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.89 1.065 2.2 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN3

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 2.645 1.88 2.785 2.8 ;
 END
 END VDD

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.355 1.12 2.68 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN4

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.105 0.275 1.245 0.645 ;
 RECT 0.555 1.54 1.735 1.68 ;
 RECT 1.105 0.645 2.36 0.785 ;
 RECT 2.065 0.52 2.36 0.645 ;
 RECT 2.065 0.27 2.205 0.52 ;
 RECT 1.595 0.785 1.735 1.54 ;
 RECT 0.595 1.68 0.745 2.545 ;
 END
 ANTENNADIFFAREA 0.526 ;
 END QN

 OBS
 LAYER PO ;
 RECT 0.72 1.14 0.98 1.37 ;
 RECT 0.88 0.105 0.98 1.14 ;
 RECT 0.88 1.37 0.98 2.755 ;
 RECT 1.205 1.14 1.465 1.37 ;
 RECT 1.365 0.105 1.465 1.14 ;
 RECT 1.365 1.37 1.465 2.745 ;
 RECT 1.85 0.105 1.95 1.065 ;
 RECT 1.85 1.295 1.95 2.75 ;
 RECT 1.85 1.065 2.08 1.295 ;
 RECT 2.345 0.105 2.445 1.12 ;
 RECT 2.345 1.35 2.445 2.755 ;
 RECT 2.345 1.12 2.575 1.35 ;
 LAYER CO ;
 RECT 2.65 1.95 2.78 2.08 ;
 RECT 1.11 0.325 1.24 0.455 ;
 RECT 0.605 1.815 0.735 1.945 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 2.07 0.325 2.2 0.455 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 0.605 2.345 0.735 2.475 ;
 RECT 0.605 1.545 0.735 1.675 ;
 RECT 0.77 1.19 0.9 1.32 ;
 RECT 1.9 1.115 2.03 1.245 ;
 RECT 1.255 1.19 1.385 1.32 ;
 RECT 1.59 0.325 1.72 0.455 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 2.395 1.17 2.525 1.3 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 2.655 0.325 2.785 0.455 ;
 RECT 0.63 0.325 0.76 0.455 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 2.65 2.225 2.78 2.355 ;
 RECT 0.605 2.085 0.735 2.215 ;
 END
END NOR4X0

MACRO NOR4X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 0.68 1.095 1.07 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.535 0.745 1.88 1.08 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.8 0.745 5.165 1.08 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END IN3

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.04 0.84 4.36 1.08 ;
 END
 ANTENNAGATEAREA 0.096 ;
 END IN4

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 1.71 0.08 1.85 0.555 ;
 RECT 0.31 0.08 0.45 0.755 ;
 RECT 4.975 0.08 5.115 0.555 ;
 RECT 3.05 0.08 3.19 0.59 ;
 RECT 0.77 0.08 0.91 0.505 ;
 RECT 4.035 0.08 4.175 0.505 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 3.135 2.355 3.275 2.8 ;
 RECT 1.71 1.935 1.85 2.8 ;
 RECT 4.975 1.495 5.115 2.8 ;
 RECT 2.11 1.6 2.25 2.8 ;
 END
 END VDD

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.56 0.68 3.8 0.92 ;
 RECT 3.635 0.92 3.775 1.795 ;
 RECT 3.635 0.31 3.775 0.68 ;
 END
 ANTENNADIFFAREA 0.479 ;
 END QN

 OBS
 LAYER PO ;
 RECT 2.835 0.14 2.935 2.07 ;
 RECT 2.685 2.07 2.935 2.3 ;
 RECT 3.21 1.155 3.515 1.385 ;
 RECT 3.415 0.14 3.515 1.155 ;
 RECT 3.415 1.385 3.515 2.785 ;
 RECT 2.365 0.14 2.465 0.88 ;
 RECT 2.365 1.11 2.465 2.01 ;
 RECT 2.235 0.88 2.465 1.11 ;
 RECT 4.29 1.07 4.39 2.38 ;
 RECT 4.29 0.105 4.39 0.84 ;
 RECT 4.13 0.84 4.39 1.07 ;
 RECT 4.76 0.975 4.86 2.38 ;
 RECT 4.76 0.105 4.86 0.745 ;
 RECT 4.76 0.745 4.99 0.975 ;
 RECT 1.025 0.105 1.125 0.84 ;
 RECT 0.865 0.84 1.125 1.07 ;
 RECT 1.025 1.07 1.125 2.375 ;
 RECT 1.495 0.105 1.595 0.745 ;
 RECT 1.495 0.975 1.595 2.38 ;
 RECT 1.495 0.745 1.725 0.975 ;
 LAYER CO ;
 RECT 0.915 0.89 1.045 1.02 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 1.715 0.325 1.845 0.455 ;
 RECT 1.545 0.795 1.675 0.925 ;
 RECT 1.715 2.01 1.845 2.14 ;
 RECT 2.735 2.12 2.865 2.25 ;
 RECT 3.14 2.405 3.27 2.535 ;
 RECT 2.275 0.93 2.405 1.06 ;
 RECT 2.115 1.65 2.245 1.78 ;
 RECT 2.585 1.58 2.715 1.71 ;
 RECT 3.055 0.36 3.185 0.49 ;
 RECT 3.26 1.205 3.39 1.335 ;
 RECT 2.115 0.36 2.245 0.49 ;
 RECT 3.64 0.36 3.77 0.49 ;
 RECT 3.64 1.58 3.77 1.71 ;
 RECT 4.98 1.545 5.11 1.675 ;
 RECT 4.04 1.545 4.17 1.675 ;
 RECT 4.04 0.325 4.17 0.455 ;
 RECT 4.51 0.325 4.64 0.455 ;
 RECT 4.18 0.89 4.31 1.02 ;
 RECT 4.81 0.795 4.94 0.925 ;
 RECT 4.98 1.545 5.11 1.675 ;
 RECT 4.98 0.325 5.11 0.455 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 0.775 1.545 0.905 1.675 ;
 RECT 1.245 0.325 1.375 0.455 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 0.775 0.325 0.905 0.455 ;
 LAYER M1 ;
 RECT 2.58 0.495 2.72 1.245 ;
 RECT 2.58 1.385 2.72 1.78 ;
 RECT 2.065 0.355 2.72 0.495 ;
 RECT 3.21 1.155 3.44 1.245 ;
 RECT 2.58 1.245 3.44 1.385 ;
 RECT 2.73 2.185 2.87 2.3 ;
 RECT 4.5 0.505 4.64 1.48 ;
 RECT 4.035 1.62 4.175 2.045 ;
 RECT 2.695 2.045 4.175 2.185 ;
 RECT 4.495 0.275 4.655 0.505 ;
 RECT 4.035 1.48 4.645 1.62 ;
 RECT 1.235 0.505 1.375 1.32 ;
 RECT 0.77 1.46 0.91 1.835 ;
 RECT 1.23 0.275 1.39 0.505 ;
 RECT 0.77 1.32 2.41 1.46 ;
 RECT 2.27 0.88 2.41 1.32 ;
 END
END NOR4X1

MACRO OR2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 2.56 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 2.56 2.96 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 1.71 1.66 1.85 2.8 ;
 END
 END VDD

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.33 2.325 1.57 2.66 ;
 END
 ANTENNAGATEAREA 0.111 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.66 0.83 1.095 1.08 ;
 END
 ANTENNAGATEAREA 0.111 ;
 END IN1

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 2.56 0.08 ;
 RECT 0.77 0.08 0.91 0.505 ;
 RECT 1.71 0.08 1.85 0.505 ;
 RECT 0.31 0.08 0.45 0.755 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.63 0.78 2.44 0.92 ;
 RECT 1.63 0.68 1.88 0.78 ;
 RECT 2.3 0.92 2.44 2.585 ;
 RECT 2.3 0.22 2.44 0.78 ;
 END
 ANTENNADIFFAREA 0.496 ;
 END Q

 OBS
 LAYER PO ;
 RECT 2.075 0.105 2.175 1.14 ;
 RECT 2.075 1.37 2.175 2.77 ;
 RECT 1.97 1.14 2.2 1.37 ;
 RECT 1.025 0.105 1.125 0.84 ;
 RECT 0.865 0.84 1.125 1.07 ;
 RECT 1.025 1.07 1.125 2.635 ;
 RECT 1.495 0.105 1.595 2.425 ;
 RECT 1.37 2.425 1.6 2.655 ;
 LAYER CO ;
 RECT 2.305 0.325 2.435 0.455 ;
 RECT 2.305 0.585 2.435 0.715 ;
 RECT 2.305 2.345 2.435 2.475 ;
 RECT 1.715 2.08 1.845 2.21 ;
 RECT 1.715 1.805 1.845 1.935 ;
 RECT 0.775 2.09 0.905 2.22 ;
 RECT 0.775 1.81 0.905 1.94 ;
 RECT 1.245 0.325 1.375 0.455 ;
 RECT 1.715 0.325 1.845 0.455 ;
 RECT 1.42 2.475 1.55 2.605 ;
 RECT 0.915 0.89 1.045 1.02 ;
 RECT 2.305 1.545 2.435 1.675 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 0.775 0.325 0.905 0.455 ;
 RECT 2.305 1.805 2.435 1.935 ;
 RECT 2.305 2.065 2.435 2.195 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 2.02 1.19 2.15 1.32 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 0.775 1.545 0.905 1.675 ;
 LAYER M1 ;
 RECT 0.77 1.26 0.91 2.38 ;
 RECT 1.23 0.275 1.39 0.505 ;
 RECT 1.235 0.44 1.375 1.34 ;
 RECT 2.005 1.14 2.16 1.37 ;
 RECT 0.87 1.26 2.12 1.4 ;
 END
END OR2X1

MACRO OR2X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 0.77 0.08 0.91 0.505 ;
 RECT 2.78 0.08 2.92 0.555 ;
 RECT 1.71 0.08 1.85 0.555 ;
 RECT 0.31 0.08 0.45 0.755 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.535 0.745 1.88 1.085 ;
 END
 ANTENNAGATEAREA 0.116 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.665 0.83 1.095 1.08 ;
 END
 ANTENNAGATEAREA 0.116 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 1.71 1.66 1.85 2.8 ;
 RECT 2.785 1.495 2.925 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.3 0.805 2.545 1.065 ;
 RECT 2.3 1.065 2.44 2.585 ;
 RECT 2.3 0.275 2.44 0.805 ;
 END
 ANTENNADIFFAREA 0.616 ;
 END Q

 OBS
 LAYER PO ;
 RECT 1.025 1.07 1.125 2.585 ;
 RECT 1.025 0.105 1.125 0.84 ;
 RECT 0.865 0.84 1.125 1.07 ;
 RECT 2.56 0.105 2.66 1.18 ;
 RECT 2.56 1.28 2.66 2.74 ;
 RECT 2.075 0.105 2.175 1.14 ;
 RECT 1.97 1.14 2.2 1.18 ;
 RECT 1.97 1.28 2.2 1.37 ;
 RECT 1.97 1.18 2.66 1.28 ;
 RECT 2.075 1.37 2.175 2.755 ;
 RECT 1.495 0.105 1.595 0.745 ;
 RECT 1.495 0.975 1.595 2.585 ;
 RECT 1.495 0.745 1.725 0.975 ;
 LAYER CO ;
 RECT 0.915 0.89 1.045 1.02 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 2.79 1.545 2.92 1.675 ;
 RECT 2.79 1.545 2.92 1.675 ;
 RECT 0.775 1.81 0.905 1.94 ;
 RECT 2.305 2.065 2.435 2.195 ;
 RECT 2.79 2.08 2.92 2.21 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 2.025 1.19 2.155 1.32 ;
 RECT 2.305 0.325 2.435 0.455 ;
 RECT 0.775 2.09 0.905 2.22 ;
 RECT 1.715 0.325 1.845 0.455 ;
 RECT 2.785 0.325 2.915 0.455 ;
 RECT 1.715 2.08 1.845 2.21 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 0.775 0.325 0.905 0.455 ;
 RECT 2.79 1.805 2.92 1.935 ;
 RECT 2.305 1.805 2.435 1.935 ;
 RECT 2.305 1.545 2.435 1.675 ;
 RECT 0.775 1.545 0.905 1.675 ;
 RECT 1.715 1.805 1.845 1.935 ;
 RECT 2.305 2.345 2.435 2.475 ;
 RECT 1.245 0.325 1.375 0.455 ;
 RECT 1.545 0.795 1.675 0.925 ;
 LAYER M1 ;
 RECT 1.23 0.275 1.39 0.505 ;
 RECT 1.235 0.44 1.375 1.34 ;
 RECT 0.77 1.28 0.91 2.38 ;
 RECT 2.02 1.14 2.16 1.425 ;
 RECT 0.87 1.28 2.12 1.42 ;
 END
END OR2X2

MACRO OR2X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 0.31 0.08 0.45 0.755 ;
 RECT 2.78 0.08 2.92 0.555 ;
 RECT 1.71 0.08 1.85 0.555 ;
 RECT 3.74 0.08 3.88 0.555 ;
 RECT 0.77 0.08 0.91 0.505 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.535 0.745 1.88 1.09 ;
 END
 ANTENNAGATEAREA 0.111 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.3 0.275 2.44 0.68 ;
 RECT 2.28 0.68 2.52 0.935 ;
 RECT 2.28 0.935 3.405 0.98 ;
 RECT 2.3 0.98 3.405 1.075 ;
 RECT 2.3 1.075 2.44 2.585 ;
 RECT 3.265 0.275 3.405 0.935 ;
 RECT 3.265 1.075 3.405 2.585 ;
 END
 ANTENNADIFFAREA 1.24 ;
 END Q

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.665 0.83 1.095 1.08 ;
 END
 ANTENNAGATEAREA 0.111 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 1.71 1.66 1.85 2.8 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 2.785 1.495 2.925 2.8 ;
 RECT 3.74 1.495 3.88 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 1.495 0.975 1.595 2.535 ;
 RECT 1.495 0.105 1.595 0.745 ;
 RECT 1.495 0.745 1.725 0.975 ;
 RECT 2.075 0.105 2.175 1.12 ;
 RECT 3.525 0.105 3.625 1.18 ;
 RECT 1.97 1.18 3.625 1.28 ;
 RECT 3.525 1.28 3.625 2.77 ;
 RECT 3.045 0.105 3.145 1.18 ;
 RECT 3.045 1.28 3.145 2.745 ;
 RECT 2.075 1.35 2.175 2.755 ;
 RECT 2.56 0.105 2.66 1.18 ;
 RECT 1.97 1.12 2.2 1.18 ;
 RECT 1.97 1.28 2.2 1.35 ;
 RECT 2.56 1.28 2.66 2.74 ;
 RECT 1.025 0.105 1.125 0.84 ;
 RECT 0.865 0.84 1.125 1.07 ;
 RECT 1.025 1.07 1.125 2.53 ;
 LAYER CO ;
 RECT 3.745 0.325 3.875 0.455 ;
 RECT 3.745 1.545 3.875 1.675 ;
 RECT 3.745 2.08 3.875 2.21 ;
 RECT 3.745 1.805 3.875 1.935 ;
 RECT 3.745 1.545 3.875 1.675 ;
 RECT 3.27 0.6 3.4 0.73 ;
 RECT 3.27 1.545 3.4 1.675 ;
 RECT 3.27 2.345 3.4 2.475 ;
 RECT 3.27 2.065 3.4 2.195 ;
 RECT 3.27 0.325 3.4 0.455 ;
 RECT 3.27 1.805 3.4 1.935 ;
 RECT 1.545 0.795 1.675 0.925 ;
 RECT 2.025 1.17 2.155 1.3 ;
 RECT 2.79 2.08 2.92 2.21 ;
 RECT 2.305 2.345 2.435 2.475 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 1.715 0.325 1.845 0.455 ;
 RECT 0.775 0.325 0.905 0.455 ;
 RECT 0.915 0.89 1.045 1.02 ;
 RECT 2.305 0.325 2.435 0.455 ;
 RECT 0.775 1.545 0.905 1.675 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 0.775 1.81 0.905 1.94 ;
 RECT 2.305 0.6 2.435 0.73 ;
 RECT 1.715 1.805 1.845 1.935 ;
 RECT 1.245 0.325 1.375 0.455 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 1.715 2.08 1.845 2.21 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 2.305 2.065 2.435 2.195 ;
 RECT 2.79 1.805 2.92 1.935 ;
 RECT 2.305 1.805 2.435 1.935 ;
 RECT 2.79 1.545 2.92 1.675 ;
 RECT 2.305 1.545 2.435 1.675 ;
 RECT 0.775 2.09 0.905 2.22 ;
 RECT 2.785 0.325 2.915 0.455 ;
 RECT 2.79 1.545 2.92 1.675 ;
 LAYER M1 ;
 RECT 1.23 0.275 1.39 0.505 ;
 RECT 1.235 0.44 1.375 1.34 ;
 RECT 0.77 1.265 0.91 2.38 ;
 RECT 2.02 1.12 2.16 1.35 ;
 RECT 0.87 1.265 2.16 1.405 ;
 END
END OR2X4

MACRO OR3X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.12 1.68 1.4 ;
 END
 ANTENNAGATEAREA 0.131 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 1.34 0.08 1.48 0.505 ;
 RECT 2.3 0.08 2.44 0.555 ;
 RECT 0.31 0.08 0.45 0.755 ;
 END
 END VSS

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.12 0.745 2.4 1.1 ;
 END
 ANTENNAGATEAREA 0.131 ;
 END IN3

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 2.39 1.8 2.53 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.76 0.66 3.085 0.93 ;
 RECT 2.945 0.93 3.085 2.245 ;
 RECT 2.945 0.275 3.085 0.66 ;
 END
 ANTENNADIFFAREA 0.529 ;
 END Q

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.805 1.12 1.16 1.4 ;
 END
 ANTENNAGATEAREA 0.131 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 0.935 1.14 1.22 1.37 ;
 RECT 1.12 0.105 1.22 1.14 ;
 RECT 1.12 1.37 1.22 2.73 ;
 RECT 2.715 0.105 2.815 1.13 ;
 RECT 2.715 1.36 2.815 2.76 ;
 RECT 2.61 1.13 2.84 1.36 ;
 RECT 1.445 1.14 1.705 1.37 ;
 RECT 1.605 0.105 1.705 1.14 ;
 RECT 1.605 1.37 1.705 2.73 ;
 RECT 2.085 0.105 2.185 0.745 ;
 RECT 2.085 0.975 2.185 2.72 ;
 RECT 2.085 0.745 2.315 0.975 ;
 LAYER CO ;
 RECT 2.95 0.605 3.08 0.735 ;
 RECT 2.395 1.965 2.525 2.095 ;
 RECT 0.985 1.19 1.115 1.32 ;
 RECT 0.865 0.325 0.995 0.455 ;
 RECT 2.95 2.065 3.08 2.195 ;
 RECT 2.95 1.545 3.08 1.675 ;
 RECT 2.95 1.805 3.08 1.935 ;
 RECT 2.95 0.325 3.08 0.455 ;
 RECT 1.495 1.19 1.625 1.32 ;
 RECT 2.135 0.795 2.265 0.925 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 0.87 1.545 1 1.675 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 2.395 2.225 2.525 2.355 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 2.66 1.18 2.79 1.31 ;
 RECT 2.305 0.325 2.435 0.455 ;
 RECT 1.83 0.325 1.96 0.455 ;
 RECT 1.345 0.325 1.475 0.455 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 0.36 1.805 0.49 1.935 ;
 LAYER M1 ;
 RECT 0.86 0.22 1 0.645 ;
 RECT 0.86 0.645 1.895 0.785 ;
 RECT 1.815 0.275 1.975 0.505 ;
 RECT 1.82 0.44 1.96 1.34 ;
 RECT 1.82 1.16 1.96 1.54 ;
 RECT 0.725 1.54 1.96 1.68 ;
 RECT 1.875 1.5 2.8 1.64 ;
 RECT 2.66 1.245 2.8 1.5 ;
 RECT 2.645 1.13 2.8 1.36 ;
 END
END OR3X1

MACRO OR3X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 1.34 0.08 1.48 0.505 ;
 RECT 0.31 0.08 0.45 0.755 ;
 RECT 2.3 0.08 2.44 0.555 ;
 RECT 3.445 0.08 3.585 0.555 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 2.39 1.55 2.53 2.8 ;
 RECT 3.445 1.485 3.585 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.805 1.12 1.18 1.4 ;
 END
 ANTENNAGATEAREA 0.131 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.1 0.745 2.37 1.08 ;
 END
 ANTENNAGATEAREA 0.131 ;
 END IN3

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.125 1.68 1.4 ;
 END
 ANTENNAGATEAREA 0.131 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.945 1.09 3.085 2.245 ;
 RECT 2.945 0.835 3.32 1.09 ;
 RECT 2.945 0.275 3.085 0.835 ;
 END
 ANTENNADIFFAREA 0.68 ;
 END Q

 OBS
 LAYER PO ;
 RECT 0.955 1.14 1.22 1.37 ;
 RECT 1.12 0.105 1.22 1.14 ;
 RECT 1.12 1.37 1.22 2.73 ;
 RECT 2.715 0.105 2.815 1.14 ;
 RECT 3.22 0.105 3.32 1.165 ;
 RECT 2.61 1.165 3.32 1.265 ;
 RECT 3.22 1.265 3.32 2.76 ;
 RECT 2.61 1.14 2.84 1.165 ;
 RECT 2.61 1.265 2.84 1.37 ;
 RECT 2.715 1.37 2.815 2.76 ;
 RECT 1.445 1.14 1.705 1.37 ;
 RECT 1.605 0.105 1.705 1.14 ;
 RECT 1.605 1.37 1.705 2.73 ;
 RECT 2.085 0.105 2.185 0.745 ;
 RECT 2.085 0.975 2.185 2.72 ;
 RECT 2.085 0.745 2.315 0.975 ;
 LAYER CO ;
 RECT 2.395 1.68 2.525 1.81 ;
 RECT 2.395 1.94 2.525 2.07 ;
 RECT 3.45 1.665 3.58 1.795 ;
 RECT 3.45 1.95 3.58 2.08 ;
 RECT 3.45 0.325 3.58 0.455 ;
 RECT 3.45 2.225 3.58 2.355 ;
 RECT 2.95 0.325 3.08 0.455 ;
 RECT 2.305 0.325 2.435 0.455 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 2.95 1.545 3.08 1.675 ;
 RECT 2.95 2.065 3.08 2.195 ;
 RECT 1.005 1.19 1.135 1.32 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 2.135 0.795 2.265 0.925 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 1.495 1.19 1.625 1.32 ;
 RECT 2.66 1.19 2.79 1.32 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 2.395 2.225 2.525 2.355 ;
 RECT 0.865 0.325 0.995 0.455 ;
 RECT 1.345 0.325 1.475 0.455 ;
 RECT 1.83 0.325 1.96 0.455 ;
 RECT 0.87 1.545 1 1.675 ;
 RECT 2.95 1.805 3.08 1.935 ;
 LAYER M1 ;
 RECT 0.86 0.26 1 0.685 ;
 RECT 0.725 1.54 1.96 1.68 ;
 RECT 1.82 1.16 1.96 1.54 ;
 RECT 0.86 0.685 1.895 0.825 ;
 RECT 1.82 0.44 1.96 1.34 ;
 RECT 1.815 0.275 1.975 0.505 ;
 RECT 2.66 1.18 2.8 1.255 ;
 RECT 2.645 1.14 2.8 1.37 ;
 RECT 1.875 1.255 2.8 1.395 ;
 END
END OR3X2

MACRO OR3X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 2.88 ;
 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.32 1.04 1.68 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.925 0.275 4.065 0.83 ;
 RECT 3.88 0.83 4.12 1.04 ;
 RECT 2.945 1.185 3.085 2.245 ;
 RECT 3.925 1.18 4.065 2.245 ;
 RECT 2.945 0.275 3.085 1.04 ;
 RECT 2.945 1.18 3.28 1.185 ;
 RECT 2.945 1.09 4.065 1.18 ;
 RECT 2.945 1.04 4.12 1.09 ;
 END
 ANTENNADIFFAREA 1.392 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 0.355 1.495 0.495 2.8 ;
 RECT 3.445 1.59 3.585 2.8 ;
 RECT 2.39 1.595 2.53 2.8 ;
 RECT 4.41 1.57 4.55 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.815 1.04 1.18 1.4 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.1 0.745 2.385 1.08 ;
 END
 ANTENNAGATEAREA 0.133 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 1.34 0.08 1.48 0.505 ;
 RECT 2.3 0.08 2.44 0.555 ;
 RECT 0.31 0.08 0.45 0.755 ;
 RECT 3.445 0.08 3.585 0.555 ;
 RECT 4.405 0.08 4.545 0.555 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 2.715 0.105 2.815 1.12 ;
 RECT 4.19 0.105 4.29 1.165 ;
 RECT 2.61 1.165 4.29 1.265 ;
 RECT 4.19 1.265 4.29 2.76 ;
 RECT 3.705 0.105 3.805 1.165 ;
 RECT 3.705 1.265 3.805 2.76 ;
 RECT 3.22 0.105 3.32 1.165 ;
 RECT 3.22 1.265 3.32 2.76 ;
 RECT 2.715 1.35 2.815 2.76 ;
 RECT 2.61 1.12 2.84 1.165 ;
 RECT 2.61 1.265 2.84 1.35 ;
 RECT 1.445 1.14 1.705 1.37 ;
 RECT 1.605 0.105 1.705 1.14 ;
 RECT 1.605 1.37 1.705 2.745 ;
 RECT 0.955 1.14 1.22 1.37 ;
 RECT 1.12 0.105 1.22 1.14 ;
 RECT 1.12 1.37 1.22 2.75 ;
 RECT 2.085 0.975 2.185 2.75 ;
 RECT 2.085 0.105 2.185 0.745 ;
 RECT 2.085 0.745 2.315 0.975 ;
 LAYER CO ;
 RECT 4.415 1.655 4.545 1.785 ;
 RECT 4.415 1.95 4.545 2.08 ;
 RECT 3.45 1.695 3.58 1.825 ;
 RECT 3.45 1.965 3.58 2.095 ;
 RECT 2.395 1.695 2.525 1.825 ;
 RECT 2.395 1.955 2.525 2.085 ;
 RECT 4.41 0.325 4.54 0.455 ;
 RECT 4.415 2.225 4.545 2.355 ;
 RECT 3.93 1.805 4.06 1.935 ;
 RECT 3.93 1.545 4.06 1.675 ;
 RECT 3.93 2.065 4.06 2.195 ;
 RECT 3.93 0.325 4.06 0.455 ;
 RECT 0.36 1.545 0.49 1.675 ;
 RECT 2.95 2.065 3.08 2.195 ;
 RECT 2.66 1.17 2.79 1.3 ;
 RECT 0.87 1.545 1 1.675 ;
 RECT 2.135 0.795 2.265 0.925 ;
 RECT 1.345 0.325 1.475 0.455 ;
 RECT 0.36 2.065 0.49 2.195 ;
 RECT 2.95 0.325 3.08 0.455 ;
 RECT 2.95 1.805 3.08 1.935 ;
 RECT 2.395 2.225 2.525 2.355 ;
 RECT 2.305 0.325 2.435 0.455 ;
 RECT 3.45 2.225 3.58 2.355 ;
 RECT 0.36 1.805 0.49 1.935 ;
 RECT 1.005 1.19 1.135 1.32 ;
 RECT 3.45 0.325 3.58 0.455 ;
 RECT 1.83 0.325 1.96 0.455 ;
 RECT 0.315 0.315 0.445 0.445 ;
 RECT 2.95 1.545 3.08 1.675 ;
 RECT 1.495 1.19 1.625 1.32 ;
 RECT 0.315 0.575 0.445 0.705 ;
 RECT 0.865 0.325 0.995 0.455 ;
 LAYER M1 ;
 RECT 0.86 0.26 1 0.685 ;
 RECT 0.725 1.54 1.96 1.68 ;
 RECT 0.86 0.685 1.895 0.825 ;
 RECT 1.82 1.16 1.96 1.54 ;
 RECT 1.82 0.44 1.96 1.34 ;
 RECT 1.815 0.275 1.975 0.505 ;
 RECT 2.66 1.18 2.8 1.255 ;
 RECT 2.645 1.12 2.8 1.35 ;
 RECT 1.875 1.255 2.8 1.395 ;
 END
END OR3X4

MACRO OR4X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.52 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.52 0.08 ;
 RECT 1.52 0.32 1.79 0.46 ;
 RECT 0.625 0.08 0.765 0.505 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 2.65 0.08 2.79 0.525 ;
 RECT 1.575 0.08 1.735 0.32 ;
 END
 END VSS

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.345 0.81 2.68 1.08 ;
 END
 ANTENNAGATEAREA 0.13 ;
 END IN4

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.1 1.07 1.405 1.4 ;
 END
 ANTENNAGATEAREA 0.13 ;
 END IN2

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.52 2.96 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 2.645 2.17 2.785 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.16 1.095 3.415 1.36 ;
 RECT 3.16 1.36 3.3 2.56 ;
 RECT 3.16 0.275 3.3 1.095 ;
 END
 ANTENNADIFFAREA 0.581 ;
 END Q

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.515 1.14 0.86 1.4 ;
 END
 ANTENNAGATEAREA 0.13 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.875 1.065 2.2 1.4 ;
 END
 ANTENNAGATEAREA 0.13 ;
 END IN3

 OBS
 LAYER PO ;
 RECT 1.205 1.14 1.465 1.37 ;
 RECT 1.365 0.09 1.465 1.14 ;
 RECT 1.365 1.37 1.465 2.79 ;
 RECT 0.675 1.14 0.98 1.37 ;
 RECT 0.88 0.09 0.98 1.14 ;
 RECT 0.88 1.37 0.98 2.79 ;
 RECT 2.915 0.09 3.015 1.14 ;
 RECT 2.915 1.37 3.015 2.79 ;
 RECT 2.81 1.14 3.04 1.37 ;
 RECT 1.85 0.09 1.95 1.065 ;
 RECT 1.85 1.295 1.95 2.79 ;
 RECT 1.85 1.065 2.08 1.295 ;
 RECT 2.345 0.09 2.445 0.83 ;
 RECT 2.345 0.83 2.59 1.06 ;
 RECT 2.345 1.06 2.445 2.79 ;
 LAYER CO ;
 RECT 3.165 2.375 3.295 2.505 ;
 RECT 0.63 0.325 0.76 0.455 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 0.725 1.19 0.855 1.32 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 0.61 1.875 0.74 2.005 ;
 RECT 2.65 2.275 2.78 2.405 ;
 RECT 2.07 0.325 2.2 0.455 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 3.165 0.59 3.295 0.72 ;
 RECT 1.255 1.19 1.385 1.32 ;
 RECT 2.41 0.88 2.54 1.01 ;
 RECT 1.59 0.325 1.72 0.455 ;
 RECT 1.9 1.115 2.03 1.245 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 3.165 0.325 3.295 0.455 ;
 RECT 3.165 1.855 3.295 1.985 ;
 RECT 2.655 0.325 2.785 0.455 ;
 RECT 1.11 0.325 1.24 0.455 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 2.86 1.19 2.99 1.32 ;
 RECT 3.165 2.115 3.295 2.245 ;
 RECT 3.165 1.595 3.295 1.725 ;
 LAYER M1 ;
 RECT 1.595 0.665 1.735 1.87 ;
 RECT 0.555 1.87 1.735 2.01 ;
 RECT 1.105 0.255 1.245 0.605 ;
 RECT 2.065 0.255 2.205 0.605 ;
 RECT 1.105 0.605 2.205 0.745 ;
 RECT 1.615 1.87 2.995 2.01 ;
 RECT 2.855 1.17 2.995 1.87 ;
 RECT 2.845 1.14 3 1.37 ;
 END
END OR4X1

MACRO OR4X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.16 BY 2.88 ;
 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.345 0.825 2.68 1.08 ;
 END
 ANTENNAGATEAREA 0.13 ;
 END IN4

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.815 1.065 2.2 1.4 ;
 END
 ANTENNAGATEAREA 0.13 ;
 END IN3

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.16 2.96 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 2.645 2.17 2.785 2.8 ;
 RECT 3.635 2.17 3.775 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.52 1.08 0.86 1.4 ;
 END
 ANTENNAGATEAREA 0.13 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 1.14 1.395 1.4 ;
 END
 ANTENNAGATEAREA 0.13 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.16 1.08 3.3 2.245 ;
 RECT 3.16 0.835 3.48 1.08 ;
 RECT 3.16 0.275 3.3 0.835 ;
 END
 ANTENNADIFFAREA 0.704 ;
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.16 0.08 ;
 RECT 0.625 0.08 0.765 0.505 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 1.575 0.08 1.735 0.505 ;
 RECT 2.65 0.08 2.79 0.505 ;
 RECT 3.64 0.08 3.78 0.505 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 3.415 0.09 3.515 1.19 ;
 RECT 2.81 1.19 3.515 1.29 ;
 RECT 3.415 1.29 3.515 2.76 ;
 RECT 2.915 0.09 3.015 1.12 ;
 RECT 2.81 1.12 3.04 1.19 ;
 RECT 2.81 1.29 3.04 1.35 ;
 RECT 2.915 1.35 3.015 2.76 ;
 RECT 0.675 1.14 0.98 1.37 ;
 RECT 0.88 0.105 0.98 1.14 ;
 RECT 0.88 1.37 0.98 2.755 ;
 RECT 1.205 1.14 1.465 1.37 ;
 RECT 1.365 0.105 1.465 1.14 ;
 RECT 1.365 1.37 1.465 2.745 ;
 RECT 1.85 0.105 1.95 1.065 ;
 RECT 1.85 1.295 1.95 2.75 ;
 RECT 1.85 1.065 2.08 1.295 ;
 RECT 2.345 0.105 2.445 0.84 ;
 RECT 2.345 1.07 2.445 2.755 ;
 RECT 2.345 0.84 2.575 1.07 ;
 LAYER CO ;
 RECT 3.645 0.325 3.775 0.455 ;
 RECT 3.64 2.225 3.77 2.355 ;
 RECT 1.59 0.325 1.72 0.455 ;
 RECT 1.9 1.115 2.03 1.245 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 1.255 1.19 1.385 1.32 ;
 RECT 0.725 1.19 0.855 1.32 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 2.395 0.89 2.525 1.02 ;
 RECT 3.165 1.805 3.295 1.935 ;
 RECT 3.165 2.065 3.295 2.195 ;
 RECT 0.63 0.325 0.76 0.455 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 3.165 0.59 3.295 0.72 ;
 RECT 3.165 0.325 3.295 0.455 ;
 RECT 0.605 1.545 0.735 1.675 ;
 RECT 2.65 2.225 2.78 2.355 ;
 RECT 2.86 1.17 2.99 1.3 ;
 RECT 1.11 0.325 1.24 0.455 ;
 RECT 2.655 0.325 2.785 0.455 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 2.07 0.325 2.2 0.455 ;
 RECT 3.165 1.545 3.295 1.675 ;
 LAYER M1 ;
 RECT 1.535 0.665 1.675 1.54 ;
 RECT 0.555 1.54 1.675 1.68 ;
 RECT 1.105 0.275 1.245 0.645 ;
 RECT 2.065 0.27 2.205 0.645 ;
 RECT 1.105 0.645 2.205 0.785 ;
 RECT 1.615 1.54 2.995 1.68 ;
 RECT 2.855 1.17 2.995 1.54 ;
 RECT 2.845 1.12 3 1.35 ;
 END
END OR4X2

MACRO OR4X4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.12 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.12 0.08 ;
 RECT 0.625 0.08 0.765 0.505 ;
 RECT 1.575 0.08 1.735 0.505 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 3.64 0.08 3.78 0.83 ;
 RECT 2.65 0.08 2.79 0.505 ;
 RECT 4.605 0.08 4.745 0.9 ;
 END
 END VSS

 PIN IN4
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.345 0.805 2.68 1.135 ;
 END
 ANTENNAGATEAREA 0.128 ;
 END IN4

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1 1.14 1.395 1.4 ;
 END
 ANTENNAGATEAREA 0.128 ;
 END IN2

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.12 2.96 ;
 RECT 4.595 1.51 4.735 2.8 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 3.635 1.47 3.775 2.8 ;
 RECT 2.645 1.82 2.785 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.115 1.325 4.255 2.245 ;
 RECT 4.115 0.275 4.255 1.185 ;
 RECT 3.16 1.185 4.255 1.325 ;
 RECT 3.16 1.4 3.3 2.585 ;
 RECT 3.16 1.325 3.505 1.4 ;
 RECT 3.16 0.275 3.3 1.135 ;
 RECT 3.16 1.135 3.505 1.185 ;
 END
 ANTENNADIFFAREA 1.382 ;
 END Q

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.52 1.14 0.86 1.4 ;
 END
 ANTENNAGATEAREA 0.128 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.89 1.065 2.205 1.4 ;
 END
 ANTENNAGATEAREA 0.128 ;
 END IN3

 OBS
 LAYER PO ;
 RECT 1.205 1.14 1.465 1.37 ;
 RECT 1.365 0.105 1.465 1.14 ;
 RECT 1.365 1.37 1.465 2.745 ;
 RECT 0.675 1.14 0.98 1.37 ;
 RECT 0.88 0.105 0.98 1.14 ;
 RECT 0.88 1.37 0.98 2.755 ;
 RECT 2.915 0.09 3.015 1.12 ;
 RECT 4.38 0.09 4.48 1.19 ;
 RECT 4.38 1.29 4.48 2.76 ;
 RECT 3.895 0.09 3.995 1.19 ;
 RECT 3.895 1.29 3.995 2.76 ;
 RECT 3.415 0.09 3.515 1.19 ;
 RECT 3.415 1.29 3.515 2.76 ;
 RECT 2.915 1.35 3.015 2.76 ;
 RECT 2.81 1.12 3.04 1.19 ;
 RECT 2.81 1.19 4.5 1.29 ;
 RECT 2.81 1.29 3.04 1.35 ;
 RECT 1.85 0.105 1.95 1.065 ;
 RECT 1.85 1.295 1.95 2.75 ;
 RECT 1.85 1.065 2.08 1.295 ;
 RECT 2.345 0.105 2.445 0.89 ;
 RECT 2.345 1.12 2.445 2.755 ;
 RECT 2.345 0.89 2.575 1.12 ;
 LAYER CO ;
 RECT 0.63 0.325 0.76 0.455 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 0.725 1.19 0.855 1.32 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 2.65 2.37 2.78 2.5 ;
 RECT 2.07 0.325 2.2 0.455 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 3.165 0.59 3.295 0.72 ;
 RECT 1.255 1.19 1.385 1.32 ;
 RECT 3.64 2.36 3.77 2.49 ;
 RECT 2.395 0.94 2.525 1.07 ;
 RECT 1.59 0.325 1.72 0.455 ;
 RECT 1.9 1.115 2.03 1.245 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 3.165 0.325 3.295 0.455 ;
 RECT 3.165 1.805 3.295 1.935 ;
 RECT 3.645 0.325 3.775 0.455 ;
 RECT 2.655 0.325 2.785 0.455 ;
 RECT 1.11 0.325 1.24 0.455 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 2.86 1.17 2.99 1.3 ;
 RECT 3.165 2.065 3.295 2.195 ;
 RECT 3.165 1.545 3.295 1.675 ;
 RECT 4.61 0.59 4.74 0.72 ;
 RECT 3.645 0.585 3.775 0.715 ;
 RECT 0.605 2.365 0.735 2.495 ;
 RECT 0.605 2.08 0.735 2.21 ;
 RECT 0.605 1.815 0.735 1.945 ;
 RECT 4.6 1.695 4.73 1.825 ;
 RECT 4.6 1.96 4.73 2.09 ;
 RECT 2.65 2.11 2.78 2.24 ;
 RECT 3.165 2.33 3.295 2.46 ;
 RECT 3.64 1.58 3.77 1.71 ;
 RECT 3.64 1.84 3.77 1.97 ;
 RECT 3.64 2.1 3.77 2.23 ;
 RECT 4.61 0.325 4.74 0.455 ;
 RECT 4.6 2.225 4.73 2.355 ;
 RECT 4.12 0.59 4.25 0.72 ;
 RECT 4.12 0.325 4.25 0.455 ;
 RECT 4.12 1.805 4.25 1.935 ;
 RECT 4.12 2.065 4.25 2.195 ;
 RECT 4.12 1.545 4.25 1.675 ;
 LAYER M1 ;
 RECT 0.6 1.54 0.74 2.63 ;
 RECT 1.595 0.665 1.735 1.54 ;
 RECT 0.6 1.54 1.735 1.68 ;
 RECT 1.105 0.275 1.245 0.645 ;
 RECT 2.065 0.27 2.205 0.645 ;
 RECT 1.105 0.645 2.205 0.785 ;
 RECT 1.615 1.54 2.995 1.68 ;
 RECT 2.855 1.17 2.995 1.54 ;
 RECT 2.845 1.12 3 1.35 ;
 END
END OR4X4

MACRO RDFFARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 21.44 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.955 0.79 3.505 1.135 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.795 1.14 1.1 1.49 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END RSTB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.18 0.865 8.465 1.08 ;
 RECT 8.18 1.08 8.46 1.1 ;
 RECT 8.18 0.82 8.46 0.865 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.565 1.5 10.705 2.295 ;
 RECT 10.565 1.09 11.105 1.5 ;
 RECT 10.565 0.525 10.705 1.09 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.615 1.485 11.755 1.79 ;
 RECT 11.615 1.095 12.065 1.485 ;
 RECT 11.615 0.43 11.755 1.095 ;
 END
 ANTENNADIFFAREA 0.471 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 21.44 2.96 ;
 RECT 6.325 2.615 6.56 2.8 ;
 RECT 2.675 2.51 2.945 2.65 ;
 RECT 4.37 2.51 4.6 2.65 ;
 RECT 8.425 2.37 8.695 2.51 ;
 RECT 13.865 2.025 14.005 2.8 ;
 RECT 0.67 1.855 0.81 2.8 ;
 RECT 11.135 2.275 11.275 2.8 ;
 RECT 12.175 2 12.315 2.8 ;
 RECT 0.265 1.64 0.425 2.8 ;
 RECT 9.62 1.94 9.76 2.8 ;
 RECT 2.74 2.65 2.88 2.8 ;
 RECT 4.415 2.65 4.555 2.8 ;
 RECT 8.49 2.51 8.63 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 21.44 0.08 ;
 RECT 8.37 0.32 8.64 0.46 ;
 RECT 16.275 0.22 16.525 0.36 ;
 RECT 4.38 0.555 4.63 0.695 ;
 RECT 2.74 0.08 2.88 0.32 ;
 RECT 13.865 0.08 14.005 0.815 ;
 RECT 0.265 0.08 0.425 0.84 ;
 RECT 7.53 0.08 7.67 0.78 ;
 RECT 1.645 0.08 1.785 0.8 ;
 RECT 6.39 0.08 6.53 0.78 ;
 RECT 11.135 0.08 11.275 0.575 ;
 RECT 0.705 0.08 0.845 0.79 ;
 RECT 19.04 0.08 19.18 0.65 ;
 RECT 12.225 0.08 12.365 0.865 ;
 RECT 9.62 0.08 9.76 0.785 ;
 RECT 8.435 0.46 8.575 0.525 ;
 RECT 8.435 0.08 8.575 0.32 ;
 RECT 16.32 0.08 16.46 0.22 ;
 RECT 4.445 0.08 4.585 0.555 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 19.895 1.4 20.235 1.765 ;
 RECT 16.275 1.47 16.505 1.61 ;
 RECT 16.325 2.31 20.05 2.385 ;
 RECT 16.32 2.225 20.05 2.31 ;
 RECT 16.32 1.61 16.46 2.225 ;
 RECT 18.995 1.395 19.135 2.225 ;
 RECT 19.91 1.765 20.05 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.78 0.75 15.285 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 17.18 2.09 18.315 2.19 ;
 RECT 16.025 1.76 17.28 1.86 ;
 RECT 16.605 0.965 16.705 1.145 ;
 RECT 18.215 0.275 18.315 0.865 ;
 RECT 17.935 0.965 18.035 1.145 ;
 RECT 17.745 1.245 17.845 1.86 ;
 RECT 16.605 1.145 18.035 1.245 ;
 RECT 17.935 0.865 18.315 0.965 ;
 RECT 16.605 0.735 16.835 0.965 ;
 RECT 3.085 1.76 3.185 2.34 ;
 RECT 2.965 1.53 3.195 1.76 ;
 RECT 12.51 0.385 12.61 2.405 ;
 RECT 12.41 2.405 12.64 2.635 ;
 RECT 12.82 1.835 12.92 2.425 ;
 RECT 12.81 1.605 13.04 1.835 ;
 RECT 17.03 0.865 17.755 0.965 ;
 RECT 17.03 0.735 17.26 0.865 ;
 RECT 17.655 0.275 17.755 0.865 ;
 RECT 2.995 0.1 5.69 0.2 ;
 RECT 5.59 0.42 5.69 0.95 ;
 RECT 5.39 0.2 5.69 0.42 ;
 RECT 2.995 0.2 3.095 0.97 ;
 RECT 8.175 0.33 8.275 0.865 ;
 RECT 8.175 0.865 8.465 1.08 ;
 RECT 8.175 1.08 8.275 2.235 ;
 RECT 8.755 0.33 8.855 1.27 ;
 RECT 8.455 1.27 8.855 1.49 ;
 RECT 8.755 1.49 8.855 2.235 ;
 RECT 6.65 0.37 6.75 2.28 ;
 RECT 6.54 2.28 6.77 2.51 ;
 RECT 5.515 1.445 5.615 2.035 ;
 RECT 5.43 2.035 5.66 2.265 ;
 RECT 3.92 1.34 4.15 1.45 ;
 RECT 3.92 0.38 4.02 1.24 ;
 RECT 3.92 1.45 4.02 2.345 ;
 RECT 5.015 0.38 5.115 1.24 ;
 RECT 5.015 1.34 5.115 2.42 ;
 RECT 3.92 1.24 5.115 1.34 ;
 RECT 18.69 0.275 18.79 1.025 ;
 RECT 18.69 1.255 18.79 1.86 ;
 RECT 18.69 1.025 18.97 1.255 ;
 RECT 4.225 0.84 4.47 0.87 ;
 RECT 4.225 0.97 4.47 1.06 ;
 RECT 4.225 0.38 4.325 0.84 ;
 RECT 4.7 0.38 4.8 0.87 ;
 RECT 4.225 0.87 4.8 0.97 ;
 RECT 6.12 0.37 6.22 1.21 ;
 RECT 6.12 1.42 6.22 2.16 ;
 RECT 6.12 1.21 6.405 1.42 ;
 RECT 13.305 0.205 13.405 0.925 ;
 RECT 11.4 0.105 14.775 0.205 ;
 RECT 11.4 0.205 11.5 0.87 ;
 RECT 14.545 0.205 14.775 0.4 ;
 RECT 11.4 1.085 11.5 2.755 ;
 RECT 11.255 0.87 11.5 1.085 ;
 RECT 13.18 0.925 13.41 1.135 ;
 RECT 3.395 0.38 3.495 0.865 ;
 RECT 3.395 1.095 3.495 2.36 ;
 RECT 3.275 0.865 3.505 1.095 ;
 RECT 2.5 0.38 2.6 1.23 ;
 RECT 2.5 1.46 2.6 2.34 ;
 RECT 2.5 1.23 2.73 1.46 ;
 RECT 2.18 1.095 2.28 2.325 ;
 RECT 1.91 0.38 2.01 0.995 ;
 RECT 2.05 2.325 2.28 2.555 ;
 RECT 1.91 0.995 2.28 1.095 ;
 RECT 19.295 0.27 19.395 0.745 ;
 RECT 19.295 0.975 19.395 1.855 ;
 RECT 19.15 0.745 19.395 0.975 ;
 RECT 6.95 1.06 7.05 2.68 ;
 RECT 7.26 0.37 7.36 0.96 ;
 RECT 9.13 2.475 9.36 2.68 ;
 RECT 6.95 0.96 7.36 1.06 ;
 RECT 6.95 2.68 9.36 2.78 ;
 RECT 0.975 0.35 1.075 1.255 ;
 RECT 0.845 1.255 1.075 1.485 ;
 RECT 0.975 1.485 1.075 2.485 ;
 RECT 13.35 2.605 14.7 2.695 ;
 RECT 13.35 1.425 13.45 2.605 ;
 RECT 13.355 2.695 14.7 2.705 ;
 RECT 12.815 0.385 12.915 1.325 ;
 RECT 14.47 2.475 14.7 2.605 ;
 RECT 12.815 1.325 13.45 1.425 ;
 RECT 9.715 1.16 10.01 1.22 ;
 RECT 9.91 0.365 10.01 1.16 ;
 RECT 9.91 1.39 10.01 2.47 ;
 RECT 9.715 1.32 10.01 1.39 ;
 RECT 9.715 1.22 10.92 1.32 ;
 RECT 10.82 0.105 10.92 1.22 ;
 RECT 10.82 1.32 10.92 2.75 ;
 RECT 4.69 1.75 4.79 2.42 ;
 RECT 4.56 1.53 4.79 1.63 ;
 RECT 4.56 1.73 4.79 1.75 ;
 RECT 4.22 1.73 4.32 2.34 ;
 RECT 4.22 1.63 4.79 1.73 ;
 RECT 16.025 0.145 16.125 0.945 ;
 RECT 14.125 0.945 16.125 1.045 ;
 RECT 16.025 1.045 16.125 1.76 ;
 RECT 13.65 0.385 13.75 1.215 ;
 RECT 13.65 1.215 13.925 1.27 ;
 RECT 13.65 1.425 13.75 2.425 ;
 RECT 13.65 1.37 13.925 1.425 ;
 RECT 14.125 1.045 14.225 1.27 ;
 RECT 13.65 1.27 14.225 1.37 ;
 RECT 14.125 1.37 14.225 2.425 ;
 RECT 18.215 1.145 18.315 2.09 ;
 RECT 17.18 1.86 17.28 2.09 ;
 RECT 17.05 1.545 17.28 1.76 ;
 RECT 14.87 0.84 15.1 0.945 ;
 RECT 14.87 1.045 15.1 1.07 ;
 RECT 14.125 0.385 14.225 0.945 ;
 LAYER CO ;
 RECT 6.59 2.33 6.72 2.46 ;
 RECT 19.945 1.44 20.075 1.57 ;
 RECT 0.28 0.36 0.41 0.49 ;
 RECT 0.28 0.62 0.41 0.75 ;
 RECT 0.28 1.71 0.41 1.84 ;
 RECT 3.325 0.915 3.455 1.045 ;
 RECT 2.55 1.28 2.68 1.41 ;
 RECT 2.1 2.375 2.23 2.505 ;
 RECT 9.065 0.57 9.195 0.7 ;
 RECT 9.065 1.64 9.195 1.77 ;
 RECT 8.44 0.325 8.57 0.455 ;
 RECT 7.905 0.57 8.035 0.7 ;
 RECT 7.925 1.48 8.055 1.61 ;
 RECT 8.495 2.375 8.625 2.505 ;
 RECT 6.38 2.63 6.51 2.76 ;
 RECT 1.93 1.585 2.06 1.715 ;
 RECT 0.885 1.305 1.015 1.435 ;
 RECT 11.14 0.395 11.27 0.525 ;
 RECT 10.57 0.585 10.7 0.715 ;
 RECT 10.57 2.105 10.7 2.235 ;
 RECT 11.14 2.34 11.27 2.47 ;
 RECT 14.92 0.89 15.05 1.02 ;
 RECT 17.1 1.595 17.23 1.725 ;
 RECT 16.655 0.785 16.785 0.915 ;
 RECT 2.745 0.12 2.875 0.25 ;
 RECT 5.48 2.085 5.61 2.215 ;
 RECT 5.44 0.24 5.57 0.37 ;
 RECT 5.26 1.67 5.39 1.8 ;
 RECT 2.745 2.515 2.875 2.645 ;
 RECT 4.42 2.515 4.55 2.645 ;
 RECT 3.65 1.52 3.78 1.65 ;
 RECT 7.18 1.49 7.31 1.62 ;
 RECT 7.535 0.6 7.665 0.73 ;
 RECT 13.055 2.05 13.185 2.18 ;
 RECT 13.055 0.635 13.185 0.765 ;
 RECT 17.08 0.785 17.21 0.915 ;
 RECT 19.2 0.795 19.33 0.925 ;
 RECT 0.28 1.97 0.41 2.1 ;
 RECT 0.28 2.23 0.41 2.36 ;
 RECT 16.325 0.225 16.455 0.355 ;
 RECT 13.23 0.965 13.36 1.095 ;
 RECT 12.23 0.635 12.36 0.765 ;
 RECT 12.18 2.06 12.31 2.19 ;
 RECT 14.35 2.065 14.48 2.195 ;
 RECT 10.57 1.715 10.7 1.845 ;
 RECT 18.79 1.075 18.92 1.205 ;
 RECT 19.525 0.505 19.655 0.635 ;
 RECT 19.525 1.44 19.655 1.57 ;
 RECT 19.045 0.47 19.175 0.6 ;
 RECT 19 1.455 19.13 1.585 ;
 RECT 18.44 1.435 18.57 1.565 ;
 RECT 18.44 0.505 18.57 0.635 ;
 RECT 17.965 1.415 18.095 1.545 ;
 RECT 2.13 0.6 2.26 0.73 ;
 RECT 1.27 1.875 1.4 2.005 ;
 RECT 1.27 0.58 1.4 0.71 ;
 RECT 0.71 0.59 0.84 0.72 ;
 RECT 0.675 1.905 0.805 2.035 ;
 RECT 6.225 1.25 6.355 1.38 ;
 RECT 4.61 1.57 4.74 1.7 ;
 RECT 4.28 0.89 4.41 1.02 ;
 RECT 3.97 1.28 4.1 1.41 ;
 RECT 3.015 1.58 3.145 1.71 ;
 RECT 6.955 0.6 7.085 0.73 ;
 RECT 6.395 0.6 6.525 0.73 ;
 RECT 5.82 0.6 5.95 0.73 ;
 RECT 5.82 1.48 5.95 1.61 ;
 RECT 5.26 0.6 5.39 0.73 ;
 RECT 4.45 0.555 4.58 0.685 ;
 RECT 3.65 0.6 3.78 0.73 ;
 RECT 1.65 0.6 1.78 0.73 ;
 RECT 14.595 0.225 14.725 0.355 ;
 RECT 16.325 1.475 16.455 1.605 ;
 RECT 15.72 1.255 15.85 1.385 ;
 RECT 15.675 0.505 15.805 0.635 ;
 RECT 14.52 2.525 14.65 2.655 ;
 RECT 12.46 2.455 12.59 2.585 ;
 RECT 12.86 1.655 12.99 1.785 ;
 RECT 14.35 0.635 14.48 0.765 ;
 RECT 13.87 0.635 14 0.765 ;
 RECT 13.87 2.075 14 2.205 ;
 RECT 13.745 1.255 13.875 1.385 ;
 RECT 9.18 2.525 9.31 2.655 ;
 RECT 11.305 0.915 11.435 1.045 ;
 RECT 11.62 1.6 11.75 1.73 ;
 RECT 17.965 0.505 18.095 0.635 ;
 RECT 17.405 1.415 17.535 1.545 ;
 RECT 17.405 0.505 17.535 0.635 ;
 RECT 11.62 0.51 11.75 0.64 ;
 RECT 9.625 2.01 9.755 2.14 ;
 RECT 9.765 1.21 9.895 1.34 ;
 RECT 9.625 0.605 9.755 0.735 ;
 RECT 10.185 2.025 10.315 2.155 ;
 RECT 10.185 0.605 10.315 0.735 ;
 RECT 8.285 0.91 8.415 1.04 ;
 RECT 8.505 1.31 8.635 1.44 ;
 LAYER M1 ;
 RECT 17.095 0.92 17.235 1.785 ;
 RECT 17.01 0.78 17.26 0.92 ;
 RECT 13.65 1.17 13.99 1.51 ;
 RECT 5.815 0.55 5.955 1.475 ;
 RECT 5.75 1.475 6.02 1.615 ;
 RECT 19.52 0.435 19.66 1.07 ;
 RECT 18.72 1.07 19.66 1.21 ;
 RECT 19.52 1.21 19.66 1.64 ;
 RECT 13.49 1.845 13.63 2.45 ;
 RECT 12.455 2.385 12.595 2.45 ;
 RECT 12.455 2.45 13.63 2.59 ;
 RECT 12.455 2.59 12.595 2.65 ;
 RECT 14.345 0.585 14.485 1.705 ;
 RECT 13.49 1.705 14.485 1.845 ;
 RECT 14.345 1.845 14.485 2.265 ;
 RECT 14.495 0.235 16.135 0.36 ;
 RECT 14.495 0.22 16.085 0.235 ;
 RECT 15.995 0.36 16.135 0.5 ;
 RECT 17.4 0.435 17.54 0.5 ;
 RECT 17.4 0.64 17.54 1.61 ;
 RECT 15.995 0.5 17.54 0.64 ;
 RECT 3.645 0.55 3.785 1.275 ;
 RECT 2.5 1.275 3.785 1.415 ;
 RECT 3.645 1.415 3.785 1.71 ;
 RECT 1.265 2.37 2.46 2.51 ;
 RECT 1.265 0.53 1.405 2.37 ;
 RECT 2.32 2.23 5 2.37 ;
 RECT 4.86 2.465 6.145 2.51 ;
 RECT 4.86 2.37 6.78 2.465 ;
 RECT 6.005 2.325 6.78 2.37 ;
 RECT 9.9 1.775 10.04 2.435 ;
 RECT 9.34 1.635 10.04 1.775 ;
 RECT 9.34 1.775 9.48 2.52 ;
 RECT 9.11 2.52 9.48 2.66 ;
 RECT 11.895 1.86 12.035 1.995 ;
 RECT 10.855 1.995 12.035 2.135 ;
 RECT 10.855 2.135 10.995 2.435 ;
 RECT 9.9 2.435 10.995 2.575 ;
 RECT 12.57 0.63 13.235 0.77 ;
 RECT 12.57 0.77 12.71 1.72 ;
 RECT 12.57 2.045 13.235 2.185 ;
 RECT 12.57 1.86 12.71 2.045 ;
 RECT 11.895 1.72 12.71 1.86 ;
 RECT 15.995 1.33 16.135 2.52 ;
 RECT 14.44 2.52 16.135 2.66 ;
 RECT 18.435 0.64 18.575 1.925 ;
 RECT 16.645 1.33 16.785 1.925 ;
 RECT 18.37 0.5 18.62 0.64 ;
 RECT 16.645 1.925 18.575 2.065 ;
 RECT 15.995 1.19 16.785 1.33 ;
 RECT 1.925 0.6 2.33 0.735 ;
 RECT 1.925 0.735 2.065 1.765 ;
 RECT 3.205 0.41 3.345 0.46 ;
 RECT 1.925 0.595 3.345 0.6 ;
 RECT 2.13 0.46 3.345 0.595 ;
 RECT 3.205 0.27 4.105 0.41 ;
 RECT 3.965 0.41 4.105 1.475 ;
 RECT 5.185 1.765 7.78 1.8 ;
 RECT 5.185 1.665 5.61 1.765 ;
 RECT 5.255 0.545 5.395 1.665 ;
 RECT 9.34 0.365 9.48 1.205 ;
 RECT 5.47 1.805 8.92 1.905 ;
 RECT 5.185 1.8 8.92 1.805 ;
 RECT 8.78 0.365 8.92 1.8 ;
 RECT 8.78 0.225 9.48 0.365 ;
 RECT 7.64 1.905 8.92 1.94 ;
 RECT 9.34 1.205 9.965 1.345 ;
 RECT 18.76 0.36 18.9 0.79 ;
 RECT 17.96 0.36 18.1 1.41 ;
 RECT 17.895 1.41 18.165 1.55 ;
 RECT 17.96 0.22 18.9 0.36 ;
 RECT 18.76 0.79 19.38 0.93 ;
 RECT 6.175 1.21 6.405 1.245 ;
 RECT 6.175 1.385 6.405 1.42 ;
 RECT 6.175 1.245 7.36 1.385 ;
 RECT 7.13 1.385 7.36 1.625 ;
 RECT 6.95 0.55 7.09 1.245 ;
 RECT 7.575 1.065 7.715 1.305 ;
 RECT 7.25 0.925 8.04 0.99 ;
 RECT 7.25 0.99 8.035 1.065 ;
 RECT 7.9 0.515 8.04 0.925 ;
 RECT 7.92 1.445 8.06 1.66 ;
 RECT 6.67 0.38 6.81 0.93 ;
 RECT 7.25 0.38 7.39 0.925 ;
 RECT 6.67 0.24 7.39 0.38 ;
 RECT 6.105 0.93 6.81 1.07 ;
 RECT 4.775 0.375 4.915 1.26 ;
 RECT 6.105 0.375 6.245 0.93 ;
 RECT 4.605 1.26 4.915 1.4 ;
 RECT 4.605 1.4 4.745 1.77 ;
 RECT 4.775 0.235 6.245 0.375 ;
 RECT 8.5 1.26 8.64 1.305 ;
 RECT 8.5 1.445 8.64 1.495 ;
 RECT 7.575 1.305 8.64 1.445 ;
 RECT 5.14 2.085 7.445 2.09 ;
 RECT 5.43 2.045 7.445 2.08 ;
 RECT 3.01 2.08 7.445 2.085 ;
 RECT 3.01 1.945 5.28 2.08 ;
 RECT 5.14 2.185 5.66 2.22 ;
 RECT 4.275 0.835 4.415 1.945 ;
 RECT 3.01 1.715 3.15 1.945 ;
 RECT 2.94 1.575 3.215 1.715 ;
 RECT 5.14 2.09 9.2 2.185 ;
 RECT 7.305 2.185 9.2 2.23 ;
 RECT 9.06 0.52 9.2 2.09 ;
 RECT 13.18 0.925 13.41 0.955 ;
 RECT 12.855 0.955 13.41 1.095 ;
 RECT 13.18 1.095 13.41 1.135 ;
 RECT 12.855 1.095 12.995 1.835 ;
 RECT 10.18 0.385 10.32 2.21 ;
 RECT 10.845 0.385 10.985 0.75 ;
 RECT 10.18 0.245 10.985 0.385 ;
 RECT 11.3 0.89 11.44 1.095 ;
 RECT 10.845 0.75 11.44 0.89 ;
 RECT 15.715 0.64 15.855 0.78 ;
 RECT 15.715 0.92 15.855 1.455 ;
 RECT 15.61 0.5 15.855 0.64 ;
 RECT 15.715 0.78 16.85 0.92 ;
 END
END RDFFARX1

MACRO RDFFARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 23.04 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.055 0.815 3.505 1.135 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.75 1.44 1.11 1.75 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END RSTB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.18 0.815 8.55 1.12 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.025 1.09 11.43 1.5 ;
 RECT 11.29 1.5 11.43 1.785 ;
 RECT 11.29 0.51 11.43 1.09 ;
 END
 ANTENNADIFFAREA 0.584 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.34 1.12 12.705 1.465 ;
 RECT 12.34 1.465 12.48 1.79 ;
 RECT 12.34 0.48 12.48 1.12 ;
 END
 ANTENNADIFFAREA 0.626 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 23.04 2.96 ;
 RECT 6.325 2.615 6.56 2.8 ;
 RECT 10.745 2.21 11.02 2.35 ;
 RECT 8.425 2.37 8.695 2.51 ;
 RECT 2.675 2.51 2.945 2.65 ;
 RECT 12.765 2.21 13.04 2.35 ;
 RECT 4.37 2.51 4.6 2.65 ;
 RECT 11.79 2.21 12.065 2.35 ;
 RECT 9.62 1.94 9.76 2.8 ;
 RECT 14.94 2.025 15.08 2.8 ;
 RECT 0.265 1.64 0.425 2.8 ;
 RECT 0.67 1.905 0.81 2.8 ;
 RECT 13.25 2 13.39 2.8 ;
 RECT 10.815 2.35 10.955 2.8 ;
 RECT 8.49 2.51 8.63 2.8 ;
 RECT 2.74 2.65 2.88 2.8 ;
 RECT 12.835 2.35 12.975 2.8 ;
 RECT 4.415 2.65 4.555 2.8 ;
 RECT 11.86 2.35 12 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 23.04 0.08 ;
 RECT 17.9 0.22 18.15 0.36 ;
 RECT 8.37 0.51 8.64 0.65 ;
 RECT 4.38 0.555 4.63 0.695 ;
 RECT 10.73 0.08 10.87 0.575 ;
 RECT 11.86 0.08 12 0.575 ;
 RECT 2.74 0.08 2.88 0.32 ;
 RECT 6.39 0.08 6.53 0.78 ;
 RECT 12.83 0.08 12.97 0.575 ;
 RECT 20.665 0.08 20.805 0.65 ;
 RECT 1.645 0.08 1.785 0.8 ;
 RECT 14.94 0.08 15.08 0.815 ;
 RECT 9.62 0.08 9.76 0.785 ;
 RECT 0.705 0.08 0.845 0.79 ;
 RECT 0.265 0.08 0.425 0.84 ;
 RECT 7.53 0.08 7.67 0.78 ;
 RECT 13.3 0.08 13.44 0.865 ;
 RECT 17.945 0.08 18.085 0.22 ;
 RECT 8.435 0.65 8.575 0.67 ;
 RECT 8.435 0.08 8.575 0.51 ;
 RECT 4.445 0.08 4.585 0.555 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 21.48 1.4 21.905 1.765 ;
 RECT 17.9 1.47 18.13 1.61 ;
 RECT 17.95 2.31 21.685 2.385 ;
 RECT 17.945 2.225 21.685 2.31 ;
 RECT 17.945 1.61 18.085 2.225 ;
 RECT 20.62 1.395 20.76 2.225 ;
 RECT 21.535 1.765 21.675 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 16.115 0.81 16.495 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 19.84 1.145 19.94 2.09 ;
 RECT 18.805 1.86 18.905 2.09 ;
 RECT 18.675 1.545 18.905 1.76 ;
 RECT 17.65 1.76 18.905 1.86 ;
 RECT 18.805 2.09 19.94 2.19 ;
 RECT 3.395 0.38 3.495 0.865 ;
 RECT 3.395 1.095 3.495 2.36 ;
 RECT 3.275 0.865 3.505 1.095 ;
 RECT 0.975 0.35 1.075 1.465 ;
 RECT 0.845 1.465 1.075 1.695 ;
 RECT 0.975 1.695 1.075 2.485 ;
 RECT 8.175 0.28 8.275 0.865 ;
 RECT 8.175 0.865 8.465 1.08 ;
 RECT 8.175 1.08 8.275 2.235 ;
 RECT 4.69 1.75 4.79 2.44 ;
 RECT 4.56 1.53 4.79 1.63 ;
 RECT 4.56 1.73 4.79 1.75 ;
 RECT 4.22 1.73 4.32 2.34 ;
 RECT 4.22 1.63 4.79 1.73 ;
 RECT 3.92 1.34 4.15 1.45 ;
 RECT 3.92 0.38 4.02 1.24 ;
 RECT 3.92 1.45 4.02 2.345 ;
 RECT 5.015 0.38 5.115 1.24 ;
 RECT 5.015 1.34 5.115 2.435 ;
 RECT 3.92 1.24 5.115 1.34 ;
 RECT 20.315 0.275 20.415 1.025 ;
 RECT 20.315 1.255 20.415 1.86 ;
 RECT 20.315 1.025 20.595 1.255 ;
 RECT 5.515 1.445 5.615 2.035 ;
 RECT 5.43 2.035 5.66 2.265 ;
 RECT 13.585 0.385 13.685 2.405 ;
 RECT 13.485 2.405 13.715 2.635 ;
 RECT 13.895 1.835 13.995 2.425 ;
 RECT 13.885 1.605 14.115 1.835 ;
 RECT 18.23 0.965 18.33 1.145 ;
 RECT 19.84 0.275 19.94 0.865 ;
 RECT 18.23 1.145 19.66 1.245 ;
 RECT 19.56 0.965 19.66 1.145 ;
 RECT 19.37 1.245 19.47 1.86 ;
 RECT 18.23 0.735 18.46 0.965 ;
 RECT 19.56 0.865 19.94 0.965 ;
 RECT 8.755 0.28 8.855 1.27 ;
 RECT 8.755 1.49 8.855 2.235 ;
 RECT 8.455 1.27 8.855 1.49 ;
 RECT 6.12 0.37 6.22 1.21 ;
 RECT 6.12 1.21 6.405 1.42 ;
 RECT 6.12 1.42 6.22 2.16 ;
 RECT 2.18 1.095 2.28 2.325 ;
 RECT 1.91 0.38 2.01 0.995 ;
 RECT 2.05 2.325 2.28 2.555 ;
 RECT 1.91 0.995 2.28 1.095 ;
 RECT 20.92 0.27 21.02 0.745 ;
 RECT 20.92 0.975 21.02 1.855 ;
 RECT 20.775 0.745 21.02 0.975 ;
 RECT 6.95 1.06 7.05 2.68 ;
 RECT 7.26 0.37 7.36 0.96 ;
 RECT 9.13 2.475 9.36 2.68 ;
 RECT 6.95 0.96 7.36 1.06 ;
 RECT 6.95 2.68 9.36 2.78 ;
 RECT 6.65 0.37 6.75 2.28 ;
 RECT 6.54 2.28 6.77 2.51 ;
 RECT 18.655 0.865 19.38 0.965 ;
 RECT 18.655 0.735 18.885 0.865 ;
 RECT 19.28 0.275 19.38 0.865 ;
 RECT 4.225 0.38 4.325 0.84 ;
 RECT 4.225 0.87 4.8 0.97 ;
 RECT 4.7 0.38 4.8 0.87 ;
 RECT 4.225 0.84 4.47 0.87 ;
 RECT 4.225 0.97 4.47 1.06 ;
 RECT 2.995 0.1 5.69 0.2 ;
 RECT 5.59 0.42 5.69 0.95 ;
 RECT 5.39 0.2 5.69 0.42 ;
 RECT 2.995 0.2 3.095 0.97 ;
 RECT 3.085 1.76 3.185 2.34 ;
 RECT 2.965 1.53 3.195 1.76 ;
 RECT 12.125 1.085 12.225 1.25 ;
 RECT 11.9 0.985 12.225 1.085 ;
 RECT 12.125 0.105 12.225 0.87 ;
 RECT 11.9 0.87 12.225 0.885 ;
 RECT 12.615 0.205 12.715 0.885 ;
 RECT 14.38 0.205 14.48 0.925 ;
 RECT 11.9 0.885 12.715 0.985 ;
 RECT 12.125 1.35 12.225 2.75 ;
 RECT 12.61 1.35 12.71 2.75 ;
 RECT 12.615 0.105 15.85 0.205 ;
 RECT 15.62 0.205 15.85 0.4 ;
 RECT 12.125 1.25 12.71 1.35 ;
 RECT 14.255 0.925 14.485 1.135 ;
 RECT 13.89 0.385 13.99 1.325 ;
 RECT 14.425 2.605 15.775 2.695 ;
 RECT 15.545 2.475 15.775 2.605 ;
 RECT 14.425 1.425 14.525 2.605 ;
 RECT 13.89 1.325 14.525 1.425 ;
 RECT 14.43 2.695 15.775 2.705 ;
 RECT 2.5 0.38 2.6 1.23 ;
 RECT 2.5 1.46 2.6 2.34 ;
 RECT 2.5 1.23 2.73 1.46 ;
 RECT 9.91 0.365 10.01 1.16 ;
 RECT 9.715 1.16 10.01 1.22 ;
 RECT 9.91 1.39 10.01 2.47 ;
 RECT 9.715 1.32 10.01 1.39 ;
 RECT 11.545 0.105 11.645 0.86 ;
 RECT 11.075 0.86 11.645 0.96 ;
 RECT 11.545 0.96 11.645 1.22 ;
 RECT 11.075 0.095 11.175 0.86 ;
 RECT 9.715 1.22 11.645 1.32 ;
 RECT 11.545 1.32 11.645 2.75 ;
 RECT 11.075 1.32 11.175 2.75 ;
 RECT 14.725 1.215 15 1.27 ;
 RECT 14.725 1.37 15 1.425 ;
 RECT 14.725 1.27 15.3 1.37 ;
 RECT 15.2 1.045 15.3 1.27 ;
 RECT 15.2 1.37 15.3 2.425 ;
 RECT 17.65 1.045 17.75 1.76 ;
 RECT 14.725 0.385 14.825 1.215 ;
 RECT 14.725 1.425 14.825 2.425 ;
 RECT 16.205 0.84 16.435 0.945 ;
 RECT 16.205 1.045 16.435 1.07 ;
 RECT 15.2 0.385 15.3 0.945 ;
 RECT 15.2 0.945 17.75 1.045 ;
 RECT 17.65 0.145 17.75 0.945 ;
 LAYER CO ;
 RECT 8.505 1.31 8.635 1.44 ;
 RECT 6.59 2.33 6.72 2.46 ;
 RECT 14.82 1.255 14.95 1.385 ;
 RECT 17.3 0.505 17.43 0.635 ;
 RECT 15.595 2.525 15.725 2.655 ;
 RECT 13.535 2.455 13.665 2.585 ;
 RECT 13.935 1.655 14.065 1.785 ;
 RECT 15.425 0.635 15.555 0.765 ;
 RECT 6.225 1.25 6.355 1.38 ;
 RECT 9.065 0.555 9.195 0.685 ;
 RECT 14.305 0.965 14.435 1.095 ;
 RECT 6.955 0.6 7.085 0.73 ;
 RECT 6.395 0.6 6.525 0.73 ;
 RECT 5.82 0.6 5.95 0.73 ;
 RECT 5.82 1.48 5.95 1.61 ;
 RECT 5.26 0.6 5.39 0.73 ;
 RECT 12.84 2.215 12.97 2.345 ;
 RECT 10.735 0.395 10.865 0.525 ;
 RECT 10.82 2.215 10.95 2.345 ;
 RECT 16.255 0.89 16.385 1.02 ;
 RECT 18.705 0.785 18.835 0.915 ;
 RECT 20.825 0.795 20.955 0.925 ;
 RECT 20.415 1.075 20.545 1.205 ;
 RECT 21.15 0.505 21.28 0.635 ;
 RECT 21.15 1.44 21.28 1.57 ;
 RECT 20.67 0.47 20.8 0.6 ;
 RECT 20.625 1.455 20.755 1.585 ;
 RECT 20.065 1.435 20.195 1.565 ;
 RECT 20.065 0.505 20.195 0.635 ;
 RECT 19.59 1.415 19.72 1.545 ;
 RECT 19.59 0.505 19.72 0.635 ;
 RECT 19.03 1.415 19.16 1.545 ;
 RECT 19.03 0.505 19.16 0.635 ;
 RECT 0.28 0.36 0.41 0.49 ;
 RECT 0.28 0.62 0.41 0.75 ;
 RECT 0.28 1.71 0.41 1.84 ;
 RECT 0.28 1.97 0.41 2.1 ;
 RECT 0.28 2.23 0.41 2.36 ;
 RECT 17.95 0.225 18.08 0.355 ;
 RECT 5.48 2.085 5.61 2.215 ;
 RECT 5.44 0.24 5.57 0.37 ;
 RECT 4.61 1.57 4.74 1.7 ;
 RECT 4.28 0.89 4.41 1.02 ;
 RECT 3.97 1.28 4.1 1.41 ;
 RECT 3.015 1.58 3.145 1.71 ;
 RECT 3.325 0.915 3.455 1.045 ;
 RECT 2.55 1.28 2.68 1.41 ;
 RECT 2.1 2.375 2.23 2.505 ;
 RECT 9.065 1.64 9.195 1.77 ;
 RECT 8.44 0.515 8.57 0.645 ;
 RECT 7.925 0.515 8.055 0.645 ;
 RECT 7.925 1.48 8.055 1.61 ;
 RECT 8.495 2.375 8.625 2.505 ;
 RECT 6.38 2.63 6.51 2.76 ;
 RECT 1.93 1.585 2.06 1.715 ;
 RECT 2.13 0.6 2.26 0.73 ;
 RECT 1.27 1.875 1.4 2.005 ;
 RECT 1.27 0.58 1.4 0.71 ;
 RECT 0.71 0.59 0.84 0.72 ;
 RECT 15.425 2.065 15.555 2.195 ;
 RECT 9.18 2.525 9.31 2.655 ;
 RECT 11.95 0.915 12.08 1.045 ;
 RECT 12.345 1.6 12.475 1.73 ;
 RECT 11.865 0.395 11.995 0.525 ;
 RECT 11.295 0.56 11.425 0.69 ;
 RECT 11.295 1.605 11.425 1.735 ;
 RECT 11.865 2.215 11.995 2.345 ;
 RECT 12.835 0.395 12.965 0.525 ;
 RECT 0.675 2 0.805 2.13 ;
 RECT 5.26 1.67 5.39 1.8 ;
 RECT 2.745 2.515 2.875 2.645 ;
 RECT 4.42 2.515 4.55 2.645 ;
 RECT 3.65 1.52 3.78 1.65 ;
 RECT 7.18 1.49 7.31 1.62 ;
 RECT 7.535 0.6 7.665 0.73 ;
 RECT 4.45 0.555 4.58 0.685 ;
 RECT 3.65 0.6 3.78 0.73 ;
 RECT 1.65 0.6 1.78 0.73 ;
 RECT 15.67 0.225 15.8 0.355 ;
 RECT 17.95 1.475 18.08 1.605 ;
 RECT 17.345 1.255 17.475 1.385 ;
 RECT 18.725 1.595 18.855 1.725 ;
 RECT 18.28 0.785 18.41 0.915 ;
 RECT 2.745 0.12 2.875 0.25 ;
 RECT 21.57 1.44 21.7 1.57 ;
 RECT 14.945 0.635 15.075 0.765 ;
 RECT 14.945 2.075 15.075 2.205 ;
 RECT 14.13 2.05 14.26 2.18 ;
 RECT 14.13 0.635 14.26 0.765 ;
 RECT 13.305 0.635 13.435 0.765 ;
 RECT 13.255 2.06 13.385 2.19 ;
 RECT 0.885 1.515 1.015 1.645 ;
 RECT 12.345 0.555 12.475 0.685 ;
 RECT 9.625 2.01 9.755 2.14 ;
 RECT 9.765 1.21 9.895 1.34 ;
 RECT 9.625 0.605 9.755 0.735 ;
 RECT 10.185 2.025 10.315 2.155 ;
 RECT 10.185 0.605 10.315 0.735 ;
 RECT 8.285 0.91 8.415 1.04 ;
 LAYER M1 ;
 RECT 17.34 0.64 17.48 0.78 ;
 RECT 17.34 0.92 17.48 1.455 ;
 RECT 17.235 0.5 17.48 0.64 ;
 RECT 17.34 0.78 18.475 0.92 ;
 RECT 21.145 0.435 21.285 1.07 ;
 RECT 21.145 1.21 21.285 1.64 ;
 RECT 20.345 1.07 21.285 1.21 ;
 RECT 14.725 1.17 15.065 1.51 ;
 RECT 17.62 0.36 17.76 0.5 ;
 RECT 15.57 0.22 17.76 0.36 ;
 RECT 17.62 0.5 19.165 0.64 ;
 RECT 19.025 0.435 19.165 0.5 ;
 RECT 19.025 0.64 19.165 1.61 ;
 RECT 3.645 0.55 3.785 1.275 ;
 RECT 2.5 1.275 3.785 1.415 ;
 RECT 3.645 1.415 3.785 1.71 ;
 RECT 1.925 0.6 2.33 0.735 ;
 RECT 1.925 0.735 2.065 1.765 ;
 RECT 3.205 0.41 3.345 0.46 ;
 RECT 1.925 0.595 3.345 0.6 ;
 RECT 2.13 0.46 3.345 0.595 ;
 RECT 3.965 0.41 4.105 1.475 ;
 RECT 3.205 0.27 4.105 0.41 ;
 RECT 7.13 1.385 7.36 1.625 ;
 RECT 6.175 1.245 7.36 1.385 ;
 RECT 6.95 0.55 7.09 1.245 ;
 RECT 6.175 1.21 6.405 1.245 ;
 RECT 6.175 1.385 6.405 1.42 ;
 RECT 18.72 0.92 18.86 1.785 ;
 RECT 18.635 0.78 18.885 0.92 ;
 RECT 5.815 0.55 5.955 1.475 ;
 RECT 5.75 1.475 6.02 1.615 ;
 RECT 17.62 1.33 17.76 2.52 ;
 RECT 15.515 2.52 17.76 2.66 ;
 RECT 20.06 0.64 20.2 1.925 ;
 RECT 18.27 1.33 18.41 1.925 ;
 RECT 19.995 0.5 20.245 0.64 ;
 RECT 18.27 1.925 20.2 2.065 ;
 RECT 17.62 1.19 18.41 1.33 ;
 RECT 20.385 0.36 20.525 0.79 ;
 RECT 19.585 0.36 19.725 1.41 ;
 RECT 19.585 0.22 20.525 0.36 ;
 RECT 19.52 1.41 19.79 1.55 ;
 RECT 20.385 0.79 21.005 0.93 ;
 RECT 7.9 0.445 8.04 0.51 ;
 RECT 7.9 0.65 8.04 0.925 ;
 RECT 7.9 1.065 8.04 1.305 ;
 RECT 7.9 1.445 8.125 1.475 ;
 RECT 7.25 0.925 8.04 1.065 ;
 RECT 7.855 1.475 8.125 1.615 ;
 RECT 7.855 0.51 8.125 0.65 ;
 RECT 7.25 0.38 7.39 0.925 ;
 RECT 6.67 0.38 6.81 0.93 ;
 RECT 6.67 0.24 7.39 0.38 ;
 RECT 6.105 0.93 6.81 1.07 ;
 RECT 6.105 0.375 6.245 0.93 ;
 RECT 4.775 0.375 4.915 1.26 ;
 RECT 4.775 0.235 6.245 0.375 ;
 RECT 4.605 1.4 4.745 1.77 ;
 RECT 4.605 1.26 4.915 1.4 ;
 RECT 8.5 1.26 8.64 1.305 ;
 RECT 8.5 1.445 8.64 1.495 ;
 RECT 7.9 1.305 8.64 1.445 ;
 RECT 13.93 1.095 14.07 1.835 ;
 RECT 14.255 0.925 14.485 0.955 ;
 RECT 14.255 1.095 14.485 1.135 ;
 RECT 13.93 0.955 14.485 1.095 ;
 RECT 1.265 2.37 2.46 2.51 ;
 RECT 1.265 0.53 1.405 2.37 ;
 RECT 2.32 2.23 5 2.37 ;
 RECT 4.86 2.465 6.145 2.51 ;
 RECT 4.86 2.37 6.78 2.465 ;
 RECT 6.005 2.325 6.78 2.37 ;
 RECT 10.46 2.07 10.6 2.435 ;
 RECT 9.9 1.775 10.04 2.435 ;
 RECT 9.9 2.435 10.6 2.575 ;
 RECT 9.34 1.635 10.04 1.775 ;
 RECT 9.34 1.775 9.48 2.52 ;
 RECT 9.11 2.52 9.48 2.66 ;
 RECT 10.46 1.93 13.11 2.07 ;
 RECT 12.97 1.86 13.11 1.93 ;
 RECT 13.645 2.045 14.31 2.185 ;
 RECT 13.645 1.86 13.785 2.045 ;
 RECT 13.645 0.63 14.31 0.77 ;
 RECT 13.645 0.77 13.785 1.72 ;
 RECT 12.97 1.72 13.785 1.86 ;
 RECT 10.18 0.775 11.15 0.915 ;
 RECT 11.01 0.36 11.15 0.775 ;
 RECT 10.18 0.55 10.32 0.775 ;
 RECT 10.18 0.915 10.32 2.21 ;
 RECT 11.57 0.36 11.71 0.75 ;
 RECT 11.01 0.22 11.71 0.36 ;
 RECT 11.945 0.89 12.085 1.095 ;
 RECT 11.57 0.75 12.085 0.89 ;
 RECT 5.185 1.765 7.78 1.8 ;
 RECT 5.185 1.665 5.61 1.765 ;
 RECT 5.255 0.545 5.395 1.665 ;
 RECT 5.185 1.8 8.92 1.805 ;
 RECT 5.47 1.805 8.92 1.905 ;
 RECT 9.34 0.365 9.48 1.205 ;
 RECT 8.78 0.365 8.92 1.8 ;
 RECT 7.64 1.905 8.92 1.94 ;
 RECT 8.78 0.225 9.48 0.365 ;
 RECT 9.34 1.205 9.965 1.345 ;
 RECT 3.01 2.08 7.445 2.085 ;
 RECT 5.14 2.085 7.445 2.09 ;
 RECT 5.43 2.045 7.445 2.08 ;
 RECT 3.01 1.945 5.28 2.08 ;
 RECT 5.14 2.185 5.66 2.22 ;
 RECT 4.275 0.835 4.415 1.945 ;
 RECT 3.01 1.715 3.15 1.945 ;
 RECT 2.94 1.575 3.215 1.715 ;
 RECT 5.14 2.09 9.2 2.185 ;
 RECT 7.305 2.185 9.2 2.23 ;
 RECT 9.06 0.505 9.2 2.09 ;
 RECT 14.565 1.845 14.705 2.45 ;
 RECT 13.53 2.385 13.67 2.45 ;
 RECT 13.53 2.45 14.705 2.59 ;
 RECT 13.53 2.59 13.67 2.65 ;
 RECT 15.42 0.585 15.56 1.705 ;
 RECT 14.565 1.705 15.56 1.845 ;
 RECT 15.42 1.845 15.56 2.265 ;
 END
END RDFFARX2

MACRO RDFFNARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 22.08 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.955 0.82 3.505 1.135 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.66 1.055 1.09 1.45 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END RSTB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.18 1.135 8.64 1.425 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 10.565 1.54 10.705 2.295 ;
 RECT 10.565 1.05 11.145 1.54 ;
 RECT 10.565 0.525 10.705 1.05 ;
 END
 ANTENNADIFFAREA 0.504 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.615 1.04 12.115 1.515 ;
 RECT 11.615 1.515 11.755 1.79 ;
 RECT 11.615 0.48 11.755 1.04 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 22.08 2.96 ;
 RECT 0.265 1.64 0.425 2.8 ;
 RECT 6.325 2.615 6.56 2.8 ;
 RECT 4.37 2.51 4.6 2.65 ;
 RECT 2.675 2.51 2.945 2.65 ;
 RECT 8.375 2.37 8.645 2.51 ;
 RECT 0.67 1.855 0.81 2.8 ;
 RECT 9.62 1.94 9.76 2.8 ;
 RECT 11.135 2.275 11.275 2.8 ;
 RECT 12.175 2 12.315 2.8 ;
 RECT 13.865 2.025 14.005 2.8 ;
 RECT 4.415 2.65 4.555 2.8 ;
 RECT 2.74 2.65 2.88 2.8 ;
 RECT 8.44 2.51 8.58 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 22.08 0.08 ;
 RECT 0.265 0.08 0.425 0.84 ;
 RECT 4.38 0.555 4.63 0.695 ;
 RECT 16.28 0.22 16.53 0.36 ;
 RECT 8.37 0.555 8.64 0.695 ;
 RECT 0.705 0.08 0.845 0.79 ;
 RECT 12.225 0.08 12.365 0.865 ;
 RECT 6.39 0.08 6.53 0.78 ;
 RECT 19.045 0.08 19.185 0.65 ;
 RECT 1.645 0.08 1.785 0.8 ;
 RECT 7.53 0.08 7.67 0.78 ;
 RECT 2.74 0.08 2.88 0.32 ;
 RECT 13.865 0.08 14.005 0.815 ;
 RECT 11.135 0.08 11.275 0.575 ;
 RECT 9.62 0.08 9.76 0.785 ;
 RECT 4.445 0.08 4.585 0.555 ;
 RECT 16.325 0.08 16.465 0.22 ;
 RECT 8.435 0.08 8.575 0.555 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 19.9 1.4 20.24 1.765 ;
 RECT 16.325 2.225 20.065 2.385 ;
 RECT 16.28 1.47 16.51 1.61 ;
 RECT 19 1.395 19.14 2.225 ;
 RECT 19.915 1.765 20.055 2.225 ;
 RECT 16.325 1.61 16.465 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.765 0.73 15.315 1.22 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 12.815 0.385 12.915 1.325 ;
 RECT 12.815 1.325 13.45 1.425 ;
 RECT 14.47 2.475 14.7 2.605 ;
 RECT 18.22 0.275 18.32 0.865 ;
 RECT 17.94 0.965 18.04 1.145 ;
 RECT 17.75 1.245 17.85 1.86 ;
 RECT 16.61 0.965 16.71 1.145 ;
 RECT 16.61 1.145 18.04 1.245 ;
 RECT 17.94 0.865 18.32 0.965 ;
 RECT 16.61 0.735 16.84 0.965 ;
 RECT 12.82 1.835 12.92 2.425 ;
 RECT 12.81 1.605 13.04 1.835 ;
 RECT 19.3 0.27 19.4 0.745 ;
 RECT 19.3 0.975 19.4 1.855 ;
 RECT 19.155 0.745 19.4 0.975 ;
 RECT 6.65 0.37 6.75 2.28 ;
 RECT 6.54 2.28 6.77 2.51 ;
 RECT 5.515 1.445 5.615 2.035 ;
 RECT 5.43 2.035 5.66 2.265 ;
 RECT 5.015 0.38 5.115 1.24 ;
 RECT 3.92 1.24 5.115 1.34 ;
 RECT 5.015 1.34 5.115 2.58 ;
 RECT 3.92 1.34 4.15 1.45 ;
 RECT 3.92 0.38 4.02 1.24 ;
 RECT 3.92 1.45 4.02 2.345 ;
 RECT 3.085 1.76 3.185 2.34 ;
 RECT 2.965 1.53 3.195 1.76 ;
 RECT 2.18 1.095 2.28 2.325 ;
 RECT 1.91 0.38 2.01 0.995 ;
 RECT 2.05 2.325 2.28 2.555 ;
 RECT 1.91 0.995 2.28 1.095 ;
 RECT 8.7 0.33 8.8 1.145 ;
 RECT 8.7 1.38 8.8 2.235 ;
 RECT 8.455 1.145 8.8 1.38 ;
 RECT 18.695 0.275 18.795 1.025 ;
 RECT 18.695 1.255 18.795 1.86 ;
 RECT 18.695 1.025 18.975 1.255 ;
 RECT 0.975 0.35 1.075 1.2 ;
 RECT 0.845 1.2 1.075 1.43 ;
 RECT 0.975 1.43 1.075 2.485 ;
 RECT 3.395 0.38 3.495 0.865 ;
 RECT 3.395 1.095 3.495 2.36 ;
 RECT 3.275 0.865 3.505 1.095 ;
 RECT 12.51 0.385 12.61 2.405 ;
 RECT 12.41 2.405 12.64 2.635 ;
 RECT 8.175 0.33 8.275 2.185 ;
 RECT 8.045 2.185 8.275 2.415 ;
 RECT 4.225 0.87 4.8 0.97 ;
 RECT 4.7 0.38 4.8 0.87 ;
 RECT 4.225 0.84 4.47 0.87 ;
 RECT 4.225 0.97 4.47 1.06 ;
 RECT 4.225 0.38 4.325 0.84 ;
 RECT 17.035 0.865 17.76 0.965 ;
 RECT 17.035 0.735 17.265 0.865 ;
 RECT 17.66 0.275 17.76 0.865 ;
 RECT 9.91 0.365 10.01 1.16 ;
 RECT 9.715 1.16 10.01 1.22 ;
 RECT 9.91 1.39 10.01 2.47 ;
 RECT 9.715 1.32 10.01 1.39 ;
 RECT 9.715 1.22 10.92 1.32 ;
 RECT 10.82 0.105 10.92 1.22 ;
 RECT 10.82 1.32 10.92 2.75 ;
 RECT 4.69 1.75 4.79 2.585 ;
 RECT 4.56 1.53 4.79 1.63 ;
 RECT 4.56 1.73 4.79 1.75 ;
 RECT 4.22 1.73 4.32 2.34 ;
 RECT 4.22 1.63 4.79 1.73 ;
 RECT 2.5 0.38 2.6 1.23 ;
 RECT 2.5 1.46 2.6 2.34 ;
 RECT 2.5 1.23 2.73 1.46 ;
 RECT 6.95 1.06 7.05 2.68 ;
 RECT 9.13 2.475 9.36 2.68 ;
 RECT 7.26 0.37 7.36 0.96 ;
 RECT 6.95 2.68 9.36 2.78 ;
 RECT 6.95 0.96 7.36 1.06 ;
 RECT 6.12 0.37 6.22 1.21 ;
 RECT 6.12 1.42 6.22 2.16 ;
 RECT 6.12 1.21 6.405 1.42 ;
 RECT 13.65 0.385 13.75 1.215 ;
 RECT 13.65 1.215 13.925 1.27 ;
 RECT 13.65 1.425 13.75 2.425 ;
 RECT 13.65 1.37 13.925 1.425 ;
 RECT 16.03 0.145 16.13 0.945 ;
 RECT 14.125 0.945 16.13 1.045 ;
 RECT 16.03 1.045 16.13 1.76 ;
 RECT 14.125 1.045 14.225 1.27 ;
 RECT 14.125 1.37 14.225 2.425 ;
 RECT 13.65 1.27 14.225 1.37 ;
 RECT 18.22 1.145 18.32 2.09 ;
 RECT 17.185 1.86 17.285 2.09 ;
 RECT 17.055 1.545 17.285 1.76 ;
 RECT 14.125 0.385 14.225 0.945 ;
 RECT 14.935 0.84 15.165 0.945 ;
 RECT 14.935 1.045 15.165 1.07 ;
 RECT 17.185 2.09 18.32 2.19 ;
 RECT 16.03 1.76 17.285 1.86 ;
 RECT 2.995 0.1 5.69 0.2 ;
 RECT 5.39 0.2 5.69 0.42 ;
 RECT 5.59 0.42 5.69 0.95 ;
 RECT 2.995 0.2 3.095 0.97 ;
 RECT 13.305 0.205 13.405 0.925 ;
 RECT 11.4 0.105 14.775 0.205 ;
 RECT 11.4 0.205 11.5 0.94 ;
 RECT 11.4 1.155 11.5 2.755 ;
 RECT 11.255 0.94 11.5 1.155 ;
 RECT 14.545 0.205 14.775 0.4 ;
 RECT 13.18 0.925 13.41 1.135 ;
 RECT 13.35 2.605 14.7 2.695 ;
 RECT 13.355 2.695 14.7 2.705 ;
 RECT 13.35 1.425 13.45 2.605 ;
 LAYER CO ;
 RECT 0.28 0.36 0.41 0.49 ;
 RECT 0.28 0.62 0.41 0.75 ;
 RECT 0.28 1.71 0.41 1.84 ;
 RECT 0.28 1.97 0.41 2.1 ;
 RECT 0.28 2.23 0.41 2.36 ;
 RECT 16.33 0.225 16.46 0.355 ;
 RECT 2.13 0.6 2.26 0.73 ;
 RECT 1.27 1.875 1.4 2.005 ;
 RECT 1.27 0.58 1.4 0.71 ;
 RECT 0.71 0.59 0.84 0.72 ;
 RECT 0.675 1.905 0.805 2.035 ;
 RECT 5.26 1.67 5.39 1.8 ;
 RECT 2.745 2.515 2.875 2.645 ;
 RECT 4.42 2.515 4.55 2.645 ;
 RECT 3.65 1.52 3.78 1.65 ;
 RECT 7.18 1.49 7.31 1.62 ;
 RECT 7.535 0.6 7.665 0.73 ;
 RECT 6.955 0.6 7.085 0.73 ;
 RECT 6.395 0.6 6.525 0.73 ;
 RECT 5.82 0.6 5.95 0.73 ;
 RECT 5.82 1.48 5.95 1.61 ;
 RECT 5.26 0.6 5.39 0.73 ;
 RECT 4.45 0.555 4.58 0.685 ;
 RECT 3.65 0.6 3.78 0.73 ;
 RECT 1.65 0.6 1.78 0.73 ;
 RECT 14.595 0.225 14.725 0.355 ;
 RECT 16.33 1.475 16.46 1.605 ;
 RECT 15.725 1.255 15.855 1.385 ;
 RECT 15.68 0.505 15.81 0.635 ;
 RECT 10.185 0.605 10.315 0.735 ;
 RECT 7.925 0.57 8.055 0.7 ;
 RECT 7.84 1.48 7.97 1.61 ;
 RECT 8.445 2.375 8.575 2.505 ;
 RECT 12.46 2.455 12.59 2.585 ;
 RECT 12.86 1.655 12.99 1.785 ;
 RECT 14.35 0.635 14.48 0.765 ;
 RECT 13.23 0.965 13.36 1.095 ;
 RECT 6.38 2.63 6.51 2.76 ;
 RECT 13.87 0.635 14 0.765 ;
 RECT 13.87 2.075 14 2.205 ;
 RECT 13.055 2.05 13.185 2.18 ;
 RECT 13.055 0.635 13.185 0.765 ;
 RECT 12.23 0.635 12.36 0.765 ;
 RECT 12.18 2.06 12.31 2.19 ;
 RECT 17.085 0.785 17.215 0.915 ;
 RECT 19.205 0.795 19.335 0.925 ;
 RECT 18.795 1.075 18.925 1.205 ;
 RECT 19.53 0.505 19.66 0.635 ;
 RECT 19.53 1.44 19.66 1.57 ;
 RECT 19.05 0.47 19.18 0.6 ;
 RECT 19.005 1.455 19.135 1.585 ;
 RECT 18.445 1.435 18.575 1.565 ;
 RECT 18.445 0.505 18.575 0.635 ;
 RECT 17.97 1.415 18.1 1.545 ;
 RECT 17.97 0.505 18.1 0.635 ;
 RECT 17.41 1.415 17.54 1.545 ;
 RECT 17.41 0.505 17.54 0.635 ;
 RECT 11.62 0.555 11.75 0.685 ;
 RECT 9.625 2.01 9.755 2.14 ;
 RECT 9.765 1.21 9.895 1.34 ;
 RECT 9.625 0.605 9.755 0.735 ;
 RECT 10.185 2.025 10.315 2.155 ;
 RECT 6.225 1.25 6.355 1.38 ;
 RECT 8.505 1.2 8.635 1.33 ;
 RECT 5.48 2.085 5.61 2.215 ;
 RECT 5.44 0.24 5.57 0.37 ;
 RECT 4.61 1.57 4.74 1.7 ;
 RECT 4.28 0.89 4.41 1.02 ;
 RECT 3.97 1.28 4.1 1.41 ;
 RECT 3.015 1.58 3.145 1.71 ;
 RECT 3.325 0.915 3.455 1.045 ;
 RECT 2.55 1.28 2.68 1.41 ;
 RECT 2.1 2.375 2.23 2.505 ;
 RECT 9.065 0.56 9.195 0.69 ;
 RECT 9.065 1.87 9.195 2 ;
 RECT 8.44 0.56 8.57 0.69 ;
 RECT 13.745 1.255 13.875 1.385 ;
 RECT 0.885 1.25 1.015 1.38 ;
 RECT 1.93 1.585 2.06 1.715 ;
 RECT 14.35 2.065 14.48 2.195 ;
 RECT 10.57 1.715 10.7 1.845 ;
 RECT 9.18 2.525 9.31 2.655 ;
 RECT 11.305 0.985 11.435 1.115 ;
 RECT 11.62 1.6 11.75 1.73 ;
 RECT 11.14 0.395 11.27 0.525 ;
 RECT 10.57 0.585 10.7 0.715 ;
 RECT 10.57 2.105 10.7 2.235 ;
 RECT 11.14 2.34 11.27 2.47 ;
 RECT 8.095 2.235 8.225 2.365 ;
 RECT 14.985 0.89 15.115 1.02 ;
 RECT 17.105 1.595 17.235 1.725 ;
 RECT 16.66 0.785 16.79 0.915 ;
 RECT 2.745 0.12 2.875 0.25 ;
 RECT 14.52 2.525 14.65 2.655 ;
 RECT 6.59 2.33 6.72 2.46 ;
 RECT 19.95 1.44 20.08 1.57 ;
 LAYER M1 ;
 RECT 3.645 0.55 3.785 1.275 ;
 RECT 3.645 1.415 3.785 1.71 ;
 RECT 2.5 1.275 3.785 1.415 ;
 RECT 13.65 1.17 13.99 1.51 ;
 RECT 6.175 1.21 6.405 1.245 ;
 RECT 6.175 1.385 6.405 1.42 ;
 RECT 6.175 1.245 7.36 1.385 ;
 RECT 6.95 0.55 7.09 1.245 ;
 RECT 7.13 1.385 7.36 1.625 ;
 RECT 17.1 0.92 17.24 1.785 ;
 RECT 17.015 0.78 17.265 0.92 ;
 RECT 16 0.36 16.14 0.5 ;
 RECT 14.495 0.22 16.14 0.36 ;
 RECT 17.405 0.435 17.545 0.5 ;
 RECT 17.405 0.64 17.545 1.61 ;
 RECT 16 0.5 17.545 0.64 ;
 RECT 1.265 2.37 2.46 2.51 ;
 RECT 1.265 0.53 1.405 2.37 ;
 RECT 2.32 2.23 5 2.37 ;
 RECT 4.86 2.465 6.145 2.51 ;
 RECT 4.86 2.37 6.78 2.465 ;
 RECT 6.005 2.325 6.78 2.37 ;
 RECT 1.925 0.6 2.33 0.735 ;
 RECT 1.925 0.735 2.065 1.765 ;
 RECT 3.205 0.41 3.345 0.46 ;
 RECT 3.965 0.41 4.105 1.475 ;
 RECT 1.925 0.595 3.345 0.6 ;
 RECT 2.13 0.46 3.345 0.595 ;
 RECT 3.205 0.27 4.105 0.41 ;
 RECT 15.72 0.64 15.86 0.78 ;
 RECT 15.72 0.92 15.86 1.455 ;
 RECT 15.72 0.78 16.855 0.92 ;
 RECT 15.615 0.5 15.86 0.64 ;
 RECT 12.855 1.095 12.995 1.835 ;
 RECT 13.18 0.925 13.41 0.955 ;
 RECT 12.855 0.955 13.41 1.095 ;
 RECT 13.18 1.095 13.41 1.135 ;
 RECT 16 1.33 16.14 2.52 ;
 RECT 14.44 2.52 16.14 2.66 ;
 RECT 18.44 0.64 18.58 1.925 ;
 RECT 16.65 1.33 16.79 1.925 ;
 RECT 18.375 0.5 18.625 0.64 ;
 RECT 16.65 1.925 18.58 2.065 ;
 RECT 16 1.19 16.79 1.33 ;
 RECT 13.49 1.845 13.63 2.45 ;
 RECT 12.455 2.385 12.595 2.45 ;
 RECT 12.455 2.59 12.595 2.65 ;
 RECT 12.455 2.45 13.63 2.59 ;
 RECT 14.345 0.585 14.485 1.705 ;
 RECT 13.49 1.705 14.485 1.845 ;
 RECT 14.345 1.845 14.485 2.265 ;
 RECT 5.185 1.765 7.78 1.8 ;
 RECT 5.185 1.665 5.61 1.765 ;
 RECT 5.255 0.545 5.395 1.665 ;
 RECT 5.185 1.8 8.92 1.805 ;
 RECT 8.78 0.365 8.92 1.8 ;
 RECT 9.34 0.365 9.48 1.205 ;
 RECT 5.47 1.805 8.92 1.905 ;
 RECT 8.78 0.225 9.48 0.365 ;
 RECT 7.64 1.905 8.92 1.94 ;
 RECT 9.34 1.205 9.965 1.345 ;
 RECT 10.18 0.385 10.32 2.21 ;
 RECT 10.845 0.385 10.985 0.75 ;
 RECT 10.18 0.245 10.985 0.385 ;
 RECT 11.3 0.89 11.44 1.165 ;
 RECT 10.845 0.75 11.44 0.89 ;
 RECT 19.525 0.435 19.665 1.07 ;
 RECT 19.525 1.21 19.665 1.64 ;
 RECT 18.725 1.07 19.665 1.21 ;
 RECT 5.815 0.55 5.955 1.475 ;
 RECT 5.75 1.475 6.02 1.615 ;
 RECT 9.9 1.775 10.04 2.435 ;
 RECT 9.34 1.635 10.04 1.775 ;
 RECT 10.855 2.135 10.995 2.435 ;
 RECT 9.9 2.435 10.995 2.575 ;
 RECT 9.34 1.775 9.48 2.52 ;
 RECT 9.11 2.52 9.48 2.66 ;
 RECT 11.895 1.86 12.035 1.995 ;
 RECT 10.855 1.995 12.035 2.135 ;
 RECT 12.57 2.045 13.235 2.185 ;
 RECT 12.57 1.86 12.71 2.045 ;
 RECT 12.57 0.77 12.71 1.72 ;
 RECT 12.57 0.63 13.235 0.77 ;
 RECT 11.895 1.72 12.71 1.86 ;
 RECT 18.765 0.36 18.905 0.79 ;
 RECT 17.965 0.36 18.105 1.41 ;
 RECT 17.965 0.22 18.905 0.36 ;
 RECT 17.9 1.41 18.17 1.55 ;
 RECT 18.765 0.79 19.385 0.93 ;
 RECT 3.01 2.08 7.445 2.085 ;
 RECT 5.14 2.085 7.445 2.09 ;
 RECT 5.43 2.045 7.445 2.08 ;
 RECT 3.01 1.945 5.28 2.08 ;
 RECT 5.14 2.185 5.66 2.22 ;
 RECT 4.275 0.835 4.415 1.945 ;
 RECT 3.01 1.715 3.15 1.945 ;
 RECT 2.94 1.575 3.215 1.715 ;
 RECT 8.09 2.23 8.23 2.435 ;
 RECT 5.14 2.09 9.2 2.185 ;
 RECT 7.305 2.185 9.2 2.23 ;
 RECT 9.06 0.505 9.2 2.09 ;
 RECT 6.67 0.38 6.81 0.93 ;
 RECT 6.67 0.24 7.39 0.38 ;
 RECT 7.25 0.38 7.39 0.925 ;
 RECT 6.105 0.93 6.81 1.07 ;
 RECT 4.775 0.375 4.915 1.26 ;
 RECT 6.105 0.375 6.245 0.93 ;
 RECT 4.605 1.26 4.915 1.4 ;
 RECT 4.605 1.4 4.745 1.77 ;
 RECT 4.775 0.235 6.245 0.375 ;
 RECT 7.835 1.065 7.975 1.48 ;
 RECT 7.835 0.515 8.06 0.785 ;
 RECT 7.835 0.785 7.975 0.925 ;
 RECT 7.785 1.48 8.025 1.62 ;
 RECT 7.25 0.925 7.975 1.065 ;
 END
END RDFFNARX1

MACRO RDFFNARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 23.04 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.06 0.82 3.505 1.115 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.82 1.12 1.12 1.395 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END RSTB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.18 1.14 8.64 1.42 ;
 END
 ANTENNAGATEAREA 0.05 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.35 1.14 11.705 1.48 ;
 RECT 11.35 1.48 11.49 1.855 ;
 RECT 11.35 0.525 11.49 1.14 ;
 END
 ANTENNADIFFAREA 0.748 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.4 1.465 12.54 1.855 ;
 RECT 12.4 1.12 12.94 1.465 ;
 RECT 12.4 0.48 12.54 1.12 ;
 END
 ANTENNADIFFAREA 0.626 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 23.04 2.96 ;
 RECT 6.325 2.615 6.56 2.8 ;
 RECT 10.74 2.275 11.01 2.415 ;
 RECT 12.815 2.275 13.085 2.415 ;
 RECT 8.375 2.37 8.645 2.51 ;
 RECT 2.675 2.51 2.945 2.65 ;
 RECT 11.855 2.275 12.125 2.415 ;
 RECT 4.37 2.51 4.6 2.65 ;
 RECT 0.265 1.64 0.425 2.8 ;
 RECT 0.67 1.855 0.81 2.8 ;
 RECT 13.25 2 13.39 2.8 ;
 RECT 14.94 2.025 15.08 2.8 ;
 RECT 9.62 1.94 9.76 2.8 ;
 RECT 10.805 2.415 10.945 2.8 ;
 RECT 12.88 2.415 13.02 2.8 ;
 RECT 8.44 2.51 8.58 2.8 ;
 RECT 2.74 2.65 2.88 2.8 ;
 RECT 11.92 2.415 12.06 2.8 ;
 RECT 4.415 2.65 4.555 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 23.04 0.08 ;
 RECT 8.37 0.565 8.64 0.705 ;
 RECT 17.34 0.22 17.59 0.36 ;
 RECT 4.38 0.555 4.63 0.695 ;
 RECT 11.92 0.08 12.06 0.575 ;
 RECT 20.105 0.08 20.245 0.65 ;
 RECT 13.3 0.08 13.44 0.865 ;
 RECT 14.94 0.08 15.08 0.815 ;
 RECT 6.39 0.08 6.53 0.78 ;
 RECT 0.265 0.08 0.425 0.84 ;
 RECT 9.62 0.08 9.76 0.785 ;
 RECT 0.705 0.08 0.845 0.79 ;
 RECT 1.645 0.08 1.785 0.8 ;
 RECT 2.74 0.08 2.88 0.32 ;
 RECT 10.79 0.08 10.93 0.575 ;
 RECT 12.87 0.08 13.01 0.575 ;
 RECT 7.53 0.08 7.67 0.78 ;
 RECT 8.435 0.08 8.575 0.565 ;
 RECT 17.385 0.08 17.525 0.22 ;
 RECT 4.445 0.08 4.585 0.555 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 20.865 1.4 21.19 1.765 ;
 RECT 17.385 2.225 21.125 2.385 ;
 RECT 17.34 1.47 17.57 1.61 ;
 RECT 20.06 1.395 20.2 2.225 ;
 RECT 20.975 1.765 21.115 2.225 ;
 RECT 17.385 1.61 17.525 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 15.86 0.82 16.18 1.1 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 11.605 1.04 11.705 1.22 ;
 RECT 11.05 0.1 11.15 0.94 ;
 RECT 9.91 0.365 10.01 1.16 ;
 RECT 9.91 1.39 10.01 2.47 ;
 RECT 11.605 1.32 11.705 2.75 ;
 RECT 11.06 1.32 11.16 2.745 ;
 RECT 11.05 0.94 11.705 1.04 ;
 RECT 0.975 0.35 1.075 1.145 ;
 RECT 0.845 1.145 1.075 1.375 ;
 RECT 0.975 1.375 1.075 2.485 ;
 RECT 3.395 0.38 3.495 0.865 ;
 RECT 3.395 1.095 3.495 2.36 ;
 RECT 3.275 0.865 3.505 1.095 ;
 RECT 3.085 1.76 3.185 2.34 ;
 RECT 2.965 1.53 3.195 1.76 ;
 RECT 8.175 0.33 8.275 2.185 ;
 RECT 8.045 2.185 8.275 2.415 ;
 RECT 19.755 0.275 19.855 1.025 ;
 RECT 19.755 1.255 19.855 1.86 ;
 RECT 19.755 1.025 20.035 1.255 ;
 RECT 6.65 0.37 6.75 2.28 ;
 RECT 6.54 2.28 6.77 2.51 ;
 RECT 5.515 1.445 5.615 2.035 ;
 RECT 5.43 2.035 5.66 2.265 ;
 RECT 4.69 1.75 4.79 2.62 ;
 RECT 4.22 1.73 4.32 2.34 ;
 RECT 4.56 1.53 4.79 1.63 ;
 RECT 4.56 1.73 4.79 1.75 ;
 RECT 4.22 1.63 4.79 1.73 ;
 RECT 8.7 0.33 8.8 1.145 ;
 RECT 8.7 1.38 8.8 2.235 ;
 RECT 8.455 1.145 8.8 1.38 ;
 RECT 2.995 0.1 5.69 0.2 ;
 RECT 5.39 0.2 5.69 0.42 ;
 RECT 5.59 0.42 5.69 0.95 ;
 RECT 2.995 0.2 3.095 0.97 ;
 RECT 13.585 0.385 13.685 2.405 ;
 RECT 13.485 2.405 13.715 2.635 ;
 RECT 13.895 1.835 13.995 2.425 ;
 RECT 13.885 1.605 14.115 1.835 ;
 RECT 6.12 0.37 6.22 1.21 ;
 RECT 6.12 1.21 6.405 1.42 ;
 RECT 6.12 1.42 6.22 2.16 ;
 RECT 2.18 1.095 2.28 2.325 ;
 RECT 1.91 0.38 2.01 0.995 ;
 RECT 2.05 2.325 2.28 2.555 ;
 RECT 1.91 0.995 2.28 1.095 ;
 RECT 20.36 0.27 20.46 0.745 ;
 RECT 20.36 0.975 20.46 1.855 ;
 RECT 20.215 0.745 20.46 0.975 ;
 RECT 18.095 0.865 18.82 0.965 ;
 RECT 18.095 0.735 18.325 0.865 ;
 RECT 18.72 0.275 18.82 0.865 ;
 RECT 3.92 1.34 4.15 1.45 ;
 RECT 3.92 0.38 4.02 1.24 ;
 RECT 3.92 1.45 4.02 2.345 ;
 RECT 5.015 0.38 5.115 1.24 ;
 RECT 3.92 1.24 5.115 1.34 ;
 RECT 5.015 1.34 5.115 2.62 ;
 RECT 14.425 2.605 15.775 2.695 ;
 RECT 14.425 1.425 14.525 2.605 ;
 RECT 14.43 2.695 15.775 2.705 ;
 RECT 13.89 0.385 13.99 1.325 ;
 RECT 15.545 2.475 15.775 2.605 ;
 RECT 13.89 1.325 14.525 1.425 ;
 RECT 2.5 0.38 2.6 1.23 ;
 RECT 2.5 1.46 2.6 2.34 ;
 RECT 2.5 1.23 2.73 1.46 ;
 RECT 6.95 1.06 7.05 2.68 ;
 RECT 7.26 0.37 7.36 0.96 ;
 RECT 9.13 2.475 9.36 2.68 ;
 RECT 6.95 0.96 7.36 1.06 ;
 RECT 6.95 2.68 9.36 2.78 ;
 RECT 17.67 0.965 17.77 1.145 ;
 RECT 19.28 0.275 19.38 0.865 ;
 RECT 17.67 1.145 19.1 1.245 ;
 RECT 19 0.965 19.1 1.145 ;
 RECT 18.81 1.245 18.91 1.86 ;
 RECT 17.67 0.735 17.9 0.965 ;
 RECT 19 0.865 19.38 0.965 ;
 RECT 12.655 0.105 15.85 0.205 ;
 RECT 14.38 0.205 14.48 0.925 ;
 RECT 12.655 0.205 12.755 0.9 ;
 RECT 12.175 0.105 12.275 0.87 ;
 RECT 12.04 0.87 12.275 0.9 ;
 RECT 12.04 0.9 12.755 1 ;
 RECT 15.62 0.205 15.85 0.4 ;
 RECT 12.175 1.085 12.275 1.2 ;
 RECT 12.175 1.2 12.765 1.3 ;
 RECT 12.175 1.3 12.275 2.755 ;
 RECT 12.665 1.3 12.765 2.745 ;
 RECT 12.04 1 12.275 1.085 ;
 RECT 14.255 0.925 14.485 1.135 ;
 RECT 14.725 1.27 15.3 1.37 ;
 RECT 14.725 1.215 15 1.27 ;
 RECT 14.725 0.385 14.825 1.215 ;
 RECT 14.725 1.37 15 1.425 ;
 RECT 14.725 1.425 14.825 2.425 ;
 RECT 15.2 1.045 15.3 1.27 ;
 RECT 15.2 1.37 15.3 2.425 ;
 RECT 17.09 0.145 17.19 0.945 ;
 RECT 15.2 0.945 17.19 1.045 ;
 RECT 17.09 1.045 17.19 1.76 ;
 RECT 19.28 1.145 19.38 2.09 ;
 RECT 18.245 1.86 18.345 2.09 ;
 RECT 18.115 1.545 18.345 1.76 ;
 RECT 15.935 0.84 16.165 0.945 ;
 RECT 15.935 1.045 16.165 1.07 ;
 RECT 15.2 0.385 15.3 0.945 ;
 RECT 18.245 2.09 19.38 2.19 ;
 RECT 17.09 1.76 18.345 1.86 ;
 RECT 4.225 0.38 4.325 0.84 ;
 RECT 4.225 0.87 4.8 0.97 ;
 RECT 4.7 0.38 4.8 0.87 ;
 RECT 4.225 0.84 4.47 0.87 ;
 RECT 4.225 0.97 4.47 1.06 ;
 RECT 9.715 1.16 10.01 1.22 ;
 RECT 9.715 1.22 11.705 1.32 ;
 RECT 9.715 1.32 10.01 1.39 ;
 RECT 11.605 0.105 11.705 0.94 ;
 LAYER CO ;
 RECT 3.65 0.6 3.78 0.73 ;
 RECT 1.65 0.6 1.78 0.73 ;
 RECT 15.67 0.225 15.8 0.355 ;
 RECT 17.39 1.475 17.52 1.605 ;
 RECT 16.785 1.255 16.915 1.385 ;
 RECT 16.74 0.505 16.87 0.635 ;
 RECT 15.595 2.525 15.725 2.655 ;
 RECT 13.535 2.455 13.665 2.585 ;
 RECT 13.935 1.655 14.065 1.785 ;
 RECT 15.425 0.635 15.555 0.765 ;
 RECT 14.945 0.635 15.075 0.765 ;
 RECT 14.945 2.075 15.075 2.205 ;
 RECT 14.82 1.255 14.95 1.385 ;
 RECT 14.305 0.965 14.435 1.095 ;
 RECT 5.26 1.67 5.39 1.8 ;
 RECT 2.745 2.515 2.875 2.645 ;
 RECT 4.42 2.515 4.55 2.645 ;
 RECT 3.65 1.52 3.78 1.65 ;
 RECT 7.18 1.49 7.31 1.62 ;
 RECT 7.535 0.6 7.665 0.73 ;
 RECT 6.955 0.6 7.085 0.73 ;
 RECT 6.395 0.6 6.525 0.73 ;
 RECT 5.82 0.6 5.95 0.73 ;
 RECT 5.82 1.48 5.95 1.61 ;
 RECT 5.26 0.6 5.39 0.73 ;
 RECT 14.13 2.05 14.26 2.18 ;
 RECT 14.13 0.635 14.26 0.765 ;
 RECT 13.305 0.635 13.435 0.765 ;
 RECT 13.255 2.06 13.385 2.19 ;
 RECT 15.425 2.065 15.555 2.195 ;
 RECT 11.355 1.675 11.485 1.805 ;
 RECT 18.145 0.785 18.275 0.915 ;
 RECT 20.265 0.795 20.395 0.925 ;
 RECT 19.855 1.075 19.985 1.205 ;
 RECT 20.59 0.505 20.72 0.635 ;
 RECT 20.59 1.44 20.72 1.57 ;
 RECT 20.11 0.47 20.24 0.6 ;
 RECT 20.065 1.455 20.195 1.585 ;
 RECT 19.505 1.435 19.635 1.565 ;
 RECT 5.48 2.085 5.61 2.215 ;
 RECT 0.28 0.36 0.41 0.49 ;
 RECT 0.28 0.62 0.41 0.75 ;
 RECT 0.28 1.71 0.41 1.84 ;
 RECT 0.28 1.97 0.41 2.1 ;
 RECT 0.28 2.23 0.41 2.36 ;
 RECT 17.39 0.225 17.52 0.355 ;
 RECT 5.44 0.24 5.57 0.37 ;
 RECT 4.61 1.57 4.74 1.7 ;
 RECT 4.28 0.89 4.41 1.02 ;
 RECT 3.97 1.28 4.1 1.41 ;
 RECT 3.015 1.58 3.145 1.71 ;
 RECT 3.325 0.915 3.455 1.045 ;
 RECT 2.55 1.28 2.68 1.41 ;
 RECT 2.1 2.375 2.23 2.505 ;
 RECT 9.065 0.57 9.195 0.7 ;
 RECT 9.065 1.845 9.195 1.975 ;
 RECT 8.44 0.57 8.57 0.7 ;
 RECT 7.925 0.57 8.055 0.7 ;
 RECT 7.86 1.48 7.99 1.61 ;
 RECT 8.445 2.375 8.575 2.505 ;
 RECT 6.38 2.63 6.51 2.76 ;
 RECT 1.93 1.585 2.06 1.715 ;
 RECT 2.13 0.6 2.26 0.73 ;
 RECT 1.27 1.875 1.4 2.005 ;
 RECT 1.27 0.58 1.4 0.71 ;
 RECT 0.71 0.59 0.84 0.72 ;
 RECT 0.675 1.905 0.805 2.035 ;
 RECT 9.18 2.525 9.31 2.655 ;
 RECT 12.09 0.915 12.22 1.045 ;
 RECT 12.405 1.675 12.535 1.805 ;
 RECT 11.925 0.395 12.055 0.525 ;
 RECT 11.355 0.585 11.485 0.715 ;
 RECT 11.925 2.28 12.055 2.41 ;
 RECT 12.875 0.395 13.005 0.525 ;
 RECT 12.885 2.28 13.015 2.41 ;
 RECT 10.795 0.395 10.925 0.525 ;
 RECT 0.885 1.195 1.015 1.325 ;
 RECT 4.45 0.555 4.58 0.685 ;
 RECT 10.81 2.28 10.94 2.41 ;
 RECT 8.095 2.235 8.225 2.365 ;
 RECT 15.985 0.89 16.115 1.02 ;
 RECT 18.165 1.595 18.295 1.725 ;
 RECT 17.72 0.785 17.85 0.915 ;
 RECT 2.745 0.12 2.875 0.25 ;
 RECT 21.01 1.44 21.14 1.57 ;
 RECT 6.225 1.25 6.355 1.38 ;
 RECT 19.505 0.505 19.635 0.635 ;
 RECT 19.03 1.415 19.16 1.545 ;
 RECT 19.03 0.505 19.16 0.635 ;
 RECT 18.47 1.415 18.6 1.545 ;
 RECT 18.47 0.505 18.6 0.635 ;
 RECT 12.405 0.555 12.535 0.685 ;
 RECT 9.625 2.01 9.755 2.14 ;
 RECT 9.765 1.21 9.895 1.34 ;
 RECT 9.625 0.605 9.755 0.735 ;
 RECT 10.185 2.025 10.315 2.155 ;
 RECT 10.185 0.605 10.315 0.735 ;
 RECT 8.505 1.2 8.635 1.33 ;
 RECT 6.59 2.33 6.72 2.46 ;
 LAYER M1 ;
 RECT 14.725 1.17 15.065 1.51 ;
 RECT 7.25 0.38 7.39 0.925 ;
 RECT 6.67 0.38 6.81 0.93 ;
 RECT 6.67 0.24 7.39 0.38 ;
 RECT 6.105 0.93 6.81 1.07 ;
 RECT 4.775 0.375 4.915 1.26 ;
 RECT 6.105 0.375 6.245 0.93 ;
 RECT 4.605 1.26 4.915 1.4 ;
 RECT 4.605 1.4 4.745 1.77 ;
 RECT 4.775 0.235 6.245 0.375 ;
 RECT 7.855 0.495 8.06 0.925 ;
 RECT 7.855 1.065 7.995 1.475 ;
 RECT 7.25 0.925 8.06 0.975 ;
 RECT 7.25 0.975 7.995 1.065 ;
 RECT 7.81 1.475 8.04 1.615 ;
 RECT 19.025 0.36 19.165 1.41 ;
 RECT 19.825 0.36 19.965 0.79 ;
 RECT 18.96 1.41 19.23 1.55 ;
 RECT 19.025 0.22 19.965 0.36 ;
 RECT 19.825 0.79 20.445 0.93 ;
 RECT 3.645 0.55 3.785 1.275 ;
 RECT 2.5 1.275 3.785 1.415 ;
 RECT 3.645 1.415 3.785 1.71 ;
 RECT 18.16 0.92 18.3 1.785 ;
 RECT 18.075 0.78 18.325 0.92 ;
 RECT 1.925 0.6 2.33 0.735 ;
 RECT 1.925 0.735 2.065 1.765 ;
 RECT 3.205 0.41 3.345 0.46 ;
 RECT 1.925 0.595 3.345 0.6 ;
 RECT 2.13 0.46 3.345 0.595 ;
 RECT 3.965 0.41 4.105 1.475 ;
 RECT 3.205 0.27 4.105 0.41 ;
 RECT 5.815 0.55 5.955 1.475 ;
 RECT 5.75 1.475 6.02 1.615 ;
 RECT 14.565 1.845 14.705 2.45 ;
 RECT 13.53 2.385 13.67 2.45 ;
 RECT 13.53 2.59 13.67 2.65 ;
 RECT 13.53 2.45 14.705 2.59 ;
 RECT 15.42 0.585 15.56 1.705 ;
 RECT 14.565 1.705 15.56 1.845 ;
 RECT 15.42 1.845 15.56 2.265 ;
 RECT 13.93 1.095 14.07 1.835 ;
 RECT 14.255 0.925 14.485 0.955 ;
 RECT 14.255 1.095 14.485 1.135 ;
 RECT 13.93 0.955 14.485 1.095 ;
 RECT 20.585 0.435 20.725 1.07 ;
 RECT 19.785 1.07 20.725 1.21 ;
 RECT 20.585 1.21 20.725 1.64 ;
 RECT 1.265 2.37 2.46 2.51 ;
 RECT 1.265 0.53 1.405 2.37 ;
 RECT 2.32 2.23 5 2.37 ;
 RECT 4.86 2.465 6.145 2.51 ;
 RECT 4.86 2.37 6.78 2.465 ;
 RECT 6.005 2.325 6.78 2.37 ;
 RECT 16.78 0.64 16.92 0.78 ;
 RECT 16.78 0.92 16.92 1.455 ;
 RECT 16.675 0.5 16.92 0.64 ;
 RECT 16.78 0.78 17.915 0.92 ;
 RECT 15.515 2.52 17.2 2.65 ;
 RECT 15.515 2.65 17.19 2.66 ;
 RECT 17.06 1.33 17.2 2.52 ;
 RECT 17.71 1.33 17.85 1.925 ;
 RECT 19.5 0.64 19.64 1.925 ;
 RECT 17.06 1.19 17.85 1.33 ;
 RECT 19.435 0.5 19.685 0.64 ;
 RECT 17.71 1.925 19.64 2.065 ;
 RECT 5.185 1.765 7.78 1.8 ;
 RECT 5.185 1.665 5.61 1.765 ;
 RECT 5.255 0.545 5.395 1.665 ;
 RECT 5.185 1.8 8.92 1.805 ;
 RECT 8.78 0.365 8.92 1.8 ;
 RECT 9.34 0.365 9.48 1.205 ;
 RECT 5.47 1.805 8.92 1.905 ;
 RECT 8.78 0.225 9.48 0.365 ;
 RECT 7.64 1.905 8.92 1.94 ;
 RECT 9.34 1.205 9.965 1.345 ;
 RECT 9.9 1.775 10.04 2.435 ;
 RECT 10.46 2.135 10.6 2.435 ;
 RECT 9.34 1.635 10.04 1.775 ;
 RECT 9.9 2.435 10.6 2.575 ;
 RECT 9.34 1.775 9.48 2.52 ;
 RECT 9.11 2.52 9.48 2.66 ;
 RECT 12.97 1.86 13.11 1.995 ;
 RECT 10.46 1.995 13.11 2.135 ;
 RECT 13.645 2.045 14.31 2.185 ;
 RECT 13.645 1.86 13.785 2.045 ;
 RECT 13.645 0.63 14.31 0.77 ;
 RECT 13.645 0.77 13.785 1.72 ;
 RECT 12.97 1.72 13.785 1.86 ;
 RECT 5.14 2.085 7.445 2.09 ;
 RECT 3.01 2.08 7.445 2.085 ;
 RECT 5.43 2.045 7.445 2.08 ;
 RECT 3.01 1.945 5.28 2.08 ;
 RECT 5.14 2.185 5.66 2.22 ;
 RECT 4.275 0.835 4.415 1.945 ;
 RECT 3.01 1.715 3.15 1.945 ;
 RECT 2.94 1.575 3.215 1.715 ;
 RECT 8.09 2.23 8.23 2.435 ;
 RECT 5.14 2.09 9.2 2.185 ;
 RECT 7.305 2.185 9.2 2.23 ;
 RECT 9.06 0.52 9.2 2.09 ;
 RECT 11.07 0.385 11.21 0.79 ;
 RECT 10.18 0.79 11.21 0.93 ;
 RECT 10.18 0.55 10.32 0.79 ;
 RECT 10.18 0.93 10.32 2.21 ;
 RECT 11.63 0.385 11.77 0.75 ;
 RECT 11.07 0.245 11.77 0.385 ;
 RECT 11.63 0.755 12.225 0.89 ;
 RECT 11.63 0.75 12.145 0.755 ;
 RECT 12.085 0.89 12.225 1.095 ;
 RECT 7.13 1.385 7.36 1.625 ;
 RECT 6.175 1.245 7.36 1.385 ;
 RECT 6.95 0.55 7.09 1.245 ;
 RECT 6.175 1.21 6.405 1.245 ;
 RECT 6.175 1.385 6.405 1.42 ;
 RECT 17.06 0.36 17.2 0.5 ;
 RECT 15.57 0.22 17.2 0.36 ;
 RECT 17.06 0.5 18.605 0.64 ;
 RECT 18.465 0.435 18.605 0.5 ;
 RECT 18.465 0.64 18.605 1.61 ;
 END
END RDFFNARX2

MACRO RSDFFARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 25.28 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.135 1.13 1.655 1.47 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.835 0.875 2.08 1.11 ;
 RECT 2.025 1.5 2.385 1.805 ;
 RECT 1.89 1.46 2.385 1.5 ;
 RECT 1.89 1.36 2.175 1.46 ;
 RECT 1.89 1.11 2.03 1.36 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.615 2.385 2.2 2.5 ;
 RECT 1.46 2.25 2.2 2.385 ;
 RECT 1.46 2.09 1.78 2.25 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.695 1.44 4.11 1.745 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END RSTB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.375 0.815 11.84 1.12 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.765 1.5 13.905 2.295 ;
 RECT 13.765 1.09 14.26 1.5 ;
 RECT 13.765 0.525 13.905 1.09 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.78 1.12 15.18 1.465 ;
 RECT 14.815 1.465 14.955 1.79 ;
 RECT 14.815 0.48 14.955 1.12 ;
 END
 ANTENNADIFFAREA 0.471 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 25.28 2.96 ;
 RECT 9.525 2.615 9.76 2.8 ;
 RECT 2.82 1.97 3.2 2.11 ;
 RECT 5.875 2.51 6.145 2.65 ;
 RECT 7.57 2.51 7.8 2.65 ;
 RECT 11.625 2.37 11.895 2.51 ;
 RECT 0.39 1.64 0.55 2.8 ;
 RECT 1.305 2.535 1.445 2.8 ;
 RECT 3.69 1.965 3.83 2.8 ;
 RECT 12.82 1.94 12.96 2.8 ;
 RECT 17.065 2.025 17.205 2.8 ;
 RECT 15.375 2 15.515 2.8 ;
 RECT 14.335 2.275 14.475 2.8 ;
 RECT 3.06 2.11 3.2 2.8 ;
 RECT 5.94 2.65 6.08 2.8 ;
 RECT 7.615 2.65 7.755 2.8 ;
 RECT 11.69 2.51 11.83 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 25.28 0.08 ;
 RECT 2.8 0.59 3.2 0.73 ;
 RECT 7.58 0.555 7.83 0.695 ;
 RECT 11.57 0.49 11.84 0.63 ;
 RECT 20.025 0.22 20.275 0.36 ;
 RECT 1.305 0.08 1.445 0.31 ;
 RECT 0.39 0.08 0.55 0.84 ;
 RECT 5.94 0.08 6.08 0.32 ;
 RECT 4.845 0.08 4.985 0.8 ;
 RECT 3.725 0.08 3.865 0.79 ;
 RECT 9.59 0.08 9.73 0.78 ;
 RECT 10.73 0.08 10.87 0.78 ;
 RECT 12.82 0.08 12.96 0.785 ;
 RECT 15.425 0.08 15.565 0.865 ;
 RECT 17.065 0.08 17.205 0.815 ;
 RECT 14.335 0.08 14.475 0.575 ;
 RECT 22.79 0.08 22.93 0.65 ;
 RECT 3.06 0.08 3.2 0.59 ;
 RECT 7.645 0.08 7.785 0.555 ;
 RECT 11.64 0.63 11.78 0.645 ;
 RECT 11.64 0.08 11.78 0.49 ;
 RECT 20.07 0.08 20.21 0.22 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 23.645 1.4 24.145 1.765 ;
 RECT 20.025 1.47 20.255 1.61 ;
 RECT 20.075 2.31 23.81 2.385 ;
 RECT 20.07 2.225 23.81 2.31 ;
 RECT 20.07 1.61 20.21 2.225 ;
 RECT 22.745 1.395 22.885 2.225 ;
 RECT 23.66 1.765 23.8 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.075 0.81 18.575 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 20.355 0.965 20.455 1.145 ;
 RECT 20.355 1.145 21.785 1.245 ;
 RECT 21.685 0.965 21.785 1.145 ;
 RECT 21.495 1.245 21.595 1.86 ;
 RECT 21.965 0.275 22.065 0.865 ;
 RECT 20.355 0.735 20.585 0.965 ;
 RECT 21.685 0.865 22.065 0.965 ;
 RECT 20.78 0.865 21.505 0.965 ;
 RECT 20.78 0.735 21.01 0.865 ;
 RECT 21.405 0.275 21.505 0.865 ;
 RECT 1.865 1.385 1.965 2.295 ;
 RECT 2.335 0.365 2.435 1.285 ;
 RECT 1.865 2.525 1.965 2.53 ;
 RECT 1.865 2.295 2.145 2.525 ;
 RECT 1.865 1.285 2.435 1.385 ;
 RECT 5.38 1.095 5.48 2.325 ;
 RECT 5.11 0.38 5.21 0.995 ;
 RECT 5.25 2.325 5.48 2.555 ;
 RECT 5.11 0.995 5.48 1.095 ;
 RECT 3.995 0.35 4.095 1.465 ;
 RECT 3.865 1.465 4.095 1.695 ;
 RECT 3.995 1.695 4.095 2.485 ;
 RECT 2.64 0.43 2.74 2.385 ;
 RECT 2.615 0.22 2.845 0.43 ;
 RECT 12.915 1.16 13.21 1.22 ;
 RECT 13.11 0.365 13.21 1.16 ;
 RECT 12.915 1.32 13.21 1.39 ;
 RECT 13.11 1.39 13.21 2.47 ;
 RECT 14.02 0.105 14.12 1.22 ;
 RECT 14.02 1.32 14.12 2.75 ;
 RECT 12.915 1.22 14.12 1.32 ;
 RECT 11.375 0.25 11.475 0.865 ;
 RECT 11.375 0.865 11.665 1.08 ;
 RECT 11.375 1.08 11.475 2.235 ;
 RECT 9.85 0.37 9.95 2.28 ;
 RECT 9.74 2.28 9.97 2.51 ;
 RECT 8.715 1.445 8.815 2.035 ;
 RECT 8.63 2.035 8.86 2.265 ;
 RECT 7.89 1.75 7.99 2.44 ;
 RECT 7.42 1.73 7.52 2.34 ;
 RECT 7.76 1.53 7.99 1.63 ;
 RECT 7.76 1.73 7.99 1.75 ;
 RECT 7.42 1.63 7.99 1.73 ;
 RECT 9.32 0.37 9.42 1.21 ;
 RECT 9.32 1.42 9.42 2.16 ;
 RECT 9.32 1.21 9.605 1.42 ;
 RECT 7.425 0.87 8 0.97 ;
 RECT 7.9 0.38 8 0.87 ;
 RECT 7.425 0.84 7.67 0.87 ;
 RECT 7.425 0.97 7.67 1.06 ;
 RECT 7.425 0.38 7.525 0.84 ;
 RECT 1.09 0.345 1.19 1.23 ;
 RECT 1.09 1.33 1.19 2.385 ;
 RECT 1.09 1.23 1.66 1.33 ;
 RECT 1.43 1.165 1.66 1.23 ;
 RECT 1.43 1.33 1.66 1.395 ;
 RECT 1.56 0.345 1.66 1.165 ;
 RECT 1.56 1.395 1.66 2.385 ;
 RECT 6.285 1.76 6.385 2.34 ;
 RECT 6.165 1.53 6.395 1.76 ;
 RECT 16.85 0.385 16.95 1.215 ;
 RECT 16.85 1.215 17.125 1.27 ;
 RECT 16.85 1.425 16.95 2.425 ;
 RECT 16.85 1.37 17.125 1.425 ;
 RECT 17.325 1.045 17.425 1.27 ;
 RECT 17.325 1.37 17.425 2.425 ;
 RECT 16.85 1.27 17.425 1.37 ;
 RECT 19.775 0.145 19.875 0.945 ;
 RECT 19.775 1.045 19.875 1.76 ;
 RECT 21.965 1.145 22.065 2.09 ;
 RECT 20.93 1.86 21.03 2.09 ;
 RECT 18.285 0.84 18.515 0.945 ;
 RECT 18.285 1.045 18.515 1.07 ;
 RECT 17.325 0.385 17.425 0.945 ;
 RECT 17.325 0.945 19.875 1.045 ;
 RECT 20.8 1.545 21.03 1.76 ;
 RECT 20.93 2.09 22.065 2.19 ;
 RECT 19.775 1.76 21.03 1.86 ;
 RECT 14.6 0.105 17.975 0.205 ;
 RECT 14.6 0.205 14.7 0.87 ;
 RECT 16.505 0.205 16.605 0.925 ;
 RECT 14.6 1.085 14.7 2.755 ;
 RECT 14.455 0.87 14.7 1.085 ;
 RECT 17.745 0.205 17.975 0.4 ;
 RECT 16.38 0.925 16.61 1.135 ;
 RECT 8.59 0.2 8.89 0.42 ;
 RECT 8.79 0.42 8.89 0.95 ;
 RECT 6.195 0.2 6.295 0.97 ;
 RECT 6.195 0.1 8.89 0.2 ;
 RECT 11.955 0.26 12.055 1.27 ;
 RECT 11.955 1.49 12.055 2.235 ;
 RECT 11.655 1.27 12.055 1.49 ;
 RECT 2.335 1.795 2.435 2.385 ;
 RECT 2.145 1.565 2.435 1.795 ;
 RECT 16.55 2.605 17.9 2.695 ;
 RECT 17.67 2.475 17.9 2.605 ;
 RECT 16.55 1.425 16.65 2.605 ;
 RECT 16.015 0.385 16.115 1.325 ;
 RECT 16.555 2.695 17.9 2.705 ;
 RECT 16.015 1.325 16.65 1.425 ;
 RECT 10.15 1.06 10.25 2.68 ;
 RECT 12.33 2.475 12.56 2.68 ;
 RECT 10.46 0.37 10.56 0.96 ;
 RECT 10.15 2.68 12.56 2.78 ;
 RECT 10.15 0.96 10.56 1.06 ;
 RECT 7.12 0.38 7.22 1.24 ;
 RECT 7.12 1.45 7.22 2.345 ;
 RECT 8.215 0.38 8.315 1.24 ;
 RECT 7.12 1.24 8.315 1.34 ;
 RECT 8.215 1.34 8.315 2.435 ;
 RECT 7.12 1.34 7.35 1.45 ;
 RECT 6.595 0.38 6.695 0.945 ;
 RECT 6.595 1.175 6.695 2.36 ;
 RECT 6.475 0.945 6.705 1.175 ;
 RECT 5.7 0.38 5.8 1.23 ;
 RECT 5.7 1.46 5.8 2.34 ;
 RECT 5.7 1.23 5.93 1.46 ;
 RECT 15.71 0.385 15.81 2.405 ;
 RECT 15.61 2.405 15.84 2.635 ;
 RECT 3.12 0.35 3.22 1.205 ;
 RECT 3.12 1.415 3.22 2.395 ;
 RECT 2.97 1.205 3.22 1.415 ;
 RECT 23.045 0.27 23.145 0.745 ;
 RECT 23.045 0.975 23.145 1.855 ;
 RECT 22.9 0.745 23.145 0.975 ;
 RECT 22.44 0.275 22.54 1.025 ;
 RECT 22.44 1.255 22.54 1.86 ;
 RECT 22.44 1.025 22.72 1.255 ;
 RECT 1.865 0.335 1.965 0.875 ;
 RECT 1.84 0.875 2.07 1.105 ;
 RECT 16.02 1.835 16.12 2.425 ;
 RECT 16.01 1.605 16.24 1.835 ;
 LAYER CO ;
 RECT 17.72 2.525 17.85 2.655 ;
 RECT 15.66 2.455 15.79 2.585 ;
 RECT 16.06 1.655 16.19 1.785 ;
 RECT 17.55 0.635 17.68 0.765 ;
 RECT 17.07 0.635 17.2 0.765 ;
 RECT 17.07 2.075 17.2 2.205 ;
 RECT 16.255 2.05 16.385 2.18 ;
 RECT 16.255 0.635 16.385 0.765 ;
 RECT 15.43 0.635 15.56 0.765 ;
 RECT 20.83 0.785 20.96 0.915 ;
 RECT 22.95 0.795 23.08 0.925 ;
 RECT 22.54 1.075 22.67 1.205 ;
 RECT 20.85 1.595 20.98 1.725 ;
 RECT 23.275 0.505 23.405 0.635 ;
 RECT 23.275 1.44 23.405 1.57 ;
 RECT 22.795 0.47 22.925 0.6 ;
 RECT 20.405 0.785 20.535 0.915 ;
 RECT 6.525 0.995 6.655 1.125 ;
 RECT 5.75 1.28 5.88 1.41 ;
 RECT 5.3 2.375 5.43 2.505 ;
 RECT 1.965 2.345 2.095 2.475 ;
 RECT 1.89 0.925 2.02 1.055 ;
 RECT 1.89 0.925 2.02 1.055 ;
 RECT 1.48 1.215 1.61 1.345 ;
 RECT 2.195 1.615 2.325 1.745 ;
 RECT 12.265 0.57 12.395 0.7 ;
 RECT 4.85 0.6 4.98 0.73 ;
 RECT 3.345 1.975 3.475 2.105 ;
 RECT 11.125 1.48 11.255 1.61 ;
 RECT 3.345 0.595 3.475 0.725 ;
 RECT 2.87 0.595 3 0.725 ;
 RECT 2.87 1.975 3 2.105 ;
 RECT 2.085 1.975 2.215 2.105 ;
 RECT 2.085 0.595 2.215 0.725 ;
 RECT 1.31 0.125 1.44 0.255 ;
 RECT 0.84 0.595 0.97 0.725 ;
 RECT 0.84 1.975 0.97 2.105 ;
 RECT 17.795 0.225 17.925 0.355 ;
 RECT 20.075 1.475 20.205 1.605 ;
 RECT 15.38 2.06 15.51 2.19 ;
 RECT 17.55 2.065 17.68 2.195 ;
 RECT 13.77 1.715 13.9 1.845 ;
 RECT 12.38 2.525 12.51 2.655 ;
 RECT 14.505 0.915 14.635 1.045 ;
 RECT 14.82 1.6 14.95 1.73 ;
 RECT 14.34 0.395 14.47 0.525 ;
 RECT 13.77 0.585 13.9 0.715 ;
 RECT 13.77 2.105 13.9 2.235 ;
 RECT 14.34 2.34 14.47 2.47 ;
 RECT 18.335 0.89 18.465 1.02 ;
 RECT 22.75 1.455 22.88 1.585 ;
 RECT 22.19 1.435 22.32 1.565 ;
 RECT 22.19 0.505 22.32 0.635 ;
 RECT 5.945 0.12 6.075 0.25 ;
 RECT 23.695 1.44 23.825 1.57 ;
 RECT 0.405 0.36 0.535 0.49 ;
 RECT 0.405 0.62 0.535 0.75 ;
 RECT 0.405 1.71 0.535 1.84 ;
 RECT 0.405 1.97 0.535 2.1 ;
 RECT 0.405 2.23 0.535 2.36 ;
 RECT 20.075 0.225 20.205 0.355 ;
 RECT 7.17 1.28 7.3 1.41 ;
 RECT 6.215 1.58 6.345 1.71 ;
 RECT 9.425 1.25 9.555 1.38 ;
 RECT 11.695 2.375 11.825 2.505 ;
 RECT 9.58 2.63 9.71 2.76 ;
 RECT 5.13 1.585 5.26 1.715 ;
 RECT 5.33 0.6 5.46 0.73 ;
 RECT 4.29 1.875 4.42 2.005 ;
 RECT 4.29 0.58 4.42 0.71 ;
 RECT 3.73 0.59 3.86 0.72 ;
 RECT 3.695 2.065 3.825 2.195 ;
 RECT 8.46 1.67 8.59 1.8 ;
 RECT 5.945 2.515 6.075 2.645 ;
 RECT 7.62 2.515 7.75 2.645 ;
 RECT 6.85 1.52 6.98 1.65 ;
 RECT 1.31 2.59 1.44 2.72 ;
 RECT 10.38 1.49 10.51 1.62 ;
 RECT 10.735 0.6 10.865 0.73 ;
 RECT 10.155 0.6 10.285 0.73 ;
 RECT 9.595 0.6 9.725 0.73 ;
 RECT 9.02 0.6 9.15 0.73 ;
 RECT 9.02 1.48 9.15 1.61 ;
 RECT 8.46 0.6 8.59 0.73 ;
 RECT 7.65 0.555 7.78 0.685 ;
 RECT 6.85 0.6 6.98 0.73 ;
 RECT 3.905 1.515 4.035 1.645 ;
 RECT 2.665 0.26 2.795 0.39 ;
 RECT 21.715 1.415 21.845 1.545 ;
 RECT 21.715 0.505 21.845 0.635 ;
 RECT 21.155 1.415 21.285 1.545 ;
 RECT 21.155 0.505 21.285 0.635 ;
 RECT 14.82 0.555 14.95 0.685 ;
 RECT 12.825 2.01 12.955 2.14 ;
 RECT 12.965 1.21 13.095 1.34 ;
 RECT 12.825 0.605 12.955 0.735 ;
 RECT 13.385 2.025 13.515 2.155 ;
 RECT 13.385 0.605 13.515 0.735 ;
 RECT 11.485 0.91 11.615 1.04 ;
 RECT 11.705 1.31 11.835 1.44 ;
 RECT 9.79 2.33 9.92 2.46 ;
 RECT 8.68 2.085 8.81 2.215 ;
 RECT 8.64 0.24 8.77 0.37 ;
 RECT 7.81 1.57 7.94 1.7 ;
 RECT 7.48 0.89 7.61 1.02 ;
 RECT 16.43 0.965 16.56 1.095 ;
 RECT 3.02 1.245 3.15 1.375 ;
 RECT 16.945 1.255 17.075 1.385 ;
 RECT 12.265 1.64 12.395 1.77 ;
 RECT 11.645 0.5 11.775 0.63 ;
 RECT 11.125 0.51 11.255 0.64 ;
 RECT 19.47 1.255 19.6 1.385 ;
 RECT 19.425 0.505 19.555 0.635 ;
 LAYER M1 ;
 RECT 16.85 1.17 17.19 1.51 ;
 RECT 16.69 1.845 16.83 2.45 ;
 RECT 15.655 2.385 15.795 2.45 ;
 RECT 15.655 2.45 16.83 2.59 ;
 RECT 15.655 2.59 15.795 2.65 ;
 RECT 17.545 0.585 17.685 1.705 ;
 RECT 16.69 1.705 17.685 1.845 ;
 RECT 17.545 1.845 17.685 2.265 ;
 RECT 16.38 0.925 16.61 0.955 ;
 RECT 16.055 0.955 16.61 1.095 ;
 RECT 16.38 1.095 16.61 1.135 ;
 RECT 16.055 1.095 16.195 1.835 ;
 RECT 13.1 1.775 13.24 2.435 ;
 RECT 12.54 1.635 13.24 1.775 ;
 RECT 12.54 1.775 12.68 2.52 ;
 RECT 12.31 2.52 12.68 2.66 ;
 RECT 14.055 2.135 14.195 2.435 ;
 RECT 13.1 2.435 14.195 2.575 ;
 RECT 15.095 1.86 15.235 1.995 ;
 RECT 14.055 1.995 15.235 2.135 ;
 RECT 15.77 0.63 16.435 0.77 ;
 RECT 15.77 0.77 15.91 1.72 ;
 RECT 15.77 2.045 16.435 2.185 ;
 RECT 15.77 1.86 15.91 2.045 ;
 RECT 15.095 1.72 15.91 1.86 ;
 RECT 9.015 0.55 9.155 1.475 ;
 RECT 8.95 1.475 9.22 1.615 ;
 RECT 10.33 1.385 10.56 1.625 ;
 RECT 9.375 1.245 10.56 1.385 ;
 RECT 10.15 0.55 10.29 1.245 ;
 RECT 9.375 1.21 9.605 1.245 ;
 RECT 9.375 1.385 9.605 1.42 ;
 RECT 8.34 2.085 10.645 2.09 ;
 RECT 6.21 2.08 10.645 2.085 ;
 RECT 8.63 2.045 10.645 2.08 ;
 RECT 8.34 2.185 8.86 2.22 ;
 RECT 6.21 1.945 8.48 2.08 ;
 RECT 7.475 0.835 7.615 1.945 ;
 RECT 6.21 1.715 6.35 1.945 ;
 RECT 6.14 1.575 6.415 1.715 ;
 RECT 8.34 2.09 12.4 2.185 ;
 RECT 10.505 2.185 12.4 2.23 ;
 RECT 12.26 0.52 12.4 2.09 ;
 RECT 5.52 2.23 8.2 2.37 ;
 RECT 8.06 2.465 9.345 2.51 ;
 RECT 4.285 2.37 5.66 2.51 ;
 RECT 4.285 0.53 4.425 2.37 ;
 RECT 8.06 2.37 9.98 2.465 ;
 RECT 9.205 2.325 9.98 2.37 ;
 RECT 6.845 0.55 6.985 1.275 ;
 RECT 5.7 1.275 6.985 1.415 ;
 RECT 6.845 1.415 6.985 1.71 ;
 RECT 2.54 1.38 2.68 1.97 ;
 RECT 2.015 0.59 2.395 0.73 ;
 RECT 2.255 0.73 2.395 0.975 ;
 RECT 2.54 1.115 2.68 1.24 ;
 RECT 2.255 0.975 2.68 1.115 ;
 RECT 2.015 1.97 2.68 2.11 ;
 RECT 2.97 1.205 3.2 1.24 ;
 RECT 2.54 1.24 3.2 1.38 ;
 RECT 2.97 1.38 3.2 1.415 ;
 RECT 22.51 0.36 22.65 0.79 ;
 RECT 21.71 0.36 21.85 1.41 ;
 RECT 21.645 1.41 21.915 1.55 ;
 RECT 21.71 0.22 22.65 0.36 ;
 RECT 22.51 0.79 23.13 0.93 ;
 RECT 19.745 0.36 19.885 0.5 ;
 RECT 17.695 0.22 19.885 0.36 ;
 RECT 19.745 0.5 21.29 0.64 ;
 RECT 21.15 0.435 21.29 0.5 ;
 RECT 21.15 0.64 21.29 1.61 ;
 RECT 13.38 0.385 13.52 2.21 ;
 RECT 14.045 0.385 14.185 0.75 ;
 RECT 13.38 0.245 14.185 0.385 ;
 RECT 14.5 0.89 14.64 1.095 ;
 RECT 14.045 0.75 14.64 0.89 ;
 RECT 8.385 1.765 10.98 1.8 ;
 RECT 8.385 1.665 8.81 1.765 ;
 RECT 8.455 0.545 8.595 1.665 ;
 RECT 11.98 0.365 12.12 1.8 ;
 RECT 8.385 1.8 12.12 1.805 ;
 RECT 8.67 1.805 12.12 1.905 ;
 RECT 12.54 0.365 12.68 1.205 ;
 RECT 10.84 1.905 12.12 1.94 ;
 RECT 11.98 0.225 12.68 0.365 ;
 RECT 12.54 1.205 13.165 1.345 ;
 RECT 5.125 0.6 5.53 0.735 ;
 RECT 5.125 0.735 5.265 1.765 ;
 RECT 6.405 0.41 6.545 0.46 ;
 RECT 5.125 0.595 6.545 0.6 ;
 RECT 5.33 0.46 6.545 0.595 ;
 RECT 7.165 0.41 7.305 1.475 ;
 RECT 6.405 0.27 7.305 0.41 ;
 RECT 11.095 0.46 11.235 0.505 ;
 RECT 11.095 0.645 11.235 0.925 ;
 RECT 11.095 1.065 11.235 1.305 ;
 RECT 11.12 1.445 11.26 1.66 ;
 RECT 10.45 0.925 11.235 1.065 ;
 RECT 11.045 0.505 11.325 0.645 ;
 RECT 10.45 0.38 10.59 0.925 ;
 RECT 9.87 0.38 10.01 0.93 ;
 RECT 9.87 0.24 10.59 0.38 ;
 RECT 9.305 0.93 10.01 1.07 ;
 RECT 7.975 0.375 8.115 1.26 ;
 RECT 9.305 0.375 9.445 0.93 ;
 RECT 7.805 1.26 8.115 1.4 ;
 RECT 7.805 1.4 7.945 1.77 ;
 RECT 7.975 0.235 9.445 0.375 ;
 RECT 11.7 1.26 11.84 1.305 ;
 RECT 11.7 1.445 11.84 1.495 ;
 RECT 11.095 1.305 11.84 1.445 ;
 RECT 3.34 0.505 3.48 1.03 ;
 RECT 3.34 1.17 3.48 2.155 ;
 RECT 5.42 1.13 5.56 1.95 ;
 RECT 4.565 1.95 5.56 2.09 ;
 RECT 4.005 0.36 4.145 1.03 ;
 RECT 4.565 0.36 4.705 1.95 ;
 RECT 3.34 1.03 4.145 1.17 ;
 RECT 4.005 0.22 4.705 0.36 ;
 RECT 5.42 0.99 6.705 1.13 ;
 RECT 0.835 0.545 0.975 0.595 ;
 RECT 0.835 0.735 0.975 2.155 ;
 RECT 1.71 0.445 1.85 0.595 ;
 RECT 0.835 0.595 1.85 0.735 ;
 RECT 1.695 0.43 2.725 0.445 ;
 RECT 1.695 0.305 2.845 0.43 ;
 RECT 2.615 0.22 2.845 0.305 ;
 RECT 23.27 0.435 23.41 1.07 ;
 RECT 22.47 1.07 23.41 1.21 ;
 RECT 23.27 1.21 23.41 1.64 ;
 RECT 19.465 0.64 19.605 0.78 ;
 RECT 19.465 0.92 19.605 1.455 ;
 RECT 19.465 0.78 20.6 0.92 ;
 RECT 19.36 0.5 19.605 0.64 ;
 RECT 19.745 1.33 19.885 2.52 ;
 RECT 17.64 2.52 19.885 2.66 ;
 RECT 22.185 0.64 22.325 1.925 ;
 RECT 20.395 1.33 20.535 1.925 ;
 RECT 22.12 0.5 22.37 0.64 ;
 RECT 20.395 1.925 22.325 2.065 ;
 RECT 19.745 1.19 20.535 1.33 ;
 RECT 20.845 0.92 20.985 1.785 ;
 RECT 20.76 0.78 21.01 0.92 ;
 END
END RSDFFARX1

MACRO RSDFFARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 26.24 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.12 1.13 1.62 1.47 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.775 1.425 2.33 1.805 ;
 RECT 1.865 0.92 2.165 1.06 ;
 RECT 2.025 1.06 2.165 1.425 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.46 2.085 1.82 2.295 ;
 RECT 1.585 2.47 2.1 2.49 ;
 RECT 1.585 2.425 2.11 2.47 ;
 RECT 1.46 2.33 2.11 2.425 ;
 RECT 1.46 2.295 2.1 2.33 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.675 1.44 4.11 1.74 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END RSTB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.375 0.8 11.81 1.12 ;
 END
 ANTENNAGATEAREA 0.066 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.23 1.09 14.735 1.5 ;
 RECT 14.52 1.5 14.66 1.855 ;
 RECT 14.52 0.5 14.66 1.09 ;
 END
 ANTENNADIFFAREA 0.598 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 15.535 1.12 15.925 1.465 ;
 RECT 15.57 1.465 15.71 1.855 ;
 RECT 15.57 0.48 15.71 1.12 ;
 END
 ANTENNADIFFAREA 0.606 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 26.24 2.96 ;
 RECT 9.525 2.615 9.76 2.8 ;
 RECT 5.875 2.51 6.145 2.65 ;
 RECT 2.8 1.97 3.2 2.11 ;
 RECT 7.57 2.51 7.8 2.65 ;
 RECT 13.97 2.275 14.235 2.415 ;
 RECT 11.625 2.37 11.895 2.51 ;
 RECT 15.025 2.275 15.3 2.415 ;
 RECT 15.995 2.275 16.265 2.415 ;
 RECT 0.39 1.64 0.55 2.8 ;
 RECT 1.305 2.565 1.445 2.8 ;
 RECT 3.69 1.955 3.83 2.8 ;
 RECT 12.82 1.94 12.96 2.8 ;
 RECT 16.445 2 16.585 2.8 ;
 RECT 18.135 2.025 18.275 2.8 ;
 RECT 5.94 2.65 6.08 2.8 ;
 RECT 3.06 2.11 3.2 2.8 ;
 RECT 7.615 2.65 7.755 2.8 ;
 RECT 14.035 2.415 14.175 2.8 ;
 RECT 11.69 2.51 11.83 2.8 ;
 RECT 15.09 2.415 15.23 2.8 ;
 RECT 16.06 2.415 16.2 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 26.24 0.08 ;
 RECT 2.8 0.59 3.2 0.73 ;
 RECT 7.58 0.555 7.83 0.695 ;
 RECT 21.095 0.22 21.345 0.36 ;
 RECT 0.39 0.08 0.55 0.84 ;
 RECT 1.305 0.08 1.445 0.36 ;
 RECT 4.845 0.08 4.985 0.8 ;
 RECT 3.725 0.08 3.865 0.79 ;
 RECT 5.94 0.08 6.08 0.32 ;
 RECT 9.59 0.08 9.73 0.78 ;
 RECT 12.82 0.08 12.96 0.785 ;
 RECT 11.635 0.08 11.775 0.65 ;
 RECT 13.96 0.08 14.1 0.575 ;
 RECT 10.73 0.08 10.87 0.78 ;
 RECT 16.04 0.08 16.18 0.575 ;
 RECT 18.135 0.08 18.275 0.815 ;
 RECT 15.09 0.08 15.23 0.575 ;
 RECT 16.495 0.08 16.635 0.865 ;
 RECT 23.86 0.08 24 0.65 ;
 RECT 3.06 0.08 3.2 0.59 ;
 RECT 7.645 0.08 7.785 0.555 ;
 RECT 21.14 0.08 21.28 0.22 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 24.62 1.385 25.115 1.75 ;
 RECT 21.13 2.225 24.88 2.385 ;
 RECT 21.095 1.47 21.325 1.61 ;
 RECT 23.815 1.395 23.955 2.225 ;
 RECT 24.73 1.75 24.87 2.225 ;
 RECT 21.14 1.61 21.28 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 19.05 0.81 19.485 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 3.12 1.415 3.22 2.395 ;
 RECT 3.12 0.35 3.22 1.205 ;
 RECT 2.97 1.205 3.22 1.415 ;
 RECT 11.955 0.205 12.055 1.27 ;
 RECT 11.955 1.49 12.055 2.235 ;
 RECT 11.655 1.27 12.055 1.49 ;
 RECT 5.38 1.095 5.48 2.325 ;
 RECT 5.11 0.38 5.21 0.995 ;
 RECT 5.25 2.325 5.48 2.555 ;
 RECT 5.11 0.995 5.48 1.095 ;
 RECT 10.15 1.06 10.25 2.68 ;
 RECT 10.46 0.37 10.56 0.96 ;
 RECT 12.33 2.475 12.56 2.68 ;
 RECT 10.15 0.96 10.56 1.06 ;
 RECT 10.15 2.68 12.56 2.78 ;
 RECT 17.09 1.835 17.19 2.425 ;
 RECT 17.08 1.605 17.31 1.835 ;
 RECT 15.355 0.105 15.455 0.87 ;
 RECT 15.21 0.87 15.455 0.88 ;
 RECT 15.21 0.88 15.925 0.98 ;
 RECT 15.825 0.205 15.925 0.88 ;
 RECT 17.575 0.205 17.675 0.925 ;
 RECT 15.355 1.085 15.455 1.21 ;
 RECT 15.355 1.31 15.455 2.75 ;
 RECT 15.83 1.31 15.93 2.75 ;
 RECT 15.21 0.98 15.455 1.085 ;
 RECT 18.815 0.205 19.045 0.4 ;
 RECT 15.825 0.105 19.045 0.205 ;
 RECT 15.355 1.21 15.93 1.31 ;
 RECT 17.45 0.925 17.68 1.135 ;
 RECT 23.51 0.275 23.61 1.025 ;
 RECT 23.51 1.255 23.61 1.86 ;
 RECT 23.51 1.025 23.79 1.255 ;
 RECT 3.995 0.35 4.095 1.465 ;
 RECT 3.865 1.465 4.095 1.695 ;
 RECT 3.995 1.695 4.095 2.485 ;
 RECT 17.62 2.605 18.97 2.695 ;
 RECT 18.74 2.475 18.97 2.605 ;
 RECT 17.62 1.425 17.72 2.605 ;
 RECT 17.085 0.385 17.185 1.325 ;
 RECT 17.625 2.695 18.97 2.705 ;
 RECT 17.085 1.325 17.72 1.425 ;
 RECT 2.64 0.44 2.74 2.385 ;
 RECT 2.63 0.23 2.86 0.44 ;
 RECT 7.425 0.87 8 0.97 ;
 RECT 7.9 0.38 8 0.87 ;
 RECT 7.425 0.84 7.67 0.87 ;
 RECT 7.425 0.97 7.67 1.06 ;
 RECT 7.425 0.38 7.525 0.84 ;
 RECT 6.285 1.76 6.385 2.34 ;
 RECT 6.165 1.53 6.395 1.76 ;
 RECT 17.92 0.385 18.02 1.215 ;
 RECT 17.92 1.215 18.195 1.27 ;
 RECT 17.92 1.425 18.02 2.425 ;
 RECT 17.92 1.37 18.195 1.425 ;
 RECT 18.395 1.045 18.495 1.27 ;
 RECT 18.395 1.37 18.495 2.425 ;
 RECT 17.92 1.27 18.495 1.37 ;
 RECT 20.845 1.045 20.945 1.76 ;
 RECT 23.035 1.145 23.135 2.09 ;
 RECT 19.195 0.84 19.425 0.945 ;
 RECT 19.195 1.045 19.425 1.07 ;
 RECT 22 1.86 22.1 2.09 ;
 RECT 18.395 0.385 18.495 0.945 ;
 RECT 18.395 0.945 20.945 1.045 ;
 RECT 20.845 0.145 20.945 0.945 ;
 RECT 21.87 1.545 22.1 1.76 ;
 RECT 22 2.09 23.135 2.19 ;
 RECT 20.845 1.76 22.1 1.86 ;
 RECT 7.12 1.45 7.22 2.345 ;
 RECT 8.215 0.38 8.315 1.24 ;
 RECT 7.12 1.24 8.315 1.34 ;
 RECT 8.215 1.34 8.315 2.46 ;
 RECT 7.12 0.38 7.22 1.24 ;
 RECT 7.12 1.34 7.35 1.45 ;
 RECT 12.915 1.16 13.21 1.22 ;
 RECT 12.915 1.22 14.875 1.32 ;
 RECT 12.915 1.32 13.21 1.39 ;
 RECT 14.775 0.98 14.875 1.22 ;
 RECT 14.775 1.32 14.875 2.745 ;
 RECT 13.11 0.365 13.21 1.16 ;
 RECT 13.11 1.39 13.21 2.47 ;
 RECT 14.3 1.32 14.4 2.755 ;
 RECT 14.775 0.105 14.875 0.88 ;
 RECT 14.27 0.88 14.875 0.98 ;
 RECT 14.27 0.095 14.37 0.88 ;
 RECT 2.145 1.565 2.435 1.795 ;
 RECT 2.335 1.795 2.435 2.385 ;
 RECT 21.425 0.965 21.525 1.145 ;
 RECT 21.425 1.145 22.855 1.245 ;
 RECT 22.755 0.965 22.855 1.145 ;
 RECT 22.565 1.245 22.665 1.86 ;
 RECT 23.035 0.275 23.135 0.865 ;
 RECT 21.425 0.735 21.655 0.965 ;
 RECT 22.755 0.865 23.135 0.965 ;
 RECT 7.89 1.75 7.99 2.475 ;
 RECT 7.76 1.53 7.99 1.63 ;
 RECT 7.76 1.73 7.99 1.75 ;
 RECT 7.42 1.73 7.52 2.34 ;
 RECT 7.42 1.63 7.99 1.73 ;
 RECT 1.395 1.165 1.66 1.23 ;
 RECT 1.09 1.23 1.66 1.33 ;
 RECT 1.395 1.33 1.66 1.395 ;
 RECT 1.56 0.345 1.66 1.165 ;
 RECT 1.56 1.395 1.66 2.385 ;
 RECT 1.09 0.345 1.19 1.23 ;
 RECT 1.09 1.33 1.19 2.385 ;
 RECT 16.78 0.385 16.88 2.405 ;
 RECT 16.68 2.405 16.91 2.635 ;
 RECT 9.32 0.37 9.42 1.21 ;
 RECT 9.32 1.21 9.605 1.42 ;
 RECT 9.32 1.42 9.42 2.16 ;
 RECT 1.865 0.335 1.965 0.875 ;
 RECT 1.865 0.875 2.095 1.105 ;
 RECT 22.475 0.275 22.575 0.865 ;
 RECT 21.85 0.735 22.08 0.865 ;
 RECT 21.85 0.865 22.575 0.965 ;
 RECT 24.115 0.27 24.215 0.745 ;
 RECT 23.97 0.745 24.215 0.975 ;
 RECT 24.115 0.975 24.215 1.855 ;
 RECT 11.375 0.205 11.475 0.865 ;
 RECT 11.375 1.08 11.475 2.235 ;
 RECT 11.375 0.865 11.665 1.08 ;
 RECT 5.7 0.38 5.8 1.23 ;
 RECT 5.7 1.46 5.8 2.34 ;
 RECT 5.7 1.23 5.93 1.46 ;
 RECT 9.85 0.37 9.95 2.28 ;
 RECT 9.74 2.28 9.97 2.51 ;
 RECT 8.715 1.445 8.815 2.035 ;
 RECT 8.63 2.035 8.86 2.265 ;
 RECT 6.595 0.38 6.695 0.945 ;
 RECT 6.595 1.175 6.695 2.36 ;
 RECT 6.475 0.945 6.705 1.175 ;
 RECT 2.335 0.365 2.435 1.285 ;
 RECT 1.865 1.385 1.965 2.285 ;
 RECT 1.86 2.285 2.09 2.515 ;
 RECT 1.865 1.285 2.435 1.385 ;
 RECT 8.59 0.2 8.89 0.42 ;
 RECT 8.79 0.42 8.89 0.95 ;
 RECT 6.195 0.2 6.295 0.97 ;
 RECT 6.195 0.1 8.89 0.2 ;
 LAYER CO ;
 RECT 5.33 0.6 5.46 0.73 ;
 RECT 4.29 1.875 4.42 2.005 ;
 RECT 4.29 0.58 4.42 0.71 ;
 RECT 3.73 0.59 3.86 0.72 ;
 RECT 3.695 2.065 3.825 2.195 ;
 RECT 8.46 1.67 8.59 1.8 ;
 RECT 5.945 2.515 6.075 2.645 ;
 RECT 7.62 2.515 7.75 2.645 ;
 RECT 6.85 1.52 6.98 1.65 ;
 RECT 1.31 2.625 1.44 2.755 ;
 RECT 0.84 0.595 0.97 0.725 ;
 RECT 0.84 1.975 0.97 2.105 ;
 RECT 18.865 0.225 18.995 0.355 ;
 RECT 21.145 1.475 21.275 1.605 ;
 RECT 20.54 1.255 20.67 1.385 ;
 RECT 20.495 0.505 20.625 0.635 ;
 RECT 18.79 2.525 18.92 2.655 ;
 RECT 14.525 1.675 14.655 1.805 ;
 RECT 12.38 2.525 12.51 2.655 ;
 RECT 18.015 1.255 18.145 1.385 ;
 RECT 10.38 1.49 10.51 1.62 ;
 RECT 10.735 0.6 10.865 0.73 ;
 RECT 15.26 0.915 15.39 1.045 ;
 RECT 15.575 1.675 15.705 1.805 ;
 RECT 15.095 0.395 15.225 0.525 ;
 RECT 14.525 0.555 14.655 0.685 ;
 RECT 15.095 2.28 15.225 2.41 ;
 RECT 16.045 0.395 16.175 0.525 ;
 RECT 16.065 2.28 16.195 2.41 ;
 RECT 13.965 0.395 14.095 0.525 ;
 RECT 14.04 2.28 14.17 2.41 ;
 RECT 19.245 0.89 19.375 1.02 ;
 RECT 21.92 1.595 22.05 1.725 ;
 RECT 16.73 2.455 16.86 2.585 ;
 RECT 17.13 1.655 17.26 1.785 ;
 RECT 21.475 0.785 21.605 0.915 ;
 RECT 5.945 0.12 6.075 0.25 ;
 RECT 24.765 1.44 24.895 1.57 ;
 RECT 0.405 0.36 0.535 0.49 ;
 RECT 0.405 0.62 0.535 0.75 ;
 RECT 0.405 1.71 0.535 1.84 ;
 RECT 0.405 1.97 0.535 2.1 ;
 RECT 0.405 2.23 0.535 2.36 ;
 RECT 21.145 0.225 21.275 0.355 ;
 RECT 11.485 0.91 11.615 1.04 ;
 RECT 9.425 1.25 9.555 1.38 ;
 RECT 2.195 1.615 2.325 1.745 ;
 RECT 12.265 1.64 12.395 1.77 ;
 RECT 11.64 0.47 11.77 0.6 ;
 RECT 11.125 0.47 11.255 0.6 ;
 RECT 11.125 1.48 11.255 1.61 ;
 RECT 11.695 2.375 11.825 2.505 ;
 RECT 3.02 1.245 3.15 1.375 ;
 RECT 10.155 0.6 10.285 0.73 ;
 RECT 9.595 0.6 9.725 0.73 ;
 RECT 9.02 0.6 9.15 0.73 ;
 RECT 9.02 1.48 9.15 1.61 ;
 RECT 8.46 0.6 8.59 0.73 ;
 RECT 7.65 0.555 7.78 0.685 ;
 RECT 6.85 0.6 6.98 0.73 ;
 RECT 4.85 0.6 4.98 0.73 ;
 RECT 3.345 1.975 3.475 2.105 ;
 RECT 3.345 0.595 3.475 0.725 ;
 RECT 2.87 0.595 3 0.725 ;
 RECT 2.87 1.975 3 2.105 ;
 RECT 2.085 1.975 2.215 2.105 ;
 RECT 2.085 0.595 2.215 0.725 ;
 RECT 1.31 0.145 1.44 0.275 ;
 RECT 18.62 0.635 18.75 0.765 ;
 RECT 18.14 0.635 18.27 0.765 ;
 RECT 18.14 2.075 18.27 2.205 ;
 RECT 17.325 2.05 17.455 2.18 ;
 RECT 17.325 0.635 17.455 0.765 ;
 RECT 16.5 0.635 16.63 0.765 ;
 RECT 16.45 2.06 16.58 2.19 ;
 RECT 18.62 2.065 18.75 2.195 ;
 RECT 21.9 0.785 22.03 0.915 ;
 RECT 24.02 0.795 24.15 0.925 ;
 RECT 23.61 1.075 23.74 1.205 ;
 RECT 24.345 0.505 24.475 0.635 ;
 RECT 24.345 1.44 24.475 1.57 ;
 RECT 3.905 1.515 4.035 1.645 ;
 RECT 11.705 1.31 11.835 1.44 ;
 RECT 9.79 2.33 9.92 2.46 ;
 RECT 8.68 2.085 8.81 2.215 ;
 RECT 8.64 0.24 8.77 0.37 ;
 RECT 7.81 1.57 7.94 1.7 ;
 RECT 7.48 0.89 7.61 1.02 ;
 RECT 7.17 1.28 7.3 1.41 ;
 RECT 6.215 1.58 6.345 1.71 ;
 RECT 17.5 0.965 17.63 1.095 ;
 RECT 2.68 0.27 2.81 0.4 ;
 RECT 12.265 0.57 12.395 0.7 ;
 RECT 23.865 0.47 23.995 0.6 ;
 RECT 23.82 1.455 23.95 1.585 ;
 RECT 23.26 1.435 23.39 1.565 ;
 RECT 23.26 0.505 23.39 0.635 ;
 RECT 22.785 1.415 22.915 1.545 ;
 RECT 22.785 0.505 22.915 0.635 ;
 RECT 22.225 1.415 22.355 1.545 ;
 RECT 22.225 0.505 22.355 0.635 ;
 RECT 15.575 0.555 15.705 0.685 ;
 RECT 12.825 2.01 12.955 2.14 ;
 RECT 12.965 1.21 13.095 1.34 ;
 RECT 12.825 0.605 12.955 0.735 ;
 RECT 13.385 2.025 13.515 2.155 ;
 RECT 13.385 0.605 13.515 0.735 ;
 RECT 6.525 0.995 6.655 1.125 ;
 RECT 5.75 1.28 5.88 1.41 ;
 RECT 5.3 2.375 5.43 2.505 ;
 RECT 1.91 2.335 2.04 2.465 ;
 RECT 1.915 0.925 2.045 1.055 ;
 RECT 1.915 0.925 2.045 1.055 ;
 RECT 1.445 1.215 1.575 1.345 ;
 RECT 9.58 2.63 9.71 2.76 ;
 RECT 5.13 1.585 5.26 1.715 ;
 LAYER M1 ;
 RECT 18.71 2.52 20.955 2.66 ;
 RECT 23.255 0.64 23.395 1.925 ;
 RECT 21.465 1.33 21.605 1.925 ;
 RECT 23.19 0.5 23.44 0.64 ;
 RECT 21.465 1.925 23.395 2.065 ;
 RECT 20.815 1.19 21.605 1.33 ;
 RECT 17.92 1.17 18.26 1.51 ;
 RECT 17.125 1.095 17.265 1.835 ;
 RECT 17.45 0.925 17.68 0.955 ;
 RECT 17.125 0.955 17.68 1.095 ;
 RECT 17.45 1.095 17.68 1.135 ;
 RECT 17.76 1.845 17.9 2.45 ;
 RECT 16.725 2.385 16.865 2.45 ;
 RECT 16.725 2.59 16.865 2.65 ;
 RECT 16.725 2.45 17.9 2.59 ;
 RECT 18.615 0.585 18.755 1.705 ;
 RECT 17.76 1.705 18.755 1.845 ;
 RECT 18.615 1.845 18.755 2.265 ;
 RECT 13.38 0.73 14.38 0.87 ;
 RECT 14.24 0.36 14.38 0.73 ;
 RECT 13.38 0.55 13.52 0.73 ;
 RECT 13.38 0.87 13.52 2.21 ;
 RECT 14.8 0.36 14.94 0.75 ;
 RECT 14.24 0.22 14.94 0.36 ;
 RECT 15.255 0.89 15.395 1.095 ;
 RECT 14.8 0.75 15.395 0.89 ;
 RECT 13.66 2.135 13.8 2.435 ;
 RECT 13.1 1.775 13.24 2.435 ;
 RECT 12.54 1.635 13.24 1.775 ;
 RECT 13.1 2.435 13.8 2.575 ;
 RECT 12.54 1.775 12.68 2.52 ;
 RECT 12.31 2.52 12.68 2.66 ;
 RECT 16.065 1.86 16.205 1.995 ;
 RECT 13.66 1.995 16.205 2.135 ;
 RECT 16.065 1.725 16.98 1.86 ;
 RECT 16.075 1.72 16.98 1.725 ;
 RECT 16.84 2.045 17.505 2.185 ;
 RECT 16.84 1.86 16.98 2.045 ;
 RECT 16.84 0.63 17.505 0.77 ;
 RECT 16.84 0.77 16.98 1.72 ;
 RECT 10.33 1.385 10.56 1.625 ;
 RECT 9.375 1.245 10.56 1.385 ;
 RECT 9.375 1.21 9.605 1.245 ;
 RECT 9.375 1.385 9.605 1.42 ;
 RECT 10.15 0.55 10.29 1.245 ;
 RECT 9.015 0.55 9.155 1.475 ;
 RECT 8.95 1.475 9.22 1.615 ;
 RECT 8.385 1.765 10.98 1.8 ;
 RECT 8.385 1.665 8.81 1.765 ;
 RECT 8.455 0.545 8.595 1.665 ;
 RECT 12.54 0.365 12.68 1.205 ;
 RECT 8.67 1.805 12.12 1.905 ;
 RECT 8.385 1.8 12.12 1.805 ;
 RECT 11.98 0.365 12.12 1.8 ;
 RECT 11.98 0.225 12.68 0.365 ;
 RECT 10.84 1.905 12.12 1.94 ;
 RECT 12.54 1.205 13.165 1.345 ;
 RECT 11.12 1.45 11.26 1.66 ;
 RECT 11.08 1.445 11.26 1.45 ;
 RECT 11.08 0.605 11.22 0.925 ;
 RECT 11.08 1.065 11.22 1.305 ;
 RECT 11.055 0.465 11.325 0.605 ;
 RECT 10.45 0.925 11.225 1.065 ;
 RECT 9.87 0.38 10.01 0.93 ;
 RECT 10.45 0.38 10.59 0.925 ;
 RECT 9.87 0.24 10.59 0.38 ;
 RECT 9.305 0.93 10.01 1.07 ;
 RECT 7.975 0.375 8.115 1.26 ;
 RECT 9.305 0.375 9.445 0.93 ;
 RECT 7.805 1.26 8.115 1.4 ;
 RECT 7.805 1.4 7.945 1.77 ;
 RECT 7.975 0.235 9.445 0.375 ;
 RECT 11.7 1.26 11.84 1.305 ;
 RECT 11.7 1.445 11.84 1.495 ;
 RECT 11.08 1.305 11.84 1.445 ;
 RECT 6.845 0.55 6.985 1.275 ;
 RECT 5.7 1.275 6.985 1.415 ;
 RECT 6.845 1.415 6.985 1.71 ;
 RECT 8.34 2.085 10.645 2.09 ;
 RECT 6.205 2.08 10.645 2.085 ;
 RECT 8.63 2.045 10.645 2.08 ;
 RECT 8.34 2.185 8.86 2.22 ;
 RECT 6.205 1.945 8.48 2.08 ;
 RECT 7.475 0.835 7.615 1.945 ;
 RECT 6.21 1.715 6.35 1.945 ;
 RECT 6.14 1.575 6.415 1.715 ;
 RECT 8.34 2.09 12.4 2.185 ;
 RECT 10.505 2.185 12.4 2.23 ;
 RECT 12.26 0.52 12.4 2.09 ;
 RECT 5.125 0.6 5.53 0.735 ;
 RECT 5.125 0.735 5.265 1.765 ;
 RECT 6.405 0.41 6.545 0.46 ;
 RECT 5.125 0.595 6.545 0.6 ;
 RECT 5.33 0.46 6.545 0.595 ;
 RECT 6.405 0.6 6.545 0.61 ;
 RECT 6.405 0.275 7.305 0.41 ;
 RECT 7.165 0.41 7.305 1.475 ;
 RECT 6.405 0.27 7.24 0.275 ;
 RECT 5.52 2.23 8.2 2.37 ;
 RECT 8.06 2.465 9.345 2.51 ;
 RECT 4.285 2.37 5.66 2.51 ;
 RECT 4.285 0.53 4.425 2.37 ;
 RECT 8.06 2.37 9.98 2.465 ;
 RECT 9.205 2.325 9.98 2.37 ;
 RECT 3.34 0.505 3.48 1.03 ;
 RECT 3.34 1.17 3.48 2.155 ;
 RECT 5.42 1.13 5.56 1.95 ;
 RECT 4.565 1.95 5.56 2.09 ;
 RECT 4.005 0.22 4.705 0.36 ;
 RECT 4.005 0.36 4.145 1.03 ;
 RECT 4.565 0.36 4.705 1.95 ;
 RECT 3.34 1.03 4.145 1.17 ;
 RECT 5.42 0.99 6.705 1.13 ;
 RECT 0.835 0.545 0.975 0.605 ;
 RECT 0.835 0.745 0.975 2.155 ;
 RECT 1.69 0.43 1.83 0.605 ;
 RECT 0.805 0.605 1.83 0.745 ;
 RECT 1.69 0.29 2.86 0.43 ;
 RECT 2.63 0.23 2.86 0.29 ;
 RECT 2.63 0.43 2.86 0.44 ;
 RECT 2.47 1.38 2.61 1.97 ;
 RECT 2.47 0.73 2.61 1.24 ;
 RECT 2.015 1.97 2.61 2.11 ;
 RECT 2.015 0.59 2.61 0.73 ;
 RECT 2.97 1.205 3.2 1.24 ;
 RECT 2.47 1.24 3.2 1.38 ;
 RECT 2.97 1.38 3.2 1.415 ;
 RECT 24.34 0.435 24.48 1.07 ;
 RECT 24.34 1.21 24.48 1.64 ;
 RECT 23.54 1.07 24.48 1.21 ;
 RECT 23.58 0.36 23.72 0.79 ;
 RECT 22.78 0.36 22.92 1.41 ;
 RECT 22.78 0.22 23.72 0.36 ;
 RECT 22.715 1.41 22.985 1.55 ;
 RECT 23.58 0.79 24.2 0.93 ;
 RECT 20.535 0.64 20.675 0.78 ;
 RECT 20.535 0.92 20.675 1.455 ;
 RECT 20.535 0.78 21.67 0.92 ;
 RECT 20.43 0.5 20.675 0.64 ;
 RECT 21.915 0.92 22.055 1.785 ;
 RECT 21.83 0.78 22.08 0.92 ;
 RECT 20.815 0.36 20.955 0.5 ;
 RECT 18.765 0.22 20.955 0.36 ;
 RECT 20.815 0.5 22.36 0.64 ;
 RECT 22.22 0.435 22.36 0.5 ;
 RECT 22.22 0.64 22.36 1.61 ;
 RECT 20.815 1.33 20.955 2.52 ;
 END
END RSDFFARX2

MACRO RSDFFNARX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 25.28 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.14 1.135 1.64 1.42 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.78 1.46 2.33 1.795 ;
 RECT 1.83 0.91 2.12 1.05 ;
 RECT 1.97 1.05 2.11 1.46 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.46 2.1 1.9 2.405 ;
 RECT 1.76 2.405 1.9 2.465 ;
 RECT 1.76 2.465 2.09 2.66 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.7 1.44 4.14 1.74 ;
 END
 ANTENNAGATEAREA 0.065 ;
 END RSTB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.38 1.13 11.84 1.555 ;
 END
 ANTENNAGATEAREA 0.042 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 13.765 1.5 13.905 2.295 ;
 RECT 13.765 1.09 14.255 1.5 ;
 RECT 13.765 0.525 13.905 1.09 ;
 END
 ANTENNADIFFAREA 0.501 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.81 1.12 15.21 1.465 ;
 RECT 14.815 1.465 14.955 1.79 ;
 RECT 14.815 0.48 14.955 1.12 ;
 END
 ANTENNADIFFAREA 0.486 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 25.28 2.96 ;
 RECT 9.525 2.615 9.76 2.8 ;
 RECT 2.8 1.97 3.2 2.11 ;
 RECT 7.57 2.51 7.8 2.65 ;
 RECT 5.875 2.51 6.145 2.65 ;
 RECT 11.575 2.37 11.845 2.51 ;
 RECT 1.305 2.58 1.445 2.8 ;
 RECT 0.39 1.64 0.55 2.8 ;
 RECT 3.69 1.905 3.83 2.8 ;
 RECT 12.82 1.94 12.96 2.8 ;
 RECT 15.375 2 15.515 2.8 ;
 RECT 17.065 2.025 17.205 2.8 ;
 RECT 14.335 2.215 14.475 2.8 ;
 RECT 3.06 2.11 3.2 2.8 ;
 RECT 7.615 2.65 7.755 2.8 ;
 RECT 5.94 2.65 6.08 2.8 ;
 RECT 11.64 2.51 11.78 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 25.28 0.08 ;
 RECT 7.58 0.555 7.83 0.695 ;
 RECT 2.8 0.59 3.2 0.73 ;
 RECT 11.57 0.555 11.84 0.695 ;
 RECT 20.025 0.22 20.275 0.36 ;
 RECT 0.39 0.08 0.55 0.84 ;
 RECT 1.305 0.08 1.445 0.315 ;
 RECT 3.725 0.08 3.865 0.79 ;
 RECT 4.845 0.08 4.985 0.8 ;
 RECT 5.94 0.08 6.08 0.32 ;
 RECT 3.06 0.08 3.2 0.59 ;
 RECT 14.335 0.08 14.475 0.575 ;
 RECT 12.82 0.08 12.96 0.785 ;
 RECT 15.425 0.08 15.565 0.865 ;
 RECT 17.065 0.08 17.205 0.815 ;
 RECT 9.59 0.08 9.73 0.78 ;
 RECT 10.73 0.08 10.87 0.63 ;
 RECT 22.79 0.08 22.93 0.65 ;
 RECT 7.645 0.08 7.785 0.555 ;
 RECT 11.635 0.695 11.775 0.705 ;
 RECT 11.635 0.08 11.775 0.555 ;
 RECT 20.07 0.08 20.21 0.22 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 23.645 1.365 24.14 1.765 ;
 RECT 20.06 2.225 23.81 2.385 ;
 RECT 20.025 1.34 20.255 1.48 ;
 RECT 22.745 1.395 22.885 2.225 ;
 RECT 23.66 1.765 23.8 2.225 ;
 RECT 20.07 1.48 20.21 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.195 0.81 18.75 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 21.965 0.275 22.065 0.865 ;
 RECT 21.685 0.965 21.785 1.145 ;
 RECT 21.495 1.245 21.595 1.86 ;
 RECT 20.355 1.145 21.785 1.245 ;
 RECT 21.685 0.865 22.065 0.965 ;
 RECT 20.355 0.735 20.585 0.965 ;
 RECT 7.425 0.87 8 0.97 ;
 RECT 7.9 0.38 8 0.87 ;
 RECT 7.425 0.84 7.67 0.87 ;
 RECT 7.425 0.97 7.67 1.06 ;
 RECT 7.425 0.38 7.525 0.84 ;
 RECT 2.335 1.795 2.435 2.385 ;
 RECT 2.145 1.565 2.435 1.795 ;
 RECT 7.12 1.34 7.35 1.45 ;
 RECT 7.12 0.38 7.22 1.24 ;
 RECT 7.12 1.45 7.22 2.345 ;
 RECT 8.215 0.38 8.315 1.24 ;
 RECT 8.215 1.34 8.315 2.57 ;
 RECT 7.12 1.24 8.315 1.34 ;
 RECT 16.02 1.835 16.12 2.425 ;
 RECT 16.01 1.605 16.24 1.835 ;
 RECT 2.64 0.43 2.74 2.385 ;
 RECT 2.63 0.22 2.86 0.43 ;
 RECT 9.32 0.37 9.42 1.21 ;
 RECT 9.32 1.21 9.605 1.42 ;
 RECT 9.32 1.42 9.42 2.16 ;
 RECT 20.78 0.865 21.505 0.965 ;
 RECT 20.78 0.735 21.01 0.865 ;
 RECT 21.405 0.275 21.505 0.865 ;
 RECT 2.335 0.365 2.435 1.285 ;
 RECT 1.865 1.385 1.965 2.455 ;
 RECT 1.84 2.455 2.07 2.685 ;
 RECT 1.865 1.285 2.435 1.385 ;
 RECT 23.045 0.27 23.145 0.745 ;
 RECT 22.9 0.745 23.145 0.975 ;
 RECT 23.045 0.975 23.145 1.855 ;
 RECT 22.44 0.275 22.54 1.025 ;
 RECT 22.44 1.025 22.72 1.255 ;
 RECT 22.44 1.255 22.54 1.86 ;
 RECT 12.915 1.16 13.21 1.22 ;
 RECT 13.11 0.365 13.21 1.16 ;
 RECT 12.915 1.32 13.21 1.39 ;
 RECT 13.11 1.39 13.21 2.47 ;
 RECT 14.02 0.105 14.12 1.22 ;
 RECT 14.02 1.32 14.12 2.79 ;
 RECT 12.915 1.22 14.12 1.32 ;
 RECT 8.715 1.445 8.815 2.035 ;
 RECT 8.63 2.035 8.86 2.265 ;
 RECT 8.59 0.2 8.89 0.42 ;
 RECT 8.79 0.42 8.89 0.95 ;
 RECT 6.195 0.2 6.295 0.97 ;
 RECT 6.195 0.1 8.89 0.2 ;
 RECT 1.865 0.335 1.965 0.865 ;
 RECT 1.865 0.865 2.095 1.095 ;
 RECT 9.85 0.37 9.95 2.28 ;
 RECT 9.74 2.28 9.97 2.51 ;
 RECT 7.89 1.75 7.99 2.57 ;
 RECT 7.76 1.53 7.99 1.63 ;
 RECT 7.76 1.73 7.99 1.75 ;
 RECT 7.42 1.73 7.52 2.34 ;
 RECT 7.42 1.63 7.99 1.73 ;
 RECT 11.89 0.325 11.99 1.295 ;
 RECT 11.89 1.53 11.99 2.23 ;
 RECT 11.655 1.295 11.99 1.53 ;
 RECT 1.395 1.165 1.66 1.23 ;
 RECT 1.09 1.23 1.66 1.33 ;
 RECT 1.395 1.33 1.66 1.395 ;
 RECT 1.56 0.345 1.66 1.165 ;
 RECT 1.56 1.395 1.66 2.385 ;
 RECT 1.09 0.345 1.19 1.23 ;
 RECT 1.09 1.33 1.19 2.385 ;
 RECT 16.85 1.215 17.125 1.27 ;
 RECT 16.85 1.37 17.125 1.425 ;
 RECT 16.85 1.27 17.425 1.37 ;
 RECT 17.325 1.045 17.425 1.27 ;
 RECT 17.325 1.37 17.425 2.425 ;
 RECT 19.775 1.045 19.875 1.76 ;
 RECT 16.85 0.385 16.95 1.215 ;
 RECT 16.85 1.425 16.95 2.425 ;
 RECT 18.285 0.84 18.515 0.945 ;
 RECT 18.285 1.045 18.515 1.07 ;
 RECT 17.325 0.385 17.425 0.945 ;
 RECT 17.325 0.945 19.875 1.045 ;
 RECT 19.775 0.145 19.875 0.945 ;
 RECT 20.93 1.86 21.03 2.09 ;
 RECT 20.8 1.545 21.03 1.76 ;
 RECT 21.965 1.145 22.065 2.09 ;
 RECT 19.775 1.76 21.03 1.86 ;
 RECT 20.93 2.09 22.065 2.19 ;
 RECT 16.55 2.605 17.9 2.695 ;
 RECT 17.67 2.475 17.9 2.605 ;
 RECT 16.55 1.425 16.65 2.605 ;
 RECT 16.015 0.385 16.115 1.325 ;
 RECT 16.555 2.695 17.9 2.705 ;
 RECT 16.015 1.325 16.65 1.425 ;
 RECT 10.15 2.655 12.575 2.755 ;
 RECT 10.15 1.06 10.25 2.655 ;
 RECT 12.33 2.475 12.56 2.655 ;
 RECT 10.46 0.37 10.56 0.96 ;
 RECT 10.15 0.96 10.56 1.06 ;
 RECT 5.38 1.095 5.48 2.325 ;
 RECT 5.11 0.38 5.21 0.995 ;
 RECT 5.25 2.325 5.48 2.555 ;
 RECT 5.11 0.995 5.48 1.095 ;
 RECT 14.6 0.105 17.975 0.205 ;
 RECT 14.6 0.205 14.7 0.87 ;
 RECT 16.505 0.205 16.605 0.925 ;
 RECT 14.6 1.085 14.7 2.79 ;
 RECT 14.41 0.87 14.7 1.085 ;
 RECT 17.745 0.205 17.975 0.4 ;
 RECT 16.38 0.925 16.61 1.135 ;
 RECT 3.995 0.35 4.095 1.465 ;
 RECT 3.865 1.465 4.095 1.695 ;
 RECT 3.995 1.695 4.095 2.485 ;
 RECT 11.375 0.33 11.475 2.125 ;
 RECT 11.245 2.125 11.475 2.355 ;
 RECT 3.12 0.35 3.22 1.205 ;
 RECT 3.12 1.415 3.22 2.395 ;
 RECT 2.97 1.205 3.22 1.415 ;
 RECT 15.71 0.385 15.81 2.405 ;
 RECT 15.61 2.405 15.84 2.635 ;
 RECT 6.285 1.76 6.385 2.34 ;
 RECT 6.165 1.53 6.395 1.76 ;
 RECT 5.7 0.38 5.8 1.23 ;
 RECT 5.7 1.46 5.8 2.34 ;
 RECT 5.7 1.23 5.93 1.46 ;
 RECT 6.595 0.38 6.695 0.945 ;
 RECT 6.595 1.175 6.695 2.36 ;
 RECT 6.475 0.945 6.705 1.175 ;
 RECT 20.355 0.965 20.455 1.145 ;
 LAYER CO ;
 RECT 15.66 2.455 15.79 2.585 ;
 RECT 16.06 1.655 16.19 1.785 ;
 RECT 17.55 0.635 17.68 0.765 ;
 RECT 14.34 2.28 14.47 2.41 ;
 RECT 11.295 2.175 11.425 2.305 ;
 RECT 3.905 1.515 4.035 1.645 ;
 RECT 17.07 0.635 17.2 0.765 ;
 RECT 17.07 2.075 17.2 2.205 ;
 RECT 16.255 2.05 16.385 2.18 ;
 RECT 16.255 0.635 16.385 0.765 ;
 RECT 15.43 0.635 15.56 0.765 ;
 RECT 15.38 2.06 15.51 2.19 ;
 RECT 17.55 2.065 17.68 2.195 ;
 RECT 7.17 1.28 7.3 1.41 ;
 RECT 6.215 1.58 6.345 1.71 ;
 RECT 6.525 0.995 6.655 1.125 ;
 RECT 5.75 1.28 5.88 1.41 ;
 RECT 5.3 2.375 5.43 2.505 ;
 RECT 1.89 2.505 2.02 2.635 ;
 RECT 1.915 0.915 2.045 1.045 ;
 RECT 7.48 0.89 7.61 1.02 ;
 RECT 16.945 1.255 17.075 1.385 ;
 RECT 3.345 1.975 3.475 2.105 ;
 RECT 3.345 0.595 3.475 0.725 ;
 RECT 2.87 1.975 3 2.105 ;
 RECT 2.085 2.075 2.215 2.205 ;
 RECT 2.085 0.595 2.215 0.725 ;
 RECT 1.31 0.135 1.44 0.265 ;
 RECT 0.84 0.595 0.97 0.725 ;
 RECT 0.84 1.975 0.97 2.105 ;
 RECT 17.795 0.225 17.925 0.355 ;
 RECT 20.075 1.345 20.205 1.475 ;
 RECT 19.47 1.255 19.6 1.385 ;
 RECT 19.425 0.505 19.555 0.635 ;
 RECT 13.77 1.655 13.9 1.785 ;
 RECT 12.38 2.525 12.51 2.655 ;
 RECT 14.46 0.915 14.59 1.045 ;
 RECT 14.82 1.54 14.95 1.67 ;
 RECT 14.34 0.395 14.47 0.525 ;
 RECT 13.77 0.585 13.9 0.715 ;
 RECT 13.77 2.045 13.9 2.175 ;
 RECT 8.46 0.6 8.59 0.73 ;
 RECT 7.65 0.555 7.78 0.685 ;
 RECT 6.85 0.6 6.98 0.73 ;
 RECT 20.83 0.785 20.96 0.915 ;
 RECT 18.335 0.89 18.465 1.02 ;
 RECT 20.85 1.595 20.98 1.725 ;
 RECT 20.405 0.785 20.535 0.915 ;
 RECT 5.945 0.12 6.075 0.25 ;
 RECT 23.695 1.47 23.825 1.6 ;
 RECT 0.405 0.39 0.535 0.52 ;
 RECT 0.405 0.65 0.535 0.78 ;
 RECT 0.405 1.735 0.535 1.865 ;
 RECT 0.405 1.995 0.535 2.125 ;
 RECT 0.405 2.255 0.535 2.385 ;
 RECT 20.075 0.225 20.205 0.355 ;
 RECT 8.64 0.24 8.77 0.37 ;
 RECT 7.81 1.57 7.94 1.7 ;
 RECT 2.195 1.615 2.325 1.745 ;
 RECT 12.265 0.56 12.395 0.69 ;
 RECT 12.265 1.87 12.395 2 ;
 RECT 11.64 0.56 11.77 0.69 ;
 RECT 11.125 0.57 11.255 0.7 ;
 RECT 11.095 1.48 11.225 1.61 ;
 RECT 11.645 2.375 11.775 2.505 ;
 RECT 9.58 2.63 9.71 2.76 ;
 RECT 5.13 1.585 5.26 1.715 ;
 RECT 5.33 0.6 5.46 0.73 ;
 RECT 4.29 1.875 4.42 2.005 ;
 RECT 4.29 0.59 4.42 0.72 ;
 RECT 3.73 0.59 3.86 0.72 ;
 RECT 3.695 2.055 3.825 2.185 ;
 RECT 8.46 1.67 8.59 1.8 ;
 RECT 5.945 2.515 6.075 2.645 ;
 RECT 7.62 2.515 7.75 2.645 ;
 RECT 6.85 1.52 6.98 1.65 ;
 RECT 1.31 2.63 1.44 2.76 ;
 RECT 10.38 1.49 10.51 1.62 ;
 RECT 10.735 0.4 10.865 0.53 ;
 RECT 10.155 0.6 10.285 0.73 ;
 RECT 9.595 0.6 9.725 0.73 ;
 RECT 9.02 0.6 9.15 0.73 ;
 RECT 9.02 1.49 9.15 1.62 ;
 RECT 2.87 0.595 3 0.725 ;
 RECT 2.68 0.26 2.81 0.39 ;
 RECT 9.425 1.25 9.555 1.38 ;
 RECT 22.95 0.795 23.08 0.925 ;
 RECT 22.54 1.075 22.67 1.205 ;
 RECT 23.275 0.505 23.405 0.635 ;
 RECT 23.275 1.44 23.405 1.57 ;
 RECT 22.795 0.47 22.925 0.6 ;
 RECT 22.75 1.455 22.88 1.585 ;
 RECT 22.19 1.435 22.32 1.565 ;
 RECT 22.19 0.505 22.32 0.635 ;
 RECT 21.715 1.415 21.845 1.545 ;
 RECT 21.715 0.505 21.845 0.635 ;
 RECT 21.155 1.415 21.285 1.545 ;
 RECT 21.155 0.505 21.285 0.635 ;
 RECT 14.82 0.555 14.95 0.685 ;
 RECT 12.825 2.01 12.955 2.14 ;
 RECT 12.965 1.21 13.095 1.34 ;
 RECT 12.825 0.605 12.955 0.735 ;
 RECT 13.385 2.025 13.515 2.155 ;
 RECT 13.385 0.605 13.515 0.735 ;
 RECT 11.695 1.35 11.825 1.48 ;
 RECT 9.79 2.33 9.92 2.46 ;
 RECT 8.68 2.085 8.81 2.215 ;
 RECT 16.43 0.965 16.56 1.095 ;
 RECT 1.445 1.215 1.575 1.345 ;
 RECT 3.02 1.245 3.15 1.375 ;
 RECT 4.85 0.6 4.98 0.73 ;
 RECT 17.72 2.525 17.85 2.655 ;
 LAYER M1 ;
 RECT 19.745 0.36 19.885 0.5 ;
 RECT 17.695 0.22 19.885 0.36 ;
 RECT 19.745 0.5 21.29 0.64 ;
 RECT 21.15 0.435 21.29 0.5 ;
 RECT 21.15 0.64 21.29 1.61 ;
 RECT 22.51 0.36 22.65 0.79 ;
 RECT 21.71 0.36 21.85 1.41 ;
 RECT 21.71 0.22 22.65 0.36 ;
 RECT 21.645 1.41 21.915 1.55 ;
 RECT 22.51 0.79 23.13 0.93 ;
 RECT 16.85 1.17 17.19 1.51 ;
 RECT 16.055 1.095 16.195 1.835 ;
 RECT 16.38 0.925 16.61 0.955 ;
 RECT 16.38 1.095 16.61 1.135 ;
 RECT 16.055 0.955 16.61 1.095 ;
 RECT 16.69 1.845 16.83 2.45 ;
 RECT 15.655 2.385 15.795 2.45 ;
 RECT 15.655 2.45 16.83 2.59 ;
 RECT 15.655 2.59 15.795 2.65 ;
 RECT 17.545 0.585 17.685 1.705 ;
 RECT 16.69 1.705 17.685 1.845 ;
 RECT 17.545 1.845 17.685 2.265 ;
 RECT 13.1 1.775 13.24 2.435 ;
 RECT 12.54 1.635 13.24 1.775 ;
 RECT 12.54 1.775 12.68 2.52 ;
 RECT 12.31 2.52 12.68 2.66 ;
 RECT 14.055 2.075 14.195 2.435 ;
 RECT 13.1 2.435 14.195 2.575 ;
 RECT 15.095 1.86 15.235 1.935 ;
 RECT 14.055 1.935 15.235 2.075 ;
 RECT 15.77 2.045 16.435 2.185 ;
 RECT 15.77 1.86 15.91 2.045 ;
 RECT 15.77 0.63 16.435 0.77 ;
 RECT 15.77 0.77 15.91 1.72 ;
 RECT 15.095 1.72 15.91 1.86 ;
 RECT 13.38 0.385 13.52 2.21 ;
 RECT 13.38 0.24 13.52 0.245 ;
 RECT 14.045 0.385 14.185 0.75 ;
 RECT 13.38 0.245 14.185 0.385 ;
 RECT 14.455 0.89 14.595 1.095 ;
 RECT 14.045 0.75 14.595 0.89 ;
 RECT 10.15 0.55 10.29 1.245 ;
 RECT 10.33 1.385 10.56 1.625 ;
 RECT 9.375 1.245 10.56 1.385 ;
 RECT 9.375 1.21 9.605 1.245 ;
 RECT 9.375 1.385 9.605 1.42 ;
 RECT 8.34 2.085 10.645 2.09 ;
 RECT 6.205 2.08 10.645 2.085 ;
 RECT 8.63 2.045 10.645 2.08 ;
 RECT 8.34 2.185 8.86 2.22 ;
 RECT 6.205 1.945 8.48 2.08 ;
 RECT 7.475 0.835 7.615 1.945 ;
 RECT 6.21 1.715 6.35 1.945 ;
 RECT 6.14 1.575 6.415 1.715 ;
 RECT 11.29 2.23 11.43 2.375 ;
 RECT 8.34 2.09 12.4 2.185 ;
 RECT 10.505 2.185 12.4 2.23 ;
 RECT 12.26 0.505 12.4 2.09 ;
 RECT 9.015 0.55 9.155 1.485 ;
 RECT 8.95 1.485 9.22 1.625 ;
 RECT 8.385 1.765 10.935 1.8 ;
 RECT 8.385 1.665 8.81 1.765 ;
 RECT 8.455 0.545 8.595 1.665 ;
 RECT 8.385 1.8 12.12 1.805 ;
 RECT 12.54 0.365 12.68 1.205 ;
 RECT 8.67 1.805 12.12 1.905 ;
 RECT 11.98 0.365 12.12 1.8 ;
 RECT 11.98 0.225 12.68 0.365 ;
 RECT 10.795 1.905 12.12 1.94 ;
 RECT 12.54 1.205 13.165 1.345 ;
 RECT 6.845 0.55 6.985 1.275 ;
 RECT 6.845 1.415 6.985 1.71 ;
 RECT 5.7 1.275 6.985 1.415 ;
 RECT 10.45 0.38 10.59 0.8 ;
 RECT 10.45 0.94 10.59 1.065 ;
 RECT 9.87 0.38 10.01 0.93 ;
 RECT 9.87 0.24 10.59 0.38 ;
 RECT 9.305 0.93 10.01 1.07 ;
 RECT 9.305 0.375 9.445 0.93 ;
 RECT 7.975 0.375 8.115 1.26 ;
 RECT 7.805 1.26 8.115 1.4 ;
 RECT 7.805 1.4 7.945 1.77 ;
 RECT 7.975 0.235 9.445 0.375 ;
 RECT 10.88 0.94 11.02 1.405 ;
 RECT 11.09 1.615 11.23 1.66 ;
 RECT 10.45 0.8 11.26 0.94 ;
 RECT 11.12 0.505 11.26 0.8 ;
 RECT 10.88 1.405 11.23 1.615 ;
 RECT 9.205 2.465 9.345 2.51 ;
 RECT 8.06 2.37 8.2 2.51 ;
 RECT 5.52 2.23 8.2 2.37 ;
 RECT 8.06 2.51 9.345 2.65 ;
 RECT 4.285 2.37 5.66 2.51 ;
 RECT 4.285 0.53 4.425 2.37 ;
 RECT 9.205 2.325 9.98 2.465 ;
 RECT 5.125 0.6 5.53 0.735 ;
 RECT 5.125 0.735 5.265 1.765 ;
 RECT 6.405 0.41 6.545 0.46 ;
 RECT 5.125 0.595 6.545 0.6 ;
 RECT 6.405 0.275 7.305 0.41 ;
 RECT 7.165 0.41 7.305 1.475 ;
 RECT 6.405 0.27 7.24 0.275 ;
 RECT 5.33 0.46 6.545 0.595 ;
 RECT 6.405 0.6 6.545 0.61 ;
 RECT 2.47 0.73 2.61 1.24 ;
 RECT 2.47 1.38 2.61 1.945 ;
 RECT 2.08 2.085 2.22 2.275 ;
 RECT 2.08 1.945 2.61 2.085 ;
 RECT 2.015 0.59 2.61 0.73 ;
 RECT 2.97 1.205 3.2 1.24 ;
 RECT 2.47 1.24 3.2 1.38 ;
 RECT 2.97 1.38 3.2 1.415 ;
 RECT 3.34 0.505 3.48 1.03 ;
 RECT 3.34 1.17 3.48 2.155 ;
 RECT 5.42 1.13 5.56 1.95 ;
 RECT 4.565 1.95 5.56 2.09 ;
 RECT 4.005 0.36 4.145 1.03 ;
 RECT 4.565 0.36 4.705 1.95 ;
 RECT 3.34 1.03 4.145 1.17 ;
 RECT 4.005 0.22 4.705 0.36 ;
 RECT 5.42 0.99 6.705 1.13 ;
 RECT 1.665 0.36 1.805 0.585 ;
 RECT 0.835 0.585 1.805 0.725 ;
 RECT 0.835 0.545 0.975 0.585 ;
 RECT 0.835 0.725 0.975 2.44 ;
 RECT 1.665 0.22 2.86 0.36 ;
 RECT 2.63 0.36 2.86 0.43 ;
 RECT 23.27 0.435 23.41 1.07 ;
 RECT 22.47 1.07 23.41 1.21 ;
 RECT 23.27 1.21 23.41 1.64 ;
 RECT 20.845 0.92 20.985 1.785 ;
 RECT 20.76 0.78 21.01 0.92 ;
 RECT 19.465 0.64 19.605 0.78 ;
 RECT 19.465 0.92 19.605 1.455 ;
 RECT 19.36 0.5 19.605 0.64 ;
 RECT 19.465 0.78 20.6 0.92 ;
 RECT 19.745 1.2 19.885 2.52 ;
 RECT 17.64 2.52 19.885 2.66 ;
 RECT 20.395 1.2 20.535 1.925 ;
 RECT 22.185 0.64 22.325 1.925 ;
 RECT 19.745 1.06 20.535 1.2 ;
 RECT 20.395 1.925 22.325 2.065 ;
 RECT 22.12 0.5 22.37 0.64 ;
 END
END RSDFFNARX1

MACRO RSDFFNARX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 25.92 BY 2.88 ;
 PIN SE
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.14 1.14 1.625 1.42 ;
 END
 ANTENNAGATEAREA 0.108 ;
 END SE

 PIN SI
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.78 1.46 2.33 1.83 ;
 RECT 1.865 0.92 2.165 1.06 ;
 RECT 2.025 1.06 2.165 1.46 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END SI

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.46 2.1 1.74 2.385 ;
 RECT 1.6 2.465 2.26 2.66 ;
 RECT 1.6 2.385 1.74 2.465 ;
 END
 ANTENNAGATEAREA 0.054 ;
 END D

 PIN RSTB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.7 1.44 4.11 1.74 ;
 END
 ANTENNAGATEAREA 0.065 ;
 END RSTB

 PIN CLK
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 11.38 1.1 11.84 1.44 ;
 END
 ANTENNAGATEAREA 0.05 ;
 END CLK

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 14.455 1.09 14.975 1.5 ;
 RECT 14.52 1.5 14.66 1.855 ;
 RECT 14.52 0.525 14.66 1.09 ;
 END
 ANTENNADIFFAREA 0.642 ;
 END Q

 PIN QN
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 15.57 1.12 16.14 1.465 ;
 RECT 15.57 1.465 15.71 1.855 ;
 RECT 15.57 0.48 15.71 1.12 ;
 END
 ANTENNADIFFAREA 0.606 ;
 END QN

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 25.92 2.96 ;
 RECT 9.525 2.615 9.76 2.8 ;
 RECT 5.875 2.51 6.145 2.65 ;
 RECT 2.8 1.97 3.2 2.11 ;
 RECT 7.57 2.51 7.8 2.65 ;
 RECT 13.97 2.275 14.235 2.415 ;
 RECT 11.625 2.37 11.895 2.51 ;
 RECT 15.025 2.275 15.3 2.415 ;
 RECT 15.995 2.275 16.265 2.415 ;
 RECT 0.39 1.64 0.55 2.8 ;
 RECT 1.305 2.54 1.445 2.8 ;
 RECT 3.69 2.045 3.83 2.8 ;
 RECT 12.82 1.94 12.96 2.8 ;
 RECT 17.815 2.025 17.955 2.8 ;
 RECT 5.94 2.65 6.08 2.8 ;
 RECT 3.06 2.11 3.2 2.8 ;
 RECT 7.615 2.65 7.755 2.8 ;
 RECT 14.035 2.415 14.175 2.8 ;
 RECT 11.69 2.51 11.83 2.8 ;
 RECT 15.09 2.415 15.23 2.8 ;
 RECT 16.06 2.415 16.2 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 25.92 0.08 ;
 RECT 2.8 0.59 3.195 0.73 ;
 RECT 7.58 0.555 7.83 0.695 ;
 RECT 11.57 0.565 11.84 0.705 ;
 RECT 20.775 0.22 21.025 0.36 ;
 RECT 1.305 0.08 1.445 0.32 ;
 RECT 0.39 0.08 0.55 0.84 ;
 RECT 4.845 0.08 4.985 0.8 ;
 RECT 3.725 0.08 3.865 0.79 ;
 RECT 5.94 0.08 6.08 0.32 ;
 RECT 9.59 0.08 9.73 0.78 ;
 RECT 10.73 0.08 10.87 0.355 ;
 RECT 13.96 0.08 14.1 0.575 ;
 RECT 12.82 0.08 12.96 0.785 ;
 RECT 17.815 0.08 17.955 0.815 ;
 RECT 15.09 0.08 15.23 0.575 ;
 RECT 16.04 0.08 16.18 0.575 ;
 RECT 23.54 0.08 23.68 0.65 ;
 RECT 3.055 0.08 3.195 0.59 ;
 RECT 7.645 0.08 7.785 0.555 ;
 RECT 11.635 0.08 11.775 0.565 ;
 RECT 20.82 0.08 20.96 0.22 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 24.3 1.385 24.815 1.75 ;
 RECT 20.81 2.225 24.56 2.385 ;
 RECT 20.775 1.47 21.005 1.61 ;
 RECT 23.495 1.395 23.635 2.225 ;
 RECT 24.41 1.75 24.55 2.225 ;
 RECT 20.82 1.61 20.96 2.225 ;
 END
 END VDDG

 PIN RETN
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 18.945 0.81 19.415 1.165 ;
 END
 ANTENNAGATEAREA 0.2 ;
 END RETN

 OBS
 LAYER PO ;
 RECT 16.77 1.835 16.87 2.425 ;
 RECT 16.76 1.605 16.99 1.835 ;
 RECT 21.53 0.865 22.255 0.965 ;
 RECT 21.53 0.735 21.76 0.865 ;
 RECT 22.155 0.275 22.255 0.865 ;
 RECT 10.15 1.06 10.25 2.68 ;
 RECT 10.46 0.37 10.56 0.96 ;
 RECT 12.33 2.475 12.56 2.68 ;
 RECT 10.15 0.96 10.56 1.06 ;
 RECT 10.15 2.68 12.56 2.78 ;
 RECT 6.595 0.38 6.695 0.945 ;
 RECT 6.595 1.175 6.695 2.36 ;
 RECT 6.475 0.945 6.705 1.175 ;
 RECT 6.285 1.76 6.385 2.34 ;
 RECT 6.165 1.53 6.395 1.76 ;
 RECT 12.915 1.16 13.21 1.22 ;
 RECT 12.915 1.22 14.875 1.32 ;
 RECT 12.915 1.32 13.21 1.39 ;
 RECT 14.775 1.04 14.875 1.22 ;
 RECT 14.775 1.32 14.875 2.75 ;
 RECT 14.27 0.095 14.37 0.94 ;
 RECT 13.11 0.365 13.21 1.16 ;
 RECT 13.11 1.39 13.21 2.47 ;
 RECT 14.775 0.105 14.875 0.94 ;
 RECT 14.27 0.94 14.875 1.04 ;
 RECT 14.3 1.32 14.4 2.75 ;
 RECT 2.64 0.43 2.74 2.385 ;
 RECT 2.615 0.22 2.845 0.43 ;
 RECT 2.335 1.8 2.435 2.385 ;
 RECT 2.145 1.565 2.435 1.8 ;
 RECT 9.32 0.37 9.42 1.21 ;
 RECT 9.32 1.21 9.605 1.42 ;
 RECT 9.32 1.42 9.42 2.16 ;
 RECT 7.12 1.34 7.35 1.45 ;
 RECT 7.12 0.38 7.22 1.24 ;
 RECT 7.12 1.45 7.22 2.345 ;
 RECT 8.215 0.38 8.315 1.24 ;
 RECT 7.12 1.24 8.315 1.34 ;
 RECT 8.215 1.34 8.315 2.62 ;
 RECT 2.335 0.365 2.435 1.285 ;
 RECT 1.865 1.385 1.965 2.455 ;
 RECT 1.865 1.285 2.44 1.385 ;
 RECT 1.855 2.455 2.085 2.685 ;
 RECT 3.12 1.415 3.22 2.395 ;
 RECT 3.12 0.35 3.22 1.205 ;
 RECT 2.97 1.205 3.22 1.415 ;
 RECT 7.89 1.75 7.99 2.62 ;
 RECT 7.76 1.53 7.99 1.63 ;
 RECT 7.76 1.73 7.99 1.75 ;
 RECT 7.42 1.73 7.52 2.34 ;
 RECT 7.42 1.63 7.99 1.73 ;
 RECT 1.385 1.165 1.66 1.23 ;
 RECT 1.09 1.23 1.66 1.33 ;
 RECT 1.385 1.33 1.66 1.395 ;
 RECT 1.56 0.345 1.66 1.165 ;
 RECT 1.56 1.395 1.66 2.385 ;
 RECT 1.09 0.345 1.19 1.23 ;
 RECT 1.09 1.33 1.19 2.385 ;
 RECT 21.105 0.965 21.205 1.145 ;
 RECT 21.105 1.145 22.535 1.245 ;
 RECT 22.435 0.965 22.535 1.145 ;
 RECT 22.245 1.245 22.345 1.86 ;
 RECT 22.715 0.275 22.815 0.865 ;
 RECT 21.105 0.735 21.335 0.965 ;
 RECT 22.435 0.865 22.815 0.965 ;
 RECT 17.3 2.605 18.65 2.695 ;
 RECT 18.42 2.475 18.65 2.605 ;
 RECT 17.3 1.425 17.4 2.605 ;
 RECT 16.765 0.385 16.865 1.325 ;
 RECT 17.305 2.695 18.65 2.705 ;
 RECT 16.765 1.325 17.4 1.425 ;
 RECT 6.195 0.1 8.89 0.2 ;
 RECT 8.79 0.42 8.89 0.95 ;
 RECT 8.59 0.2 8.89 0.42 ;
 RECT 6.195 0.2 6.295 0.97 ;
 RECT 5.38 1.095 5.48 2.325 ;
 RECT 5.11 0.38 5.21 0.995 ;
 RECT 5.25 2.325 5.48 2.555 ;
 RECT 5.11 0.995 5.48 1.095 ;
 RECT 18.075 1.045 18.175 1.27 ;
 RECT 18.075 1.37 18.175 2.425 ;
 RECT 17.6 1.27 18.175 1.37 ;
 RECT 20.525 0.145 20.625 0.945 ;
 RECT 20.525 1.045 20.625 1.76 ;
 RECT 17.6 1.215 17.875 1.27 ;
 RECT 17.6 1.37 17.875 1.425 ;
 RECT 22.715 1.145 22.815 2.09 ;
 RECT 21.68 1.86 21.78 2.09 ;
 RECT 21.55 1.545 21.78 1.76 ;
 RECT 19.035 0.84 19.265 0.945 ;
 RECT 19.035 1.045 19.265 1.07 ;
 RECT 18.075 0.385 18.175 0.945 ;
 RECT 18.075 0.945 20.625 1.045 ;
 RECT 17.6 0.385 17.7 1.215 ;
 RECT 17.6 1.425 17.7 2.425 ;
 RECT 21.68 2.09 22.815 2.19 ;
 RECT 20.525 1.76 21.78 1.86 ;
 RECT 15.355 0.105 15.455 0.87 ;
 RECT 15.21 0.87 15.455 0.88 ;
 RECT 15.21 0.88 15.925 0.98 ;
 RECT 15.825 0.205 15.925 0.88 ;
 RECT 17.255 0.205 17.355 0.925 ;
 RECT 15.355 1.085 15.455 1.26 ;
 RECT 15.355 1.36 15.455 2.75 ;
 RECT 15.83 1.36 15.93 2.75 ;
 RECT 15.21 0.98 15.455 1.085 ;
 RECT 18.495 0.205 18.725 0.4 ;
 RECT 15.825 0.105 18.725 0.205 ;
 RECT 15.355 1.26 15.93 1.36 ;
 RECT 17.13 0.925 17.36 1.135 ;
 RECT 9.85 0.37 9.95 2.28 ;
 RECT 9.74 2.28 9.97 2.51 ;
 RECT 16.46 0.385 16.56 2.405 ;
 RECT 16.36 2.405 16.59 2.635 ;
 RECT 5.7 0.38 5.8 1.23 ;
 RECT 5.7 1.46 5.8 2.34 ;
 RECT 5.7 1.23 5.93 1.46 ;
 RECT 3.995 0.35 4.095 1.465 ;
 RECT 3.865 1.465 4.095 1.695 ;
 RECT 3.995 1.695 4.095 2.485 ;
 RECT 23.19 0.275 23.29 1.025 ;
 RECT 23.19 1.255 23.29 1.86 ;
 RECT 23.19 1.025 23.47 1.255 ;
 RECT 11.955 0.33 12.055 1.16 ;
 RECT 11.955 1.38 12.055 2.235 ;
 RECT 11.655 1.16 12.055 1.38 ;
 RECT 23.795 0.27 23.895 0.745 ;
 RECT 23.795 0.975 23.895 1.855 ;
 RECT 23.65 0.745 23.895 0.975 ;
 RECT 1.865 0.335 1.965 0.875 ;
 RECT 1.865 0.875 2.095 1.105 ;
 RECT 11.375 0.33 11.475 2.145 ;
 RECT 11.245 2.145 11.475 2.375 ;
 RECT 7.425 0.38 7.525 0.84 ;
 RECT 7.425 0.87 8 0.97 ;
 RECT 7.9 0.38 8 0.87 ;
 RECT 7.425 0.84 7.67 0.87 ;
 RECT 7.425 0.97 7.67 1.06 ;
 RECT 8.715 1.445 8.815 2.035 ;
 RECT 8.63 2.035 8.86 2.265 ;
 LAYER CO ;
 RECT 8.64 0.24 8.77 0.37 ;
 RECT 7.81 1.57 7.94 1.7 ;
 RECT 7.48 0.89 7.61 1.02 ;
 RECT 7.17 1.28 7.3 1.41 ;
 RECT 6.215 1.58 6.345 1.71 ;
 RECT 6.525 0.995 6.655 1.125 ;
 RECT 5.75 1.28 5.88 1.41 ;
 RECT 5.3 2.375 5.43 2.505 ;
 RECT 1.905 2.505 2.035 2.635 ;
 RECT 1.915 0.925 2.045 1.055 ;
 RECT 1.915 0.925 2.045 1.055 ;
 RECT 11.105 1.48 11.235 1.61 ;
 RECT 11.695 2.375 11.825 2.505 ;
 RECT 9.58 2.63 9.71 2.76 ;
 RECT 5.13 1.585 5.26 1.715 ;
 RECT 5.33 0.6 5.46 0.73 ;
 RECT 4.29 1.875 4.42 2.005 ;
 RECT 4.29 0.59 4.42 0.72 ;
 RECT 3.73 0.59 3.86 0.72 ;
 RECT 3.695 2.095 3.825 2.225 ;
 RECT 8.46 1.67 8.59 1.8 ;
 RECT 5.945 2.515 6.075 2.645 ;
 RECT 7.62 2.515 7.75 2.645 ;
 RECT 6.85 1.52 6.98 1.65 ;
 RECT 1.31 2.615 1.44 2.745 ;
 RECT 10.38 1.49 10.51 1.62 ;
 RECT 1.435 1.215 1.565 1.345 ;
 RECT 2.195 1.615 2.325 1.745 ;
 RECT 12.265 0.57 12.395 0.7 ;
 RECT 10.735 0.12 10.865 0.25 ;
 RECT 10.155 0.6 10.285 0.73 ;
 RECT 9.595 0.6 9.725 0.73 ;
 RECT 18.47 2.525 18.6 2.655 ;
 RECT 16.41 2.455 16.54 2.585 ;
 RECT 16.81 1.655 16.94 1.785 ;
 RECT 18.3 0.615 18.43 0.745 ;
 RECT 17.82 0.615 17.95 0.745 ;
 RECT 17.82 2.075 17.95 2.205 ;
 RECT 17.005 2.05 17.135 2.18 ;
 RECT 17.005 0.615 17.135 0.745 ;
 RECT 18.3 2.065 18.43 2.195 ;
 RECT 14.525 1.675 14.655 1.805 ;
 RECT 12.38 2.525 12.51 2.655 ;
 RECT 21.58 0.785 21.71 0.915 ;
 RECT 23.7 0.795 23.83 0.925 ;
 RECT 23.29 1.075 23.42 1.205 ;
 RECT 24.025 0.505 24.155 0.635 ;
 RECT 24.025 1.44 24.155 1.57 ;
 RECT 9.02 1.48 9.15 1.61 ;
 RECT 8.46 0.6 8.59 0.73 ;
 RECT 7.65 0.555 7.78 0.685 ;
 RECT 6.85 0.6 6.98 0.73 ;
 RECT 4.85 0.6 4.98 0.73 ;
 RECT 3.345 1.975 3.475 2.105 ;
 RECT 3.345 0.595 3.475 0.725 ;
 RECT 2.87 0.595 3 0.725 ;
 RECT 2.87 1.975 3 2.105 ;
 RECT 2.085 1.975 2.215 2.105 ;
 RECT 2.085 0.595 2.215 0.725 ;
 RECT 1.31 0.14 1.44 0.27 ;
 RECT 0.84 0.595 0.97 0.725 ;
 RECT 0.84 1.975 0.97 2.105 ;
 RECT 18.545 0.225 18.675 0.355 ;
 RECT 20.825 1.475 20.955 1.605 ;
 RECT 20.22 1.255 20.35 1.385 ;
 RECT 20.175 0.505 20.305 0.635 ;
 RECT 23.545 0.47 23.675 0.6 ;
 RECT 3.905 1.515 4.035 1.645 ;
 RECT 15.26 0.915 15.39 1.045 ;
 RECT 15.575 1.675 15.705 1.805 ;
 RECT 15.095 0.395 15.225 0.525 ;
 RECT 8.68 2.085 8.81 2.215 ;
 RECT 11.295 2.195 11.425 2.325 ;
 RECT 16.045 0.395 16.175 0.525 ;
 RECT 16.065 2.28 16.195 2.41 ;
 RECT 13.965 0.395 14.095 0.525 ;
 RECT 14.04 2.28 14.17 2.41 ;
 RECT 19.085 0.89 19.215 1.02 ;
 RECT 21.6 1.595 21.73 1.725 ;
 RECT 21.155 0.785 21.285 0.915 ;
 RECT 5.945 0.12 6.075 0.25 ;
 RECT 24.445 1.44 24.575 1.57 ;
 RECT 0.405 0.36 0.535 0.49 ;
 RECT 0.405 0.62 0.535 0.75 ;
 RECT 0.405 1.71 0.535 1.84 ;
 RECT 0.405 1.97 0.535 2.1 ;
 RECT 0.405 2.23 0.535 2.36 ;
 RECT 20.825 0.225 20.955 0.355 ;
 RECT 12.265 1.845 12.395 1.975 ;
 RECT 11.64 0.57 11.77 0.7 ;
 RECT 11.125 0.57 11.255 0.7 ;
 RECT 9.02 0.6 9.15 0.73 ;
 RECT 14.525 0.585 14.655 0.715 ;
 RECT 15.095 2.28 15.225 2.41 ;
 RECT 17.18 0.965 17.31 1.095 ;
 RECT 2.665 0.26 2.795 0.39 ;
 RECT 9.425 1.25 9.555 1.38 ;
 RECT 3.02 1.245 3.15 1.375 ;
 RECT 17.695 1.255 17.825 1.385 ;
 RECT 23.5 1.455 23.63 1.585 ;
 RECT 22.94 1.435 23.07 1.565 ;
 RECT 22.94 0.505 23.07 0.635 ;
 RECT 22.465 1.415 22.595 1.545 ;
 RECT 22.465 0.505 22.595 0.635 ;
 RECT 21.905 1.415 22.035 1.545 ;
 RECT 21.905 0.505 22.035 0.635 ;
 RECT 15.575 0.555 15.705 0.685 ;
 RECT 12.825 2.01 12.955 2.14 ;
 RECT 12.965 1.21 13.095 1.34 ;
 RECT 12.825 0.605 12.955 0.735 ;
 RECT 13.385 2.025 13.515 2.155 ;
 RECT 13.385 0.605 13.515 0.735 ;
 RECT 11.705 1.2 11.835 1.33 ;
 RECT 9.79 2.33 9.92 2.46 ;
 LAYER M1 ;
 RECT 21.145 1.925 23.075 2.065 ;
 RECT 17.13 0.925 17.36 0.955 ;
 RECT 16.805 0.955 17.36 1.095 ;
 RECT 17.13 1.095 17.36 1.135 ;
 RECT 16.805 1.095 16.945 1.835 ;
 RECT 17.6 1.17 17.94 1.51 ;
 RECT 17.44 1.845 17.58 2.45 ;
 RECT 16.405 2.385 16.545 2.45 ;
 RECT 16.405 2.45 17.58 2.59 ;
 RECT 16.405 2.59 16.545 2.65 ;
 RECT 18.295 0.55 18.435 1.705 ;
 RECT 17.44 1.705 18.435 1.845 ;
 RECT 18.295 1.845 18.435 2.265 ;
 RECT 13.66 2.135 13.8 2.435 ;
 RECT 13.1 1.775 13.24 2.435 ;
 RECT 12.54 1.635 13.24 1.775 ;
 RECT 13.1 2.435 13.8 2.575 ;
 RECT 12.54 1.775 12.68 2.52 ;
 RECT 12.31 2.52 12.68 2.66 ;
 RECT 16.065 1.725 16.66 1.86 ;
 RECT 16.065 1.86 16.205 1.995 ;
 RECT 16.075 1.72 16.66 1.725 ;
 RECT 13.66 1.995 16.205 2.135 ;
 RECT 16.52 2.045 17.185 2.185 ;
 RECT 16.52 1.86 16.66 2.045 ;
 RECT 16.52 0.75 16.66 1.72 ;
 RECT 16.52 0.61 17.205 0.75 ;
 RECT 9.015 0.55 9.155 1.475 ;
 RECT 8.95 1.475 9.22 1.615 ;
 RECT 8.385 1.765 10.925 1.8 ;
 RECT 8.385 1.665 8.81 1.765 ;
 RECT 8.455 0.545 8.595 1.665 ;
 RECT 8.385 1.8 12.12 1.805 ;
 RECT 12.54 0.365 12.68 1.205 ;
 RECT 8.67 1.805 12.12 1.905 ;
 RECT 11.98 0.365 12.12 1.8 ;
 RECT 11.98 0.225 12.68 0.365 ;
 RECT 10.785 1.905 12.12 1.94 ;
 RECT 12.54 1.205 13.165 1.345 ;
 RECT 10.33 1.385 10.56 1.625 ;
 RECT 9.375 1.245 10.56 1.385 ;
 RECT 10.15 0.55 10.29 1.245 ;
 RECT 9.375 1.21 9.605 1.245 ;
 RECT 9.375 1.385 9.605 1.42 ;
 RECT 10.45 0.38 10.59 0.71 ;
 RECT 10.45 0.85 10.59 1.065 ;
 RECT 9.87 0.38 10.01 0.93 ;
 RECT 9.87 0.24 10.59 0.38 ;
 RECT 9.305 0.93 10.01 1.07 ;
 RECT 7.975 0.375 8.115 1.26 ;
 RECT 9.305 0.375 9.445 0.93 ;
 RECT 7.805 1.26 8.115 1.4 ;
 RECT 7.805 1.4 7.945 1.77 ;
 RECT 7.975 0.235 9.445 0.375 ;
 RECT 11.1 0.85 11.24 1.66 ;
 RECT 10.45 0.71 11.26 0.85 ;
 RECT 11.12 0.515 11.26 0.71 ;
 RECT 6.845 0.55 6.985 1.275 ;
 RECT 5.7 1.275 6.985 1.415 ;
 RECT 6.845 1.415 6.985 1.71 ;
 RECT 5.52 2.23 8.2 2.37 ;
 RECT 8.06 2.465 9.345 2.51 ;
 RECT 4.285 2.37 5.66 2.51 ;
 RECT 4.285 0.53 4.425 2.37 ;
 RECT 8.06 2.37 9.98 2.465 ;
 RECT 9.205 2.325 9.98 2.37 ;
 RECT 8.34 2.085 10.645 2.09 ;
 RECT 6.205 2.08 10.645 2.085 ;
 RECT 8.63 2.045 10.645 2.08 ;
 RECT 8.34 2.185 8.86 2.22 ;
 RECT 6.205 1.945 8.48 2.08 ;
 RECT 7.475 0.835 7.615 1.945 ;
 RECT 6.21 1.715 6.35 1.945 ;
 RECT 6.14 1.575 6.415 1.715 ;
 RECT 11.29 2.23 11.43 2.395 ;
 RECT 8.34 2.09 12.4 2.185 ;
 RECT 10.505 2.185 12.4 2.23 ;
 RECT 12.26 0.52 12.4 2.09 ;
 RECT 5.125 0.6 5.53 0.735 ;
 RECT 5.125 0.735 5.265 1.765 ;
 RECT 6.405 0.6 6.545 0.61 ;
 RECT 6.405 0.41 6.545 0.46 ;
 RECT 6.405 0.275 7.305 0.41 ;
 RECT 7.165 0.41 7.305 1.475 ;
 RECT 6.405 0.27 7.24 0.275 ;
 RECT 5.125 0.595 6.545 0.6 ;
 RECT 5.33 0.46 6.545 0.595 ;
 RECT 2.47 0.73 2.61 1.24 ;
 RECT 2.47 1.38 2.61 1.97 ;
 RECT 2.015 1.97 2.61 2.11 ;
 RECT 2.015 0.59 2.61 0.73 ;
 RECT 2.97 1.205 3.2 1.24 ;
 RECT 2.47 1.24 3.2 1.38 ;
 RECT 2.97 1.38 3.2 1.415 ;
 RECT 23.26 0.36 23.4 0.79 ;
 RECT 22.46 0.36 22.6 1.41 ;
 RECT 22.395 1.41 22.665 1.55 ;
 RECT 22.46 0.22 23.4 0.36 ;
 RECT 23.26 0.79 23.88 0.93 ;
 RECT 20.495 0.36 20.635 0.5 ;
 RECT 18.445 0.22 20.635 0.36 ;
 RECT 20.495 0.5 22.04 0.64 ;
 RECT 21.9 0.435 22.04 0.5 ;
 RECT 21.9 0.64 22.04 1.61 ;
 RECT 13.38 0.73 14.38 0.87 ;
 RECT 14.24 0.36 14.38 0.73 ;
 RECT 13.38 0.55 13.52 0.73 ;
 RECT 13.38 0.87 13.52 2.21 ;
 RECT 14.8 0.36 14.94 0.75 ;
 RECT 14.24 0.22 14.94 0.36 ;
 RECT 15.255 0.89 15.395 1.095 ;
 RECT 14.8 0.75 15.395 0.89 ;
 RECT 3.34 0.505 3.48 1.03 ;
 RECT 3.34 1.17 3.48 2.155 ;
 RECT 5.42 1.13 5.56 1.95 ;
 RECT 4.565 1.95 5.56 2.09 ;
 RECT 4.565 0.36 4.705 1.95 ;
 RECT 4.005 0.36 4.145 1.03 ;
 RECT 3.34 1.03 4.145 1.17 ;
 RECT 4.005 0.22 4.705 0.36 ;
 RECT 5.42 0.99 6.705 1.13 ;
 RECT 0.835 0.545 0.975 0.585 ;
 RECT 0.835 0.725 0.975 2.155 ;
 RECT 1.64 0.36 1.78 0.585 ;
 RECT 0.83 0.585 1.78 0.725 ;
 RECT 1.635 0.22 2.845 0.36 ;
 RECT 2.615 0.36 2.845 0.43 ;
 RECT 24.02 0.435 24.16 1.07 ;
 RECT 23.22 1.07 24.16 1.21 ;
 RECT 24.02 1.21 24.16 1.64 ;
 RECT 20.215 0.64 20.355 0.78 ;
 RECT 20.215 0.92 20.355 1.455 ;
 RECT 20.11 0.5 20.355 0.64 ;
 RECT 20.215 0.78 21.35 0.92 ;
 RECT 21.595 0.92 21.735 1.785 ;
 RECT 21.51 0.78 21.76 0.92 ;
 RECT 20.495 1.33 20.635 2.52 ;
 RECT 18.39 2.52 20.635 2.66 ;
 RECT 22.935 0.64 23.075 1.925 ;
 RECT 21.145 1.33 21.285 1.925 ;
 RECT 22.87 0.5 23.12 0.64 ;
 RECT 20.495 1.19 21.285 1.33 ;
 END
END RSDFFNARX2

MACRO TNBUFFX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 2.88 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.105 1.155 1.715 1.405 ;
 END
 ANTENNAGATEAREA 0.155 ;
 END ENB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 2.39 2.355 2.53 2.8 ;
 RECT 1.26 2.05 1.4 2.8 ;
 RECT 4.055 2.37 4.195 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 1.26 0.08 1.4 0.825 ;
 RECT 4.055 0.08 4.195 0.7 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 3.16 0.08 3.3 0.74 ;
 RECT 2.685 0.74 3.3 0.88 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.37 0.225 3.005 0.445 ;
 RECT 2.685 0.445 3.005 0.6 ;
 END
 ANTENNAGATEAREA 0.102 ;
 END INP

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.145 1.76 4.73 2.18 ;
 RECT 4.53 0.585 4.705 0.725 ;
 RECT 4.535 0.515 4.675 0.585 ;
 RECT 4.535 0.725 4.705 0.79 ;
 RECT 4.565 0.79 4.705 1.76 ;
 END
 ANTENNADIFFAREA 0.476 ;
 END Z

 OBS
 LAYER PO ;
 RECT 1.875 0.28 1.975 1.68 ;
 RECT 1.045 1.385 1.145 1.68 ;
 RECT 1.045 1.78 1.145 2.58 ;
 RECT 1.515 1.78 1.615 2.57 ;
 RECT 1.045 0.4 1.145 1.155 ;
 RECT 1.045 1.155 1.29 1.385 ;
 RECT 1.045 1.68 1.975 1.78 ;
 RECT 2.405 0.41 2.505 1.09 ;
 RECT 2.175 1.09 2.505 1.205 ;
 RECT 2.175 1.205 2.275 2.79 ;
 RECT 2.405 0.18 2.615 0.41 ;
 RECT 3.01 1.205 3.11 1.61 ;
 RECT 2.985 0.495 3.085 1.105 ;
 RECT 3.01 1.61 3.28 1.84 ;
 RECT 3.01 1.84 3.11 2.58 ;
 RECT 2.985 1.105 3.11 1.205 ;
 RECT 4.175 0.86 4.415 1.09 ;
 RECT 4.315 0.09 4.415 0.86 ;
 RECT 3.46 1.44 3.91 1.655 ;
 RECT 3.46 1.425 4.415 1.44 ;
 RECT 3.6 1.31 4.415 1.425 ;
 RECT 4.315 1.44 4.415 2.79 ;
 LAYER CO ;
 RECT 4.535 0.59 4.665 0.72 ;
 RECT 4.535 2.045 4.665 2.175 ;
 RECT 4.06 0.5 4.19 0.63 ;
 RECT 4.06 2.44 4.19 2.57 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 2.735 0.745 2.865 0.875 ;
 RECT 1.12 1.205 1.25 1.335 ;
 RECT 3.5 1.475 3.63 1.605 ;
 RECT 2.445 0.23 2.575 0.36 ;
 RECT 3.11 1.66 3.24 1.79 ;
 RECT 3.235 2.23 3.365 2.36 ;
 RECT 3.445 0.745 3.575 0.875 ;
 RECT 2.76 1.95 2.89 2.08 ;
 RECT 2.395 2.405 2.525 2.535 ;
 RECT 1.625 0.6 1.755 0.73 ;
 RECT 2.095 0.535 2.225 0.665 ;
 RECT 1.845 1.95 1.975 2.08 ;
 RECT 1.265 2.12 1.395 2.25 ;
 RECT 1.265 0.625 1.395 0.755 ;
 RECT 0.795 0.625 0.925 0.755 ;
 RECT 0.795 2.12 0.925 2.25 ;
 RECT 4.215 0.91 4.345 1.04 ;
 LAYER M1 ;
 RECT 0.79 0.555 0.93 1.555 ;
 RECT 0.79 1.695 0.93 2.32 ;
 RECT 0.79 1.555 1.835 1.655 ;
 RECT 1.695 1.695 3.31 1.795 ;
 RECT 0.79 1.655 3.31 1.695 ;
 RECT 2.09 0.46 2.23 0.595 ;
 RECT 2.09 0.595 2.545 0.735 ;
 RECT 2.405 0.735 2.545 1.095 ;
 RECT 3.44 0.675 3.58 0.865 ;
 RECT 3.44 1.005 3.915 1.095 ;
 RECT 2.405 1.095 3.915 1.235 ;
 RECT 3.775 1.235 3.915 2.225 ;
 RECT 3.165 2.225 3.915 2.365 ;
 RECT 3.44 0.865 4.395 1.005 ;
 RECT 4.145 1.005 4.395 1.045 ;
 RECT 2.09 1.015 2.23 1.375 ;
 RECT 1.62 0.53 1.76 0.875 ;
 RECT 1.62 0.875 2.23 1.015 ;
 RECT 3.495 1.515 3.635 1.945 ;
 RECT 2.09 1.375 3.635 1.515 ;
 RECT 1.665 1.945 3.635 2.085 ;
 END
END TNBUFFX1

MACRO TNBUFFX16
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 13.12 BY 2.88 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.84 0.225 3.155 0.615 ;
 END
 ANTENNAGATEAREA 0.29 ;
 END INP

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.105 1.13 1.715 1.47 ;
 END
 ANTENNAGATEAREA 0.311 ;
 END ENB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 13.12 2.96 ;
 RECT 2.2 2.38 2.34 2.8 ;
 RECT 3.03 2.355 3.17 2.8 ;
 RECT 5.21 2.37 5.35 2.8 ;
 RECT 12.735 2.37 12.875 2.8 ;
 RECT 11.795 2.37 11.935 2.8 ;
 RECT 10.855 2.37 10.995 2.8 ;
 RECT 9.915 2.37 10.055 2.8 ;
 RECT 8.975 2.37 9.115 2.8 ;
 RECT 8.035 2.37 8.175 2.8 ;
 RECT 7.095 2.37 7.235 2.8 ;
 RECT 6.155 2.37 6.295 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.26 2.05 1.4 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 13.12 0.08 ;
 RECT 3.105 0.77 3.57 0.91 ;
 RECT 6.09 0.305 6.365 0.445 ;
 RECT 7.035 0.305 7.31 0.445 ;
 RECT 7.975 0.305 8.25 0.445 ;
 RECT 8.915 0.305 9.19 0.445 ;
 RECT 9.855 0.305 10.13 0.445 ;
 RECT 10.795 0.305 11.07 0.445 ;
 RECT 11.735 0.305 12.01 0.445 ;
 RECT 12.675 0.305 12.95 0.445 ;
 RECT 4.18 0.08 4.32 0.955 ;
 RECT 3.43 0.08 3.57 0.77 ;
 RECT 5.21 0.08 5.35 0.7 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.26 0.08 1.4 0.825 ;
 RECT 6.155 0.08 6.295 0.305 ;
 RECT 7.1 0.08 7.24 0.305 ;
 RECT 8.04 0.08 8.18 0.305 ;
 RECT 8.98 0.08 9.12 0.305 ;
 RECT 9.92 0.08 10.06 0.305 ;
 RECT 10.86 0.08 11 0.305 ;
 RECT 11.8 0.08 11.94 0.305 ;
 RECT 12.74 0.08 12.88 0.305 ;
 END
 END VSS

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 12.62 0.725 12.76 2.04 ;
 RECT 12.175 2.18 12.475 2.365 ;
 RECT 12.175 1.975 12.475 2.04 ;
 RECT 5.58 2.04 12.76 2.18 ;
 RECT 5.62 0.585 12.76 0.725 ;
 END
 ANTENNADIFFAREA 4.85 ;
 END Z

 OBS
 LAYER PO ;
 RECT 2.23 1.18 2.33 1.68 ;
 RECT 2.345 0.28 2.445 1.08 ;
 RECT 1.875 0.28 1.975 1.08 ;
 RECT 1.045 1.36 1.145 1.68 ;
 RECT 1.045 1.78 1.145 2.58 ;
 RECT 1.515 1.78 1.615 2.78 ;
 RECT 1.985 1.78 2.085 2.78 ;
 RECT 1.045 0.4 1.145 1.13 ;
 RECT 1.045 1.13 1.29 1.36 ;
 RECT 1.875 1.08 2.445 1.18 ;
 RECT 1.045 1.68 2.33 1.78 ;
 RECT 2.815 1.095 2.92 1.105 ;
 RECT 2.82 0.41 2.92 1.095 ;
 RECT 3.285 1.205 3.385 2.79 ;
 RECT 3.48 0.495 3.58 1.105 ;
 RECT 2.815 1.205 2.915 2.79 ;
 RECT 2.815 1.105 3.58 1.205 ;
 RECT 2.82 0.18 3.06 0.41 ;
 RECT 3.76 1.76 4.03 1.84 ;
 RECT 3.76 1.84 3.86 2.79 ;
 RECT 3.76 1.205 3.86 1.61 ;
 RECT 4.29 1.205 4.39 1.66 ;
 RECT 4.435 0.49 4.535 1.105 ;
 RECT 3.965 0.495 4.065 1.105 ;
 RECT 3.755 1.66 4.39 1.76 ;
 RECT 4.29 1.76 4.39 2.79 ;
 RECT 3.755 1.61 4.03 1.66 ;
 RECT 3.76 1.105 4.535 1.205 ;
 RECT 4.575 1.44 5.025 1.655 ;
 RECT 4.715 1.31 12.62 1.425 ;
 RECT 8.945 1.19 9.155 1.31 ;
 RECT 7.065 1.19 7.275 1.31 ;
 RECT 4.575 1.425 12.62 1.44 ;
 RECT 12.3 1.19 12.51 1.31 ;
 RECT 10.345 1.19 10.555 1.31 ;
 RECT 12.52 1.44 12.62 2.79 ;
 RECT 12.05 1.44 12.15 2.79 ;
 RECT 11.58 1.44 11.68 2.79 ;
 RECT 11.11 1.44 11.21 2.79 ;
 RECT 10.64 1.44 10.74 2.79 ;
 RECT 10.17 1.44 10.27 2.79 ;
 RECT 9.7 1.44 9.8 2.79 ;
 RECT 9.23 1.44 9.33 2.79 ;
 RECT 8.76 1.44 8.86 2.79 ;
 RECT 8.29 1.44 8.39 2.79 ;
 RECT 7.82 1.44 7.92 2.79 ;
 RECT 7.35 1.44 7.45 2.79 ;
 RECT 6.88 1.44 6.98 2.79 ;
 RECT 6.41 1.44 6.51 2.79 ;
 RECT 5.94 1.44 6.04 2.79 ;
 RECT 5.47 1.19 5.68 1.31 ;
 RECT 5.47 1.44 5.57 2.79 ;
 RECT 10.705 0.97 10.915 1.09 ;
 RECT 9.515 0.97 9.725 1.09 ;
 RECT 7.925 0.97 8.135 1.09 ;
 RECT 5.86 0.97 6.07 1.09 ;
 RECT 11.87 0.97 12.08 1.09 ;
 RECT 12.055 0.09 12.155 0.84 ;
 RECT 11.585 0.09 11.685 0.84 ;
 RECT 11.115 0.09 11.215 0.84 ;
 RECT 10.645 0.09 10.745 0.84 ;
 RECT 10.175 0.09 10.275 0.84 ;
 RECT 9.705 0.09 9.805 0.84 ;
 RECT 9.235 0.09 9.335 0.84 ;
 RECT 8.765 0.09 8.865 0.84 ;
 RECT 8.295 0.09 8.395 0.84 ;
 RECT 7.825 0.09 7.925 0.84 ;
 RECT 7.355 0.09 7.455 0.84 ;
 RECT 6.885 0.09 6.985 0.84 ;
 RECT 6.41 0.09 6.51 0.84 ;
 RECT 5.94 0.09 6.04 0.84 ;
 RECT 5.47 0.09 5.57 0.84 ;
 RECT 12.525 0.09 12.625 0.84 ;
 RECT 5.47 0.84 12.625 0.97 ;
 LAYER CO ;
 RECT 4.615 1.475 4.745 1.605 ;
 RECT 2.89 0.23 3.02 0.36 ;
 RECT 3.86 1.66 3.99 1.79 ;
 RECT 4.55 2.08 4.68 2.21 ;
 RECT 4 2.405 4.13 2.535 ;
 RECT 4.655 0.845 4.785 0.975 ;
 RECT 3.715 0.845 3.845 0.975 ;
 RECT 3.505 2.08 3.635 2.21 ;
 RECT 3.035 2.405 3.165 2.535 ;
 RECT 2.565 0.535 2.695 0.665 ;
 RECT 2.095 0.79 2.225 0.92 ;
 RECT 1.625 0.535 1.755 0.665 ;
 RECT 2.205 2.43 2.335 2.56 ;
 RECT 1.735 2.105 1.865 2.235 ;
 RECT 1.265 2.12 1.395 2.25 ;
 RECT 1.265 0.625 1.395 0.755 ;
 RECT 0.795 0.625 0.925 0.755 ;
 RECT 0.795 2.12 0.925 2.25 ;
 RECT 5.9 0.91 6.03 1.04 ;
 RECT 12.34 1.24 12.47 1.37 ;
 RECT 10.385 1.24 10.515 1.37 ;
 RECT 11.91 0.91 12.04 1.04 ;
 RECT 10.745 0.91 10.875 1.04 ;
 RECT 9.555 0.91 9.685 1.04 ;
 RECT 8.985 1.24 9.115 1.37 ;
 RECT 7.105 1.24 7.235 1.37 ;
 RECT 7.965 0.91 8.095 1.04 ;
 RECT 5.51 1.24 5.64 1.37 ;
 RECT 8.045 0.31 8.175 0.44 ;
 RECT 8.985 0.31 9.115 0.44 ;
 RECT 12.275 0.59 12.405 0.72 ;
 RECT 7.575 0.59 7.705 0.72 ;
 RECT 7.105 0.31 7.235 0.44 ;
 RECT 11.805 0.31 11.935 0.44 ;
 RECT 6.63 0.59 6.76 0.72 ;
 RECT 11.335 0.59 11.465 0.72 ;
 RECT 6.16 0.31 6.29 0.44 ;
 RECT 10.865 0.31 10.995 0.44 ;
 RECT 5.69 0.59 5.82 0.72 ;
 RECT 10.395 0.59 10.525 0.72 ;
 RECT 9.925 0.31 10.055 0.44 ;
 RECT 9.455 0.59 9.585 0.72 ;
 RECT 8.515 0.59 8.645 0.72 ;
 RECT 12.745 0.31 12.875 0.44 ;
 RECT 12.27 2.045 12.4 2.175 ;
 RECT 11.8 2.44 11.93 2.57 ;
 RECT 11.33 2.045 11.46 2.175 ;
 RECT 10.86 2.44 10.99 2.57 ;
 RECT 10.39 2.045 10.52 2.175 ;
 RECT 9.92 2.44 10.05 2.57 ;
 RECT 9.45 2.045 9.58 2.175 ;
 RECT 8.51 2.045 8.64 2.175 ;
 RECT 8.04 2.44 8.17 2.57 ;
 RECT 7.57 2.045 7.7 2.175 ;
 RECT 6.63 2.045 6.76 2.175 ;
 RECT 6.16 2.44 6.29 2.57 ;
 RECT 5.69 2.045 5.82 2.175 ;
 RECT 12.74 2.44 12.87 2.57 ;
 RECT 8.98 2.44 9.11 2.57 ;
 RECT 7.1 2.44 7.23 2.57 ;
 RECT 5.215 0.5 5.345 0.63 ;
 RECT 5.215 2.44 5.345 2.57 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 2.565 2.08 2.695 2.21 ;
 RECT 4.185 0.775 4.315 0.905 ;
 RECT 3.175 0.775 3.305 0.905 ;
 RECT 1.12 1.18 1.25 1.31 ;
 LAYER M1 ;
 RECT 12.335 1.18 12.475 1.645 ;
 RECT 10.38 1.18 10.52 1.645 ;
 RECT 7.1 1.18 7.24 1.645 ;
 RECT 8.98 1.18 9.12 1.645 ;
 RECT 5.505 1.19 5.645 1.645 ;
 RECT 5.505 1.645 12.475 1.785 ;
 RECT 0.79 0.555 0.93 1.655 ;
 RECT 0.79 1.795 0.93 2.32 ;
 RECT 0.79 1.655 4.055 1.795 ;
 RECT 2.56 0.6 2.7 1.095 ;
 RECT 1.62 0.46 2.7 0.6 ;
 RECT 1.62 0.6 1.76 0.735 ;
 RECT 2.56 1.095 5.065 1.235 ;
 RECT 4.925 1.235 5.065 2.4 ;
 RECT 4.625 0.78 5.065 0.865 ;
 RECT 4.625 1.005 5.065 1.095 ;
 RECT 3.9 2.4 5.065 2.54 ;
 RECT 3.71 0.775 3.85 1.095 ;
 RECT 10.695 1.005 10.925 1.045 ;
 RECT 9.505 1.005 9.735 1.045 ;
 RECT 7.915 1.005 8.145 1.045 ;
 RECT 5.85 1.005 6.08 1.045 ;
 RECT 4.625 0.905 12.09 1.005 ;
 RECT 11.86 1.005 12.09 1.045 ;
 RECT 4.625 0.865 12.085 0.905 ;
 RECT 2.09 0.74 2.23 1.375 ;
 RECT 1.665 2.215 2.89 2.24 ;
 RECT 4.61 1.515 4.75 2.075 ;
 RECT 1.665 2.075 4.75 2.215 ;
 RECT 2.09 1.375 4.75 1.515 ;
 END
END TNBUFFX16

MACRO TNBUFFX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.105 1.155 1.715 1.405 ;
 END
 ANTENNAGATEAREA 0.155 ;
 END ENB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 1.26 2.05 1.4 2.8 ;
 RECT 2.39 2.355 2.53 2.8 ;
 RECT 4.055 2.37 4.195 2.8 ;
 RECT 5 2.37 5.14 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 4.935 0.305 5.21 0.445 ;
 RECT 2.685 0.74 3.3 0.88 ;
 RECT 1.26 0.08 1.4 0.825 ;
 RECT 4.055 0.08 4.195 0.7 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 5 0.08 5.14 0.305 ;
 RECT 3.16 0.08 3.3 0.74 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.37 0.225 3.02 0.445 ;
 RECT 2.72 0.445 3.02 0.6 ;
 END
 ANTENNAGATEAREA 0.102 ;
 END INP

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.465 0.585 5.225 0.725 ;
 RECT 4.415 2.04 5.225 2.18 ;
 RECT 4.415 2.18 4.765 2.43 ;
 RECT 5.085 0.725 5.225 2.04 ;
 END
 ANTENNADIFFAREA 0.606 ;
 END Z

 OBS
 LAYER PO ;
 RECT 1.875 0.28 1.975 1.68 ;
 RECT 1.045 1.385 1.145 1.68 ;
 RECT 1.045 1.78 1.145 2.58 ;
 RECT 1.515 1.78 1.615 2.57 ;
 RECT 1.045 0.4 1.145 1.155 ;
 RECT 1.045 1.155 1.29 1.385 ;
 RECT 1.045 1.68 1.975 1.78 ;
 RECT 2.405 0.41 2.505 1.09 ;
 RECT 2.175 1.09 2.505 1.205 ;
 RECT 2.175 1.205 2.275 2.79 ;
 RECT 2.405 0.18 2.615 0.41 ;
 RECT 3.01 1.205 3.11 1.61 ;
 RECT 2.985 0.495 3.085 1.105 ;
 RECT 3.01 1.61 3.28 1.84 ;
 RECT 3.01 1.84 3.11 2.58 ;
 RECT 2.985 1.105 3.11 1.205 ;
 RECT 4.785 0.09 4.885 0.84 ;
 RECT 4.705 0.97 4.915 1.09 ;
 RECT 4.315 0.09 4.415 0.84 ;
 RECT 4.315 0.84 4.915 0.97 ;
 RECT 3.46 1.44 3.91 1.655 ;
 RECT 3.46 1.425 4.885 1.44 ;
 RECT 3.6 1.31 4.885 1.425 ;
 RECT 4.785 1.44 4.885 2.79 ;
 RECT 4.315 1.44 4.415 2.79 ;
 LAYER CO ;
 RECT 5.005 0.31 5.135 0.44 ;
 RECT 4.535 0.59 4.665 0.72 ;
 RECT 5.005 2.44 5.135 2.57 ;
 RECT 4.535 2.045 4.665 2.175 ;
 RECT 4.06 0.5 4.19 0.63 ;
 RECT 4.06 2.44 4.19 2.57 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 2.735 0.745 2.865 0.875 ;
 RECT 1.12 1.205 1.25 1.335 ;
 RECT 3.5 1.475 3.63 1.605 ;
 RECT 2.445 0.23 2.575 0.36 ;
 RECT 3.11 1.66 3.24 1.79 ;
 RECT 3.235 2.23 3.365 2.36 ;
 RECT 3.445 0.745 3.575 0.875 ;
 RECT 2.76 1.95 2.89 2.08 ;
 RECT 2.395 2.405 2.525 2.535 ;
 RECT 1.625 0.6 1.755 0.73 ;
 RECT 2.095 0.535 2.225 0.665 ;
 RECT 1.845 1.95 1.975 2.08 ;
 RECT 1.265 2.12 1.395 2.25 ;
 RECT 1.265 0.625 1.395 0.755 ;
 RECT 0.795 0.625 0.925 0.755 ;
 RECT 0.795 2.12 0.925 2.25 ;
 RECT 4.745 0.91 4.875 1.04 ;
 LAYER M1 ;
 RECT 0.79 0.555 0.93 1.555 ;
 RECT 0.79 1.695 0.93 2.32 ;
 RECT 0.79 1.555 1.835 1.655 ;
 RECT 1.695 1.695 3.31 1.795 ;
 RECT 0.79 1.655 3.31 1.695 ;
 RECT 2.09 0.46 2.23 0.595 ;
 RECT 2.09 0.595 2.545 0.735 ;
 RECT 2.405 0.735 2.545 1.095 ;
 RECT 3.44 0.675 3.58 0.865 ;
 RECT 3.44 1.005 3.915 1.095 ;
 RECT 2.405 1.095 3.915 1.235 ;
 RECT 3.775 1.235 3.915 2.225 ;
 RECT 3.165 2.225 3.915 2.365 ;
 RECT 3.44 0.865 4.945 1.005 ;
 RECT 4.675 1.005 4.945 1.045 ;
 RECT 2.09 1.015 2.23 1.375 ;
 RECT 1.62 0.53 1.76 0.875 ;
 RECT 1.62 0.875 2.23 1.015 ;
 RECT 3.495 1.515 3.635 1.945 ;
 RECT 2.09 1.375 3.635 1.515 ;
 RECT 1.665 1.945 3.635 2.085 ;
 END
END TNBUFFX2

MACRO TNBUFFX32
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 23.68 BY 2.88 ;
 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.74 0.225 5.115 0.635 ;
 END
 ANTENNAGATEAREA 0.58 ;
 END INP

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.105 1.13 1.715 1.43 ;
 END
 ANTENNAGATEAREA 0.551 ;
 END ENB

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 8.595 0.585 22.98 0.725 ;
 RECT 8.555 2.04 23.01 2.18 ;
 RECT 22.67 2.18 23.01 2.185 ;
 RECT 22.67 1.755 23.01 2.04 ;
 RECT 22.76 0.725 22.9 1.755 ;
 END
 ANTENNADIFFAREA 9.698 ;
 END Z

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 23.68 2.96 ;
 RECT 8.185 2.37 8.325 2.8 ;
 RECT 23.27 2.37 23.41 2.8 ;
 RECT 22.29 2.37 22.43 2.8 ;
 RECT 21.35 2.37 21.49 2.8 ;
 RECT 20.41 2.37 20.55 2.8 ;
 RECT 19.47 2.37 19.61 2.8 ;
 RECT 18.53 2.37 18.67 2.8 ;
 RECT 17.59 2.37 17.73 2.8 ;
 RECT 16.65 2.37 16.79 2.8 ;
 RECT 15.71 2.37 15.85 2.8 ;
 RECT 14.77 2.37 14.91 2.8 ;
 RECT 13.83 2.37 13.97 2.8 ;
 RECT 12.89 2.37 13.03 2.8 ;
 RECT 11.95 2.37 12.09 2.8 ;
 RECT 11.01 2.37 11.15 2.8 ;
 RECT 10.07 2.37 10.21 2.8 ;
 RECT 9.13 2.37 9.27 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 RECT 1.26 2.05 1.4 2.8 ;
 RECT 2.2 2.38 2.34 2.8 ;
 RECT 3.145 2.355 3.285 2.8 ;
 RECT 3.975 2.355 4.115 2.8 ;
 RECT 4.915 2.355 5.055 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 23.68 0.08 ;
 RECT 5.26 0.08 5.4 0.955 ;
 RECT 9.065 0.305 9.34 0.445 ;
 RECT 10.01 0.305 10.285 0.445 ;
 RECT 10.95 0.305 11.225 0.445 ;
 RECT 11.89 0.305 12.165 0.445 ;
 RECT 12.83 0.305 13.105 0.445 ;
 RECT 13.77 0.305 14.045 0.445 ;
 RECT 14.71 0.305 14.985 0.445 ;
 RECT 15.65 0.305 15.925 0.445 ;
 RECT 16.59 0.305 16.865 0.445 ;
 RECT 17.53 0.305 17.805 0.445 ;
 RECT 18.47 0.305 18.745 0.445 ;
 RECT 19.41 0.305 19.685 0.445 ;
 RECT 20.345 0.305 20.62 0.445 ;
 RECT 21.285 0.305 21.56 0.445 ;
 RECT 22.23 0.305 22.505 0.445 ;
 RECT 6.2 0.08 6.34 0.955 ;
 RECT 7.14 0.08 7.28 0.955 ;
 RECT 8.185 0.08 8.325 0.7 ;
 RECT 23.235 0.08 23.375 0.51 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 1.26 0.08 1.4 0.825 ;
 RECT 4.32 0.08 4.46 0.955 ;
 RECT 9.13 0.08 9.27 0.305 ;
 RECT 10.075 0.08 10.215 0.305 ;
 RECT 11.015 0.08 11.155 0.305 ;
 RECT 11.955 0.08 12.095 0.305 ;
 RECT 12.895 0.08 13.035 0.305 ;
 RECT 13.835 0.08 13.975 0.305 ;
 RECT 14.775 0.08 14.915 0.305 ;
 RECT 15.715 0.08 15.855 0.305 ;
 RECT 16.655 0.08 16.795 0.305 ;
 RECT 17.595 0.08 17.735 0.305 ;
 RECT 18.535 0.08 18.675 0.305 ;
 RECT 19.475 0.08 19.615 0.305 ;
 RECT 20.41 0.08 20.55 0.305 ;
 RECT 21.35 0.08 21.49 0.305 ;
 RECT 22.295 0.08 22.435 0.305 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 22.085 1.19 22.295 1.31 ;
 RECT 20.845 1.19 21.055 1.31 ;
 RECT 18.965 1.19 19.175 1.31 ;
 RECT 23.015 1.44 23.115 2.79 ;
 RECT 22.545 1.44 22.645 2.79 ;
 RECT 22.075 1.44 22.175 2.79 ;
 RECT 21.605 1.44 21.705 2.79 ;
 RECT 21.135 1.44 21.235 2.79 ;
 RECT 20.665 1.44 20.765 2.79 ;
 RECT 20.195 1.44 20.295 2.79 ;
 RECT 19.725 1.44 19.825 2.79 ;
 RECT 19.255 1.44 19.355 2.79 ;
 RECT 18.785 1.44 18.885 2.79 ;
 RECT 18.315 1.44 18.415 2.79 ;
 RECT 11.92 1.19 12.13 1.31 ;
 RECT 13.32 1.19 13.53 1.31 ;
 RECT 17.085 1.19 17.295 1.31 ;
 RECT 15.275 1.19 15.485 1.31 ;
 RECT 13.145 1.44 13.245 2.79 ;
 RECT 12.675 1.44 12.775 2.79 ;
 RECT 12.205 1.44 12.305 2.79 ;
 RECT 11.735 1.44 11.835 2.79 ;
 RECT 11.265 1.44 11.365 2.79 ;
 RECT 10.795 1.44 10.895 2.79 ;
 RECT 10.325 1.44 10.425 2.79 ;
 RECT 9.855 1.44 9.955 2.79 ;
 RECT 9.385 1.44 9.485 2.79 ;
 RECT 8.915 1.44 9.015 2.79 ;
 RECT 8.445 1.44 8.545 2.79 ;
 RECT 17.845 1.44 17.945 2.79 ;
 RECT 17.375 1.44 17.475 2.79 ;
 RECT 15.025 1.44 15.125 2.79 ;
 RECT 14.555 1.44 14.655 2.79 ;
 RECT 10.9 0.97 11.11 1.09 ;
 RECT 13.68 0.97 13.89 1.09 ;
 RECT 13.15 0.09 13.25 0.84 ;
 RECT 11.27 0.09 11.37 0.84 ;
 RECT 10.8 0.09 10.9 0.84 ;
 RECT 8.835 0.97 9.045 1.09 ;
 RECT 12.49 0.97 12.7 1.09 ;
 RECT 19.505 0.97 19.715 1.09 ;
 RECT 18.23 0.97 18.44 1.09 ;
 RECT 17.475 0.97 17.685 1.09 ;
 RECT 16.32 0.97 16.53 1.09 ;
 RECT 14.845 0.97 15.055 1.09 ;
 RECT 15.03 0.09 15.13 0.84 ;
 RECT 14.56 0.09 14.66 0.84 ;
 RECT 14.09 0.09 14.19 0.84 ;
 RECT 13.62 0.09 13.72 0.84 ;
 RECT 12.68 0.09 12.78 0.84 ;
 RECT 12.21 0.09 12.31 0.84 ;
 RECT 11.74 0.09 11.84 0.84 ;
 RECT 23.02 0.09 23.12 0.84 ;
 RECT 22.55 0.09 22.65 0.84 ;
 RECT 22.08 0.09 22.18 0.84 ;
 RECT 21.61 0.09 21.71 0.84 ;
 RECT 21.14 0.09 21.24 0.84 ;
 RECT 20.67 0.09 20.77 0.84 ;
 RECT 20.2 0.09 20.3 0.84 ;
 RECT 19.73 0.09 19.83 0.84 ;
 RECT 19.26 0.09 19.36 0.84 ;
 RECT 18.79 0.09 18.89 0.84 ;
 RECT 18.32 0.09 18.42 0.84 ;
 RECT 17.85 0.09 17.95 0.84 ;
 RECT 17.38 0.09 17.48 0.84 ;
 RECT 16.91 0.09 17.01 0.84 ;
 RECT 16.44 0.09 16.54 0.84 ;
 RECT 15.97 0.09 16.07 0.84 ;
 RECT 15.5 0.09 15.6 0.84 ;
 RECT 10.33 0.09 10.43 0.84 ;
 RECT 9.86 0.09 9.96 0.84 ;
 RECT 9.385 0.09 9.485 0.84 ;
 RECT 8.915 0.09 9.015 0.84 ;
 RECT 8.445 0.09 8.545 0.84 ;
 RECT 21.29 0.97 21.5 1.09 ;
 RECT 8.445 0.84 23.12 0.97 ;
 RECT 2.23 1.195 2.33 1.68 ;
 RECT 3.285 0.28 3.385 1.095 ;
 RECT 2.815 0.28 2.915 1.095 ;
 RECT 2.345 0.28 2.445 1.095 ;
 RECT 1.875 0.28 1.975 1.095 ;
 RECT 1.045 1.36 1.145 1.68 ;
 RECT 1.045 1.78 1.145 2.58 ;
 RECT 2.925 1.78 3.025 2.78 ;
 RECT 2.455 1.78 2.555 2.78 ;
 RECT 1.985 1.78 2.085 2.78 ;
 RECT 1.515 1.78 1.615 2.78 ;
 RECT 1.045 0.4 1.145 1.13 ;
 RECT 1.045 1.13 1.29 1.36 ;
 RECT 1.875 1.095 3.385 1.195 ;
 RECT 1.045 1.68 3.025 1.78 ;
 RECT 5.045 0.41 5.145 1.105 ;
 RECT 4.575 0.495 4.675 1.105 ;
 RECT 5.515 0.495 5.615 1.105 ;
 RECT 4.105 0.49 4.205 1.105 ;
 RECT 5.17 1.205 5.27 2.79 ;
 RECT 4.7 1.205 4.8 2.79 ;
 RECT 4.23 1.205 4.33 2.79 ;
 RECT 3.76 1.205 3.86 2.79 ;
 RECT 4.86 0.18 5.145 0.41 ;
 RECT 3.76 1.105 5.615 1.205 ;
 RECT 5.64 1.84 5.74 2.79 ;
 RECT 5.64 1.76 5.915 1.84 ;
 RECT 7.05 1.205 7.15 1.66 ;
 RECT 6.58 1.205 6.68 1.66 ;
 RECT 6.11 1.205 6.21 1.66 ;
 RECT 6.455 0.49 6.555 1.105 ;
 RECT 7.395 0.495 7.495 1.105 ;
 RECT 5.985 0.495 6.085 1.105 ;
 RECT 6.925 0.49 7.025 1.105 ;
 RECT 7.05 1.76 7.15 2.79 ;
 RECT 6.58 1.76 6.68 2.79 ;
 RECT 6.11 1.76 6.21 2.79 ;
 RECT 5.64 1.61 5.915 1.66 ;
 RECT 5.985 1.105 7.495 1.205 ;
 RECT 5.64 1.66 7.15 1.76 ;
 RECT 7.34 1.44 7.79 1.655 ;
 RECT 7.34 1.425 23.115 1.44 ;
 RECT 16.905 1.44 17.005 2.79 ;
 RECT 16.435 1.44 16.535 2.79 ;
 RECT 15.965 1.44 16.065 2.79 ;
 RECT 15.495 1.44 15.595 2.79 ;
 RECT 14.085 1.44 14.185 2.79 ;
 RECT 13.615 1.44 13.715 2.79 ;
 RECT 10.04 1.19 10.25 1.31 ;
 RECT 8.445 1.19 8.655 1.31 ;
 RECT 7.675 1.31 23.115 1.425 ;
 LAYER CO ;
 RECT 15.25 0.59 15.38 0.72 ;
 RECT 10.55 0.59 10.68 0.72 ;
 RECT 10.08 0.31 10.21 0.44 ;
 RECT 20.42 0.31 20.55 0.44 ;
 RECT 14.78 0.31 14.91 0.44 ;
 RECT 4.45 2.08 4.58 2.21 ;
 RECT 3.51 2.08 3.64 2.21 ;
 RECT 9.135 0.31 9.265 0.44 ;
 RECT 19.01 0.59 19.14 0.72 ;
 RECT 2.095 0.51 2.225 0.64 ;
 RECT 1.625 0.78 1.755 0.91 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 7.145 0.775 7.275 0.905 ;
 RECT 6.205 0.775 6.335 0.905 ;
 RECT 5.265 0.775 5.395 0.905 ;
 RECT 1.12 1.18 1.25 1.31 ;
 RECT 20.415 2.44 20.545 2.57 ;
 RECT 7.38 1.475 7.51 1.605 ;
 RECT 11.96 1.24 12.09 1.37 ;
 RECT 4.9 0.23 5.03 0.36 ;
 RECT 5.745 1.66 5.875 1.79 ;
 RECT 7.27 2.08 7.4 2.21 ;
 RECT 6.8 2.405 6.93 2.535 ;
 RECT 6.33 2.08 6.46 2.21 ;
 RECT 5.86 2.405 5.99 2.535 ;
 RECT 7.615 0.845 7.745 0.975 ;
 RECT 6.675 0.845 6.805 0.975 ;
 RECT 4.325 0.775 4.455 0.905 ;
 RECT 5.735 0.845 5.865 0.975 ;
 RECT 4.795 0.845 4.925 0.975 ;
 RECT 3.855 0.845 3.985 0.975 ;
 RECT 5.39 2.08 5.52 2.21 ;
 RECT 4.92 2.405 5.05 2.535 ;
 RECT 3.035 0.51 3.165 0.64 ;
 RECT 2.565 0.78 2.695 0.91 ;
 RECT 3.15 2.405 3.28 2.535 ;
 RECT 2.675 2.105 2.805 2.235 ;
 RECT 2.205 2.43 2.335 2.56 ;
 RECT 1.735 2.105 1.865 2.235 ;
 RECT 1.265 2.12 1.395 2.25 ;
 RECT 1.265 0.625 1.395 0.755 ;
 RECT 0.795 0.625 0.925 0.755 ;
 RECT 0.795 2.12 0.925 2.25 ;
 RECT 23.24 0.32 23.37 0.45 ;
 RECT 8.875 0.91 9.005 1.04 ;
 RECT 22.125 1.24 22.255 1.37 ;
 RECT 20.885 1.24 21.015 1.37 ;
 RECT 21.355 2.44 21.485 2.57 ;
 RECT 20.885 2.045 21.015 2.175 ;
 RECT 12.53 0.91 12.66 1.04 ;
 RECT 15.315 1.24 15.445 1.37 ;
 RECT 18.535 2.44 18.665 2.57 ;
 RECT 18.065 2.045 18.195 2.175 ;
 RECT 19.545 0.91 19.675 1.04 ;
 RECT 18.27 0.91 18.4 1.04 ;
 RECT 17.515 0.91 17.645 1.04 ;
 RECT 16.36 0.91 16.49 1.04 ;
 RECT 14.885 0.91 15.015 1.04 ;
 RECT 13.72 0.91 13.85 1.04 ;
 RECT 9.605 0.59 9.735 0.72 ;
 RECT 14.31 0.59 14.44 0.72 ;
 RECT 13.84 0.31 13.97 0.44 ;
 RECT 8.665 0.59 8.795 0.72 ;
 RECT 17.125 1.24 17.255 1.37 ;
 RECT 23.275 2.425 23.405 2.555 ;
 RECT 15.715 2.44 15.845 2.57 ;
 RECT 11.955 2.44 12.085 2.57 ;
 RECT 10.075 2.44 10.205 2.57 ;
 RECT 8.19 0.5 8.32 0.63 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 19.005 1.24 19.135 1.37 ;
 RECT 13.36 1.24 13.49 1.37 ;
 RECT 21.33 0.91 21.46 1.04 ;
 RECT 17.125 2.045 17.255 2.175 ;
 RECT 16.655 2.44 16.785 2.57 ;
 RECT 16.185 2.045 16.315 2.175 ;
 RECT 15.245 2.045 15.375 2.175 ;
 RECT 14.775 2.44 14.905 2.57 ;
 RECT 14.305 2.045 14.435 2.175 ;
 RECT 13.835 2.44 13.965 2.57 ;
 RECT 13.365 2.045 13.495 2.175 ;
 RECT 12.895 2.44 13.025 2.57 ;
 RECT 12.425 2.045 12.555 2.175 ;
 RECT 11.485 2.045 11.615 2.175 ;
 RECT 11.015 2.44 11.145 2.57 ;
 RECT 10.545 2.045 10.675 2.175 ;
 RECT 9.605 2.045 9.735 2.175 ;
 RECT 9.135 2.44 9.265 2.57 ;
 RECT 8.665 2.045 8.795 2.175 ;
 RECT 19.475 2.44 19.605 2.57 ;
 RECT 17.595 2.44 17.725 2.57 ;
 RECT 19.95 0.59 20.08 0.72 ;
 RECT 3.98 2.405 4.11 2.535 ;
 RECT 3.505 0.78 3.635 0.91 ;
 RECT 8.19 2.44 8.32 2.57 ;
 RECT 18.54 0.31 18.67 0.44 ;
 RECT 13.37 0.59 13.5 0.72 ;
 RECT 19.48 0.31 19.61 0.44 ;
 RECT 22.77 0.59 22.9 0.72 ;
 RECT 18.07 0.59 18.2 0.72 ;
 RECT 12.9 0.31 13.03 0.44 ;
 RECT 17.6 0.31 17.73 0.44 ;
 RECT 22.3 0.31 22.43 0.44 ;
 RECT 17.13 0.59 17.26 0.72 ;
 RECT 12.43 0.59 12.56 0.72 ;
 RECT 21.83 0.59 21.96 0.72 ;
 RECT 16.66 0.31 16.79 0.44 ;
 RECT 11.49 0.59 11.62 0.72 ;
 RECT 15.72 0.31 15.85 0.44 ;
 RECT 22.765 2.045 22.895 2.175 ;
 RECT 22.295 2.44 22.425 2.57 ;
 RECT 21.825 2.045 21.955 2.175 ;
 RECT 19.945 2.045 20.075 2.175 ;
 RECT 19.005 2.045 19.135 2.175 ;
 RECT 10.08 1.24 10.21 1.37 ;
 RECT 10.94 0.91 11.07 1.04 ;
 RECT 8.485 1.24 8.615 1.37 ;
 RECT 21.36 0.31 21.49 0.44 ;
 RECT 16.19 0.59 16.32 0.72 ;
 RECT 11.02 0.31 11.15 0.44 ;
 RECT 11.96 0.31 12.09 0.44 ;
 RECT 20.89 0.59 21.02 0.72 ;
 LAYER M1 ;
 RECT 0.79 0.555 0.93 1.655 ;
 RECT 0.79 1.795 0.93 2.32 ;
 RECT 0.79 1.655 5.94 1.795 ;
 RECT 22.12 1.18 22.26 1.645 ;
 RECT 20.88 1.18 21.02 1.645 ;
 RECT 19 1.18 19.14 1.645 ;
 RECT 17.12 1.18 17.26 1.645 ;
 RECT 15.31 1.18 15.45 1.645 ;
 RECT 13.355 1.18 13.495 1.645 ;
 RECT 10.075 1.18 10.215 1.645 ;
 RECT 11.955 1.18 12.095 1.645 ;
 RECT 8.48 1.19 8.62 1.645 ;
 RECT 8.48 1.645 22.26 1.785 ;
 RECT 6.245 1.515 6.385 2.075 ;
 RECT 3.245 1.375 6.385 1.515 ;
 RECT 1.665 2.215 3.005 2.24 ;
 RECT 3.5 0.71 3.64 0.845 ;
 RECT 2.56 0.71 2.7 0.845 ;
 RECT 1.62 0.71 1.76 0.845 ;
 RECT 3.245 0.985 3.385 1.375 ;
 RECT 1.62 0.845 3.64 0.985 ;
 RECT 1.665 2.1 7.515 2.215 ;
 RECT 2.865 2.075 7.515 2.1 ;
 RECT 7.375 1.425 7.515 2.075 ;
 RECT 2.205 0.355 3.99 0.455 ;
 RECT 2.845 0.455 3.99 0.495 ;
 RECT 3.85 0.495 3.99 1.095 ;
 RECT 2.845 0.495 3.285 0.645 ;
 RECT 2.205 0.315 3.285 0.355 ;
 RECT 2.985 0.31 3.285 0.315 ;
 RECT 2.025 0.505 2.345 0.645 ;
 RECT 2.205 0.455 2.345 0.505 ;
 RECT 7.6 0.775 7.81 0.865 ;
 RECT 7.6 1.005 7.81 1.095 ;
 RECT 5.79 2.4 7.81 2.54 ;
 RECT 3.85 1.095 7.81 1.235 ;
 RECT 7.67 1.235 7.81 2.4 ;
 RECT 6.67 0.775 6.81 1.095 ;
 RECT 5.73 0.775 5.87 1.095 ;
 RECT 4.79 0.775 4.93 1.095 ;
 RECT 19.495 1.005 19.725 1.045 ;
 RECT 18.22 1.005 18.45 1.045 ;
 RECT 17.465 1.005 17.695 1.045 ;
 RECT 16.31 1.005 16.54 1.045 ;
 RECT 14.835 1.005 15.065 1.045 ;
 RECT 13.67 1.005 13.9 1.045 ;
 RECT 12.48 1.005 12.71 1.045 ;
 RECT 10.89 1.005 11.12 1.045 ;
 RECT 8.825 1.005 9.055 1.045 ;
 RECT 21.28 1.005 21.51 1.045 ;
 RECT 7.6 0.865 21.58 1.005 ;
 END
END TNBUFFX32

MACRO TNBUFFX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.4 BY 2.88 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.105 1.155 1.715 1.405 ;
 END
 ANTENNAGATEAREA 0.191 ;
 END ENB

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.4 2.96 ;
 RECT 1.26 2.05 1.4 2.8 ;
 RECT 2.405 2.355 2.545 2.8 ;
 RECT 4.055 2.37 4.195 2.8 ;
 RECT 5.94 2.37 6.08 2.8 ;
 RECT 5 2.37 5.14 2.8 ;
 RECT 0.3 1.74 0.44 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.4 0.08 ;
 RECT 4.935 0.305 5.21 0.445 ;
 RECT 5.88 0.305 6.155 0.445 ;
 RECT 2.685 0.805 3.295 0.945 ;
 RECT 1.26 0.08 1.4 0.825 ;
 RECT 4.055 0.08 4.195 0.7 ;
 RECT 0.3 0.08 0.44 0.775 ;
 RECT 5 0.08 5.14 0.305 ;
 RECT 5.945 0.08 6.085 0.305 ;
 RECT 3.155 0.08 3.295 0.805 ;
 END
 END VSS

 PIN INP
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.37 0.225 3.015 0.445 ;
 RECT 2.715 0.445 3.015 0.62 ;
 END
 ANTENNAGATEAREA 0.145 ;
 END INP

 PIN Z
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.47 2.04 5.96 2.18 ;
 RECT 4.465 0.585 5.96 0.725 ;
 RECT 5.375 2.18 5.725 2.43 ;
 RECT 5.82 0.725 5.96 2.04 ;
 END
 ANTENNADIFFAREA 1.214 ;
 END Z

 OBS
 LAYER PO ;
 RECT 1.875 0.28 1.975 1.68 ;
 RECT 1.045 1.385 1.145 1.68 ;
 RECT 1.045 1.78 1.145 2.58 ;
 RECT 1.515 1.78 1.615 2.78 ;
 RECT 1.045 0.4 1.145 1.155 ;
 RECT 1.045 1.155 1.29 1.385 ;
 RECT 1.045 1.68 1.975 1.78 ;
 RECT 2.185 1.09 2.505 1.205 ;
 RECT 2.405 0.41 2.505 1.09 ;
 RECT 2.185 1.205 2.285 2.79 ;
 RECT 2.405 0.18 2.615 0.41 ;
 RECT 3.01 1.205 3.11 1.61 ;
 RECT 2.985 0.495 3.085 1.105 ;
 RECT 3.01 1.61 3.28 1.84 ;
 RECT 3.01 1.84 3.11 2.79 ;
 RECT 2.985 1.105 3.11 1.205 ;
 RECT 4.785 0.09 4.885 0.84 ;
 RECT 4.705 0.97 4.915 1.09 ;
 RECT 5.73 0.09 5.83 0.84 ;
 RECT 5.255 0.09 5.355 0.84 ;
 RECT 4.315 0.09 4.415 0.84 ;
 RECT 4.315 0.84 5.83 0.97 ;
 RECT 3.46 1.44 3.91 1.655 ;
 RECT 5.455 1.19 5.665 1.31 ;
 RECT 3.46 1.425 5.825 1.44 ;
 RECT 3.6 1.31 5.825 1.425 ;
 RECT 5.725 1.44 5.825 2.79 ;
 RECT 5.255 1.44 5.355 2.79 ;
 RECT 4.785 1.44 4.885 2.79 ;
 RECT 4.315 1.19 4.525 1.31 ;
 RECT 4.315 1.44 4.415 2.79 ;
 LAYER CO ;
 RECT 5.495 1.24 5.625 1.37 ;
 RECT 4.355 1.24 4.485 1.37 ;
 RECT 5.95 0.31 6.08 0.44 ;
 RECT 5.475 0.59 5.605 0.72 ;
 RECT 5.005 0.31 5.135 0.44 ;
 RECT 4.535 0.59 4.665 0.72 ;
 RECT 5.475 2.045 5.605 2.175 ;
 RECT 5.005 2.44 5.135 2.57 ;
 RECT 4.535 2.045 4.665 2.175 ;
 RECT 5.945 2.44 6.075 2.57 ;
 RECT 4.06 0.5 4.19 0.63 ;
 RECT 4.06 2.44 4.19 2.57 ;
 RECT 0.305 0.59 0.435 0.72 ;
 RECT 0.305 0.33 0.435 0.46 ;
 RECT 0.305 2.345 0.435 2.475 ;
 RECT 0.305 2.085 0.435 2.215 ;
 RECT 0.305 1.825 0.435 1.955 ;
 RECT 2.735 0.81 2.865 0.94 ;
 RECT 1.12 1.205 1.25 1.335 ;
 RECT 3.5 1.475 3.63 1.605 ;
 RECT 2.445 0.23 2.575 0.36 ;
 RECT 3.11 1.66 3.24 1.79 ;
 RECT 3.235 2.405 3.365 2.535 ;
 RECT 3.445 0.845 3.575 0.975 ;
 RECT 2.76 2.08 2.89 2.21 ;
 RECT 2.41 2.405 2.54 2.535 ;
 RECT 1.625 0.78 1.755 0.91 ;
 RECT 2.095 0.535 2.225 0.665 ;
 RECT 1.845 2.08 1.975 2.21 ;
 RECT 1.265 2.12 1.395 2.25 ;
 RECT 1.265 0.625 1.395 0.755 ;
 RECT 0.795 0.625 0.925 0.755 ;
 RECT 0.795 2.12 0.925 2.25 ;
 RECT 4.745 0.91 4.875 1.04 ;
 LAYER M1 ;
 RECT 5.49 1.18 5.63 1.645 ;
 RECT 4.35 1.19 4.49 1.645 ;
 RECT 4.35 1.645 5.63 1.785 ;
 RECT 0.79 0.555 0.93 1.555 ;
 RECT 0.79 1.695 0.93 2.32 ;
 RECT 0.79 1.555 1.835 1.655 ;
 RECT 1.695 1.695 3.31 1.795 ;
 RECT 0.79 1.655 3.31 1.695 ;
 RECT 3.44 0.775 3.58 0.865 ;
 RECT 3.44 1.005 3.915 1.095 ;
 RECT 2.37 1.095 3.915 1.235 ;
 RECT 3.775 1.235 3.915 2.4 ;
 RECT 3.165 2.4 3.915 2.54 ;
 RECT 2.09 0.595 2.545 0.735 ;
 RECT 2.405 0.735 2.545 1.095 ;
 RECT 2.09 0.46 2.23 0.595 ;
 RECT 3.44 0.865 4.945 1.005 ;
 RECT 4.675 1.005 4.945 1.045 ;
 RECT 2.09 1.015 2.23 1.375 ;
 RECT 1.62 0.71 1.76 0.875 ;
 RECT 1.62 0.875 2.23 1.015 ;
 RECT 3.495 1.515 3.635 2.075 ;
 RECT 2.09 1.375 3.635 1.515 ;
 RECT 1.665 2.075 3.635 2.215 ;
 END
END TNBUFFX4

MACRO LSDNSSX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8 0.08 ;
 RECT 0.615 0.08 0.755 0.54 ;
 RECT 3.075 0.08 3.215 0.59 ;
 RECT 1.95 0.08 2.09 0.57 ;
 RECT 7.385 0.08 7.525 0.89 ;
 RECT 4.065 0.08 4.205 0.59 ;
 RECT 5.03 0.08 5.17 0.59 ;
 RECT 6 0.08 6.14 0.59 ;
 RECT 6.955 0.08 7.095 0.59 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.36 0.84 0.66 1.14 ;
 END
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8 2.96 ;
 RECT 0.615 1.625 0.755 2.8 ;
 RECT 3.115 1.725 3.255 2.8 ;
 RECT 7.385 1.935 7.525 2.8 ;
 RECT 1.955 1.725 2.095 2.8 ;
 RECT 4.065 1.725 4.205 2.8 ;
 RECT 5.03 1.725 5.17 2.8 ;
 RECT 6 1.725 6.14 2.8 ;
 RECT 6.955 1.725 7.095 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.485 1.445 6.625 2.35 ;
 RECT 6.485 0.4 6.625 1.035 ;
 RECT 3.595 1.095 6.78 1.235 ;
 RECT 6.29 1.235 6.78 1.445 ;
 RECT 6.29 1.035 6.78 1.095 ;
 RECT 3.595 1.235 3.735 2.35 ;
 RECT 3.595 0.4 3.735 1.095 ;
 RECT 4.56 1.235 4.7 2.35 ;
 RECT 4.56 0.4 4.7 1.095 ;
 RECT 5.53 1.235 5.67 2.35 ;
 RECT 5.53 0.4 5.67 1.095 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 0.87 0.1 0.97 1.17 ;
 RECT 0.87 1.4 0.97 2.785 ;
 RECT 0.755 1.17 0.985 1.4 ;
 RECT 0.4 0.1 0.5 0.91 ;
 RECT 0.4 1.14 0.5 1.955 ;
 RECT 0.345 0.91 0.575 1.14 ;
 RECT 5.315 0.2 5.415 2.655 ;
 RECT 6.27 0.2 6.37 2.655 ;
 RECT 6.74 0.2 6.84 2.755 ;
 RECT 5.785 2.655 6.37 2.755 ;
 RECT 5.785 0.2 5.885 2.655 ;
 RECT 5.315 0.1 5.885 0.2 ;
 RECT 4.815 0.2 4.915 2.655 ;
 RECT 4.345 0.2 4.445 2.655 ;
 RECT 3.85 0.2 3.95 2.655 ;
 RECT 3.38 0.2 3.48 0.945 ;
 RECT 3.38 1.175 3.48 2.755 ;
 RECT 6.27 0.1 6.84 0.2 ;
 RECT 4.815 2.655 5.415 2.755 ;
 RECT 4.345 0.1 4.915 0.2 ;
 RECT 3.85 2.655 4.445 2.755 ;
 RECT 3.38 0.1 3.95 0.2 ;
 RECT 3.25 0.945 3.48 1.175 ;
 RECT 1.73 0.1 1.83 1.015 ;
 RECT 1.73 1.115 1.83 2.785 ;
 RECT 2.84 0.1 2.94 1.015 ;
 RECT 2.84 1.115 2.94 2.785 ;
 RECT 1.315 1.015 2.94 1.115 ;
 RECT 2.21 0.1 2.31 1.015 ;
 RECT 2.21 1.115 2.31 2.785 ;
 RECT 1.315 0.945 1.545 1.015 ;
 RECT 1.315 1.115 1.545 1.175 ;
 LAYER CO ;
 RECT 1.475 2.31 1.605 2.44 ;
 RECT 1.095 2.065 1.225 2.195 ;
 RECT 7.39 0.43 7.52 0.56 ;
 RECT 7.39 0.69 7.52 0.82 ;
 RECT 2.545 2.135 2.675 2.265 ;
 RECT 1.96 1.795 2.09 1.925 ;
 RECT 1.955 0.39 2.085 0.52 ;
 RECT 2.545 1.75 2.675 1.88 ;
 RECT 1.96 2.31 2.09 2.44 ;
 RECT 2.545 0.47 2.675 0.6 ;
 RECT 0.805 1.22 0.935 1.35 ;
 RECT 7.39 2.265 7.52 2.395 ;
 RECT 7.39 2.005 7.52 2.135 ;
 RECT 3.12 1.795 3.25 1.925 ;
 RECT 3.12 2.31 3.25 2.44 ;
 RECT 1.095 0.45 1.225 0.58 ;
 RECT 0.62 2.31 0.75 2.44 ;
 RECT 3.08 0.39 3.21 0.52 ;
 RECT 1.095 1.615 1.225 1.745 ;
 RECT 0.62 0.34 0.75 0.47 ;
 RECT 0.62 1.735 0.75 1.865 ;
 RECT 0.395 0.96 0.525 1.09 ;
 RECT 0.15 1.535 0.28 1.665 ;
 RECT 0.15 0.33 0.28 0.46 ;
 RECT 3.3 0.995 3.43 1.125 ;
 RECT 6.96 0.39 7.09 0.52 ;
 RECT 6.49 1.75 6.62 1.88 ;
 RECT 6.96 1.795 7.09 1.925 ;
 RECT 6.96 2.31 7.09 2.44 ;
 RECT 6.49 0.47 6.62 0.6 ;
 RECT 6.49 2.135 6.62 2.265 ;
 RECT 6.005 0.39 6.135 0.52 ;
 RECT 5.535 1.75 5.665 1.88 ;
 RECT 6.005 1.795 6.135 1.925 ;
 RECT 6.005 2.31 6.135 2.44 ;
 RECT 5.535 0.47 5.665 0.6 ;
 RECT 5.535 2.135 5.665 2.265 ;
 RECT 5.035 0.39 5.165 0.52 ;
 RECT 4.565 1.75 4.695 1.88 ;
 RECT 5.035 1.795 5.165 1.925 ;
 RECT 5.035 2.31 5.165 2.44 ;
 RECT 4.565 0.47 4.695 0.6 ;
 RECT 4.565 2.135 4.695 2.265 ;
 RECT 3.6 0.47 3.73 0.6 ;
 RECT 3.6 2.135 3.73 2.265 ;
 RECT 4.07 0.39 4.2 0.52 ;
 RECT 3.6 1.75 3.73 1.88 ;
 RECT 4.07 1.795 4.2 1.925 ;
 RECT 4.07 2.31 4.2 2.44 ;
 RECT 1.365 0.995 1.495 1.125 ;
 RECT 1.47 0.39 1.6 0.52 ;
 RECT 1.475 1.795 1.605 1.925 ;
 LAYER M1 ;
 RECT 1.09 0.345 1.23 0.99 ;
 RECT 1.09 1.13 1.23 2.29 ;
 RECT 1.09 0.99 1.56 1.13 ;
 RECT 1.47 1.325 2.965 1.465 ;
 RECT 2.54 0.4 2.68 1.325 ;
 RECT 2.54 1.465 2.68 2.35 ;
 RECT 2.825 1.14 2.965 1.325 ;
 RECT 1.47 1.465 1.61 2.51 ;
 RECT 1.7 0.85 1.84 1.325 ;
 RECT 1.465 0.32 1.605 0.71 ;
 RECT 1.465 0.71 1.84 0.85 ;
 RECT 3.295 0.925 3.435 1 ;
 RECT 3.295 1.14 3.435 1.195 ;
 RECT 2.825 1 3.435 1.14 ;
 RECT 0.08 0.66 0.22 1.285 ;
 RECT 0.08 1.425 0.285 1.435 ;
 RECT 0.145 0.26 0.285 0.52 ;
 RECT 0.08 0.52 0.285 0.66 ;
 RECT 0.145 1.435 0.285 1.74 ;
 RECT 0.08 1.285 0.94 1.425 ;
 RECT 0.8 1.15 0.94 1.285 ;
 END
END LSDNSSX8

MACRO LSDNX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.76 BY 5.76 ;
 PIN VDDH
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 5.04 5.76 5.2 ;
 RECT 3.985 3.965 4.125 5.04 ;
 RECT 3.475 4.075 3.615 5.04 ;
 END
 END VDDH

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.58 3.85 1.875 4.155 ;
 END
 ANTENNAGATEAREA 0.071 ;
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.76 2.96 ;
 RECT 1.435 2.96 1.575 3.71 ;
 RECT 2.415 2.96 2.555 3.205 ;
 RECT 2.415 2.485 2.555 2.8 ;
 END
 END VSS

 PIN VDDL
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.76 0.08 ;
 RECT 1.435 0.08 1.575 1.395 ;
 RECT 1.95 0.08 2.09 1.34 ;
 END
 PORT
 LAYER M1 ;
 RECT 0 5.68 5.76 5.84 ;
 END
 END VDDL

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.58 1.47 1.185 1.755 ;
 RECT 0.945 0.545 1.085 1.47 ;
 END
 ANTENNADIFFAREA 0.499 ;
 END Q

 OBS
 LAYER PO ;
 RECT 0.585 1.72 0.685 3.22 ;
 RECT 0.585 1.48 0.815 1.72 ;
 RECT 0.585 3.22 0.815 3.45 ;
 RECT 1.21 2.975 2.195 3.075 ;
 RECT 1.21 3.075 1.31 3.88 ;
 RECT 1.21 0.36 1.31 2.975 ;
 RECT 1.97 3.075 2.195 3.345 ;
 RECT 3.26 3.945 3.36 4.705 ;
 RECT 1.69 3.295 1.79 3.845 ;
 RECT 1.63 3.87 3.36 3.945 ;
 RECT 1.63 3.945 1.855 4.1 ;
 RECT 1.69 3.845 3.36 3.87 ;
 LAYER CO ;
 RECT 0.95 0.935 1.08 1.065 ;
 RECT 2.42 2.89 2.55 3.02 ;
 RECT 1.955 0.62 2.085 0.75 ;
 RECT 0.635 1.54 0.765 1.67 ;
 RECT 1.44 3.53 1.57 3.66 ;
 RECT 0.95 0.655 1.08 0.785 ;
 RECT 1.44 0.655 1.57 0.785 ;
 RECT 1.44 1.195 1.57 1.325 ;
 RECT 1.955 0.88 2.085 1.01 ;
 RECT 0.635 3.27 0.765 3.4 ;
 RECT 0.95 3.27 1.08 3.4 ;
 RECT 1.44 0.935 1.57 1.065 ;
 RECT 0.95 3.53 1.08 3.66 ;
 RECT 1.955 1.14 2.085 1.27 ;
 RECT 3.99 4.325 4.12 4.455 ;
 RECT 3.99 4.065 4.12 4.195 ;
 RECT 2.015 3.165 2.145 3.295 ;
 RECT 1.44 3.53 1.57 3.66 ;
 RECT 3.01 4.145 3.14 4.275 ;
 RECT 3.48 4.145 3.61 4.275 ;
 RECT 2.42 2.63 2.55 2.76 ;
 RECT 1.675 3.92 1.805 4.05 ;
 RECT 0.95 1.455 1.08 1.585 ;
 RECT 0.95 1.195 1.08 1.325 ;
 RECT 1.91 3.53 2.04 3.66 ;
 LAYER M1 ;
 RECT 0.945 3.13 1.085 3.22 ;
 RECT 0.565 3.22 1.085 3.47 ;
 RECT 0.945 3.47 1.085 3.725 ;
 RECT 1.905 3.365 2.045 3.505 ;
 RECT 1.905 3.645 2.045 3.71 ;
 RECT 1.905 3.105 2.215 3.365 ;
 RECT 1.905 3.505 3.145 3.645 ;
 RECT 3.005 3.645 3.145 4.345 ;
 END
END LSDNX1

MACRO XNOR2X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.45 1.4 4.59 2.565 ;
 RECT 4.45 1.16 4.76 1.4 ;
 RECT 4.45 0.515 4.59 1.16 ;
 END
 ANTENNADIFFAREA 0.702 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 0.665 1.55 0.805 2.8 ;
 RECT 2.09 1.825 2.23 2.8 ;
 RECT 4.94 2.12 5.08 2.8 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 3.88 2.12 4.02 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 4.945 0.08 5.085 0.82 ;
 RECT 2.075 0.08 2.215 0.82 ;
 RECT 0.665 0.08 0.805 0.775 ;
 RECT 3.9 0.08 4.04 0.82 ;
 RECT 0.215 0.08 0.355 0.755 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.27 1.16 3.465 1.32 ;
 RECT 3.27 1.32 3.64 1.58 ;
 END
 ANTENNAGATEAREA 0.136 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 0.985 1 1.4 ;
 END
 ANTENNAGATEAREA 0.136 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 0.92 2.44 2.47 2.535 ;
 RECT 0.92 2.535 2.465 2.54 ;
 RECT 2.37 0.395 2.47 2.44 ;
 RECT 0.92 1.215 1.02 2.44 ;
 RECT 0.92 0.375 1.02 0.985 ;
 RECT 0.815 0.985 1.025 1.215 ;
 RECT 3.28 0.425 3.38 0.975 ;
 RECT 3.16 0.21 3.39 0.425 ;
 RECT 3.665 0.39 3.765 2.425 ;
 RECT 3.56 2.425 3.77 2.655 ;
 RECT 3.28 1.42 3.38 2.535 ;
 RECT 1.785 0.215 1.885 2.255 ;
 RECT 2.77 0.215 2.87 1.155 ;
 RECT 2.77 1.19 3.485 1.255 ;
 RECT 3.275 1.255 3.485 1.42 ;
 RECT 2.77 1.155 3.38 1.19 ;
 RECT 1.785 0.115 2.87 0.215 ;
 RECT 2.775 1.65 2.875 2.53 ;
 RECT 2.66 1.435 2.89 1.65 ;
 RECT 4.17 0.35 4.27 1.07 ;
 RECT 4.17 1.285 4.27 2.745 ;
 RECT 4.045 1.07 4.275 1.08 ;
 RECT 4.045 1.08 4.825 1.18 ;
 RECT 4.045 1.18 4.275 1.285 ;
 RECT 4.725 0.35 4.825 1.08 ;
 RECT 4.725 1.18 4.825 2.745 ;
 LAYER CO ;
 RECT 2.095 1.875 2.225 2.005 ;
 RECT 3.21 0.25 3.34 0.38 ;
 RECT 4.455 2.385 4.585 2.515 ;
 RECT 0.67 0.595 0.8 0.725 ;
 RECT 3.315 1.24 3.445 1.37 ;
 RECT 4.095 1.11 4.225 1.24 ;
 RECT 4.455 0.625 4.585 0.755 ;
 RECT 2.995 2.115 3.125 2.245 ;
 RECT 3.885 2.17 4.015 2.3 ;
 RECT 0.855 1.035 0.985 1.165 ;
 RECT 0.67 1.62 0.8 1.75 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 2.995 1.81 3.125 1.94 ;
 RECT 4.945 2.17 5.075 2.3 ;
 RECT 3.905 0.625 4.035 0.755 ;
 RECT 3.6 2.475 3.73 2.605 ;
 RECT 2.08 0.625 2.21 0.755 ;
 RECT 4.455 1.835 4.585 1.965 ;
 RECT 4.455 2.11 4.585 2.24 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 1.535 0.625 1.665 0.755 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 1.145 1.6 1.275 1.73 ;
 RECT 2.71 1.475 2.84 1.605 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 1.535 1.81 1.665 1.94 ;
 RECT 4.95 0.625 5.08 0.755 ;
 RECT 1.145 0.595 1.275 0.725 ;
 RECT 4.455 1.56 4.585 1.69 ;
 RECT 2.995 0.625 3.125 0.755 ;
 LAYER M1 ;
 RECT 1.14 0.48 1.28 2.235 ;
 RECT 1.14 2.235 1.95 2.375 ;
 RECT 1.81 1.645 1.95 2.235 ;
 RECT 1.81 1.505 2.52 1.645 ;
 RECT 2.38 1.645 2.52 2.475 ;
 RECT 3.59 2.425 3.74 2.475 ;
 RECT 3.59 2.615 3.74 2.655 ;
 RECT 2.38 2.475 3.74 2.615 ;
 RECT 1.53 0.3 1.67 0.97 ;
 RECT 1.53 1.11 1.67 1.99 ;
 RECT 2.705 0.385 2.845 0.97 ;
 RECT 2.705 1.11 2.845 1.425 ;
 RECT 1.53 0.97 2.845 1.11 ;
 RECT 2.7 1.425 2.85 1.66 ;
 RECT 2.705 0.245 3.39 0.385 ;
 RECT 2.99 0.535 3.13 0.625 ;
 RECT 2.99 0.765 3.13 2.295 ;
 RECT 2.99 0.625 3.745 0.765 ;
 RECT 3.605 0.765 3.745 1.02 ;
 RECT 4.085 1.16 4.235 1.295 ;
 RECT 3.605 1.02 4.27 1.16 ;
 END
END XNOR2X2

MACRO XNOR3X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.68 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.2 2.375 7.5 2.66 ;
 RECT 7.36 0.44 7.5 2.375 ;
 END
 ANTENNADIFFAREA 0.468 ;
 END Q

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.04 1.075 5.445 1.4 ;
 END
 ANTENNAGATEAREA 0.129 ;
 END IN3

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.68 0.08 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 2.305 0.08 2.445 0.82 ;
 RECT 4.105 0.08 4.245 0.82 ;
 RECT 1.125 0.08 1.265 0.785 ;
 RECT 6.85 0.08 6.99 0.875 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 1.99 0.98 2.36 ;
 END
 ANTENNAGATEAREA 0.152 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.99 1.245 2.36 1.805 ;
 END
 ANTENNAGATEAREA 0.152 ;
 END IN1

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.68 2.96 ;
 RECT 6.89 1.73 7.03 2.8 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 2.18 2.35 2.32 2.8 ;
 RECT 1.125 1.515 1.265 2.8 ;
 RECT 4.11 1.89 4.25 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 5.01 1.215 6.64 1.305 ;
 RECT 5.01 1.075 5.29 1.215 ;
 RECT 5.19 0.335 5.29 1.075 ;
 RECT 5.19 1.305 6.64 1.315 ;
 RECT 6.54 0.385 6.64 1.215 ;
 RECT 6.54 1.315 6.64 2.1 ;
 RECT 5.66 1.315 5.76 2.415 ;
 RECT 5.14 1.5 5.24 2.595 ;
 RECT 6.26 2.35 6.36 2.595 ;
 RECT 5.14 2.595 6.36 2.695 ;
 RECT 6.15 2.12 6.36 2.35 ;
 RECT 3.535 1.4 3.635 2.78 ;
 RECT 2.975 0.945 3.08 0.985 ;
 RECT 2.975 0.985 3.075 1.3 ;
 RECT 2.98 0.2 3.08 0.945 ;
 RECT 1.965 0.2 2.065 1.365 ;
 RECT 1.965 1.365 2.18 1.595 ;
 RECT 1.965 1.595 2.065 2.5 ;
 RECT 2.975 1.3 3.635 1.4 ;
 RECT 1.965 0.1 3.08 0.2 ;
 RECT 3.77 0.39 3.99 0.465 ;
 RECT 3.89 0.465 3.99 2.78 ;
 RECT 3.77 0.235 3.98 0.39 ;
 RECT 3.485 0.21 3.585 0.89 ;
 RECT 3.47 0.89 3.68 1.12 ;
 RECT 4.365 0.385 4.465 1.175 ;
 RECT 4.365 1.39 4.465 2.39 ;
 RECT 4.25 1.175 4.48 1.39 ;
 RECT 2.575 0.395 2.675 2.68 ;
 RECT 0.905 0.355 1.005 2.075 ;
 RECT 0.905 2.305 1.005 2.68 ;
 RECT 0.905 2.68 2.675 2.78 ;
 RECT 0.805 2.075 1.015 2.305 ;
 RECT 5.655 0.39 5.76 0.44 ;
 RECT 5.655 0.21 5.755 0.39 ;
 RECT 5.66 0.44 5.76 0.905 ;
 RECT 5.655 0.205 6.355 0.21 ;
 RECT 5.655 0.11 6.35 0.205 ;
 RECT 6.145 0.21 6.355 0.475 ;
 RECT 7.145 0.24 7.245 1.185 ;
 RECT 6.99 1.185 7.245 1.395 ;
 RECT 7.145 1.395 7.245 2.78 ;
 RECT 2.98 1.83 3.08 2.78 ;
 RECT 2.87 1.6 3.08 1.83 ;
 LAYER CO ;
 RECT 3.51 0.94 3.64 1.07 ;
 RECT 7.365 1.555 7.495 1.685 ;
 RECT 0.845 2.125 0.975 2.255 ;
 RECT 0.655 0.605 0.785 0.735 ;
 RECT 0.655 1.525 0.785 1.655 ;
 RECT 7.365 1.91 7.495 2.04 ;
 RECT 4.115 2 4.245 2.13 ;
 RECT 3.81 0.285 3.94 0.415 ;
 RECT 6.185 0.295 6.315 0.425 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 2.01 1.415 2.14 1.545 ;
 RECT 4.11 0.625 4.24 0.755 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 6.855 0.645 6.985 0.775 ;
 RECT 7.365 0.49 7.495 0.62 ;
 RECT 1.13 0.605 1.26 0.735 ;
 RECT 4.915 0.625 5.045 0.755 ;
 RECT 3.2 0.625 3.33 0.755 ;
 RECT 5.055 1.125 5.185 1.255 ;
 RECT 1.13 1.59 1.26 1.72 ;
 RECT 1.715 0.625 1.845 0.755 ;
 RECT 2.91 1.65 3.04 1.78 ;
 RECT 6.29 1.555 6.42 1.685 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 2.185 2.42 2.315 2.55 ;
 RECT 5.88 2.025 6.01 2.155 ;
 RECT 5.41 0.625 5.54 0.755 ;
 RECT 6.19 2.17 6.32 2.3 ;
 RECT 5.88 0.625 6.01 0.755 ;
 RECT 6.29 0.64 6.42 0.77 ;
 RECT 3.2 2.05 3.33 2.18 ;
 RECT 4.3 1.215 4.43 1.345 ;
 RECT 4.765 1.95 4.895 2.08 ;
 RECT 7.04 1.225 7.17 1.355 ;
 RECT 1.715 2.07 1.845 2.2 ;
 RECT 6.895 1.855 7.025 1.985 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 2.31 0.625 2.44 0.755 ;
 RECT 5.41 1.915 5.54 2.045 ;
 LAYER M1 ;
 RECT 4.76 0.76 4.9 2.15 ;
 RECT 4.76 0.62 5.1 0.76 ;
 RECT 5.405 1.805 5.545 2.49 ;
 RECT 5.405 2.49 6.73 2.63 ;
 RECT 5.405 2.63 5.545 2.635 ;
 RECT 5.36 0.62 5.725 0.76 ;
 RECT 5.585 0.76 5.725 1.665 ;
 RECT 5.405 1.665 5.725 1.805 ;
 RECT 6.59 1.355 6.73 2.49 ;
 RECT 6.99 1.355 7.22 1.365 ;
 RECT 6.59 1.215 7.22 1.355 ;
 RECT 3.195 0.575 3.335 0.605 ;
 RECT 3.195 0.745 3.335 2.265 ;
 RECT 3.185 0.605 3.965 0.745 ;
 RECT 3.825 0.745 3.965 1.205 ;
 RECT 4.29 1.165 4.61 1.205 ;
 RECT 4.47 0.395 4.61 1.165 ;
 RECT 4.29 1.35 4.48 1.4 ;
 RECT 4.29 1.345 4.61 1.35 ;
 RECT 3.825 1.205 4.61 1.345 ;
 RECT 5.875 0.395 6.015 2.21 ;
 RECT 4.47 0.255 6.015 0.395 ;
 RECT 1.71 0.515 1.85 2.025 ;
 RECT 1.71 2.165 1.85 2.295 ;
 RECT 2.52 1.61 2.66 2.025 ;
 RECT 2.52 2.165 2.66 2.415 ;
 RECT 2.905 1.61 3.045 1.835 ;
 RECT 1.71 2.025 2.66 2.165 ;
 RECT 3.475 1.12 3.615 2.415 ;
 RECT 3.475 0.89 3.65 1.12 ;
 RECT 2.52 1.47 3.055 1.61 ;
 RECT 2.52 2.415 3.62 2.555 ;
 RECT 0.65 0.51 0.79 1.06 ;
 RECT 0.65 1.2 0.79 1.775 ;
 RECT 0.65 1.06 1.56 1.2 ;
 RECT 1.42 0.365 1.56 1.06 ;
 RECT 1.42 0.225 2.13 0.365 ;
 RECT 1.99 0.365 2.13 0.965 ;
 RECT 3.8 0.235 3.95 0.265 ;
 RECT 3.8 0.405 3.95 0.465 ;
 RECT 2.62 0.265 3.95 0.405 ;
 RECT 1.99 0.965 2.76 1.105 ;
 RECT 2.62 0.405 2.76 0.965 ;
 RECT 6.175 0.245 6.425 0.475 ;
 RECT 6.285 0.475 6.425 2.12 ;
 RECT 6.18 2.12 6.425 2.35 ;
 RECT 6.185 0.22 6.425 0.245 ;
 END
END XNOR3X1

MACRO XNOR3X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.32 BY 2.88 ;
 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.05 1.365 2.36 1.72 ;
 END
 ANTENNAGATEAREA 0.152 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.04 1.075 5.445 1.4 ;
 END
 ANTENNAGATEAREA 0.128 ;
 END IN3

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.36 1.16 7.64 1.4 ;
 RECT 7.36 1.4 7.5 2.655 ;
 RECT 7.36 0.535 7.5 1.16 ;
 END
 ANTENNADIFFAREA 0.64 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.32 2.96 ;
 RECT 4.11 1.89 4.25 2.8 ;
 RECT 1.125 1.515 1.265 2.8 ;
 RECT 6.89 1.73 7.03 2.8 ;
 RECT 2.18 2.35 2.32 2.8 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 7.865 1.73 8.005 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.32 0.08 ;
 RECT 4.105 0.08 4.245 0.82 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 6.85 0.08 6.99 0.875 ;
 RECT 2.305 0.08 2.445 0.82 ;
 RECT 1.125 0.08 1.265 0.785 ;
 RECT 7.86 0.08 8 0.875 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 2.075 0.98 2.36 ;
 END
 ANTENNAGATEAREA 0.152 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 5.01 1.215 6.64 1.305 ;
 RECT 5.01 1.075 5.29 1.215 ;
 RECT 5.19 0.335 5.29 1.075 ;
 RECT 5.19 1.305 6.64 1.315 ;
 RECT 6.54 0.385 6.64 1.215 ;
 RECT 6.54 1.315 6.64 2.1 ;
 RECT 5.66 1.315 5.76 2.45 ;
 RECT 1.965 0.2 2.065 1.365 ;
 RECT 1.965 1.365 2.265 1.595 ;
 RECT 1.965 1.595 2.065 2.5 ;
 RECT 3.535 1.4 3.635 2.78 ;
 RECT 2.975 0.945 3.08 0.985 ;
 RECT 2.975 0.985 3.075 1.3 ;
 RECT 2.98 0.2 3.08 0.945 ;
 RECT 2.975 1.3 3.635 1.4 ;
 RECT 1.965 0.1 3.08 0.2 ;
 RECT 6.99 1.185 7.245 1.25 ;
 RECT 6.99 1.35 7.245 1.395 ;
 RECT 6.99 1.25 7.74 1.35 ;
 RECT 7.64 0.19 7.74 1.25 ;
 RECT 7.64 1.35 7.74 2.78 ;
 RECT 7.145 0.195 7.245 1.185 ;
 RECT 7.145 1.395 7.245 2.78 ;
 RECT 3.77 0.39 3.99 0.465 ;
 RECT 3.89 0.465 3.99 2.78 ;
 RECT 3.77 0.235 3.98 0.39 ;
 RECT 5.14 1.5 5.24 2.635 ;
 RECT 6.26 2.35 6.36 2.635 ;
 RECT 5.14 2.635 6.36 2.735 ;
 RECT 6.15 2.12 6.36 2.35 ;
 RECT 5.655 0.39 5.76 0.44 ;
 RECT 5.655 0.21 5.755 0.39 ;
 RECT 5.66 0.44 5.76 0.905 ;
 RECT 5.655 0.205 6.355 0.21 ;
 RECT 5.655 0.11 6.35 0.205 ;
 RECT 6.145 0.21 6.355 0.475 ;
 RECT 0.905 0.355 1.005 2.075 ;
 RECT 0.905 2.305 1.005 2.68 ;
 RECT 2.575 0.395 2.675 2.68 ;
 RECT 0.805 2.075 1.015 2.305 ;
 RECT 0.905 2.68 2.675 2.78 ;
 RECT 2.98 1.83 3.08 2.78 ;
 RECT 2.87 1.6 3.08 1.83 ;
 RECT 3.485 0.21 3.585 0.89 ;
 RECT 3.47 0.89 3.68 1.12 ;
 RECT 4.365 0.385 4.465 1.175 ;
 RECT 4.365 1.39 4.465 2.465 ;
 RECT 4.25 1.175 4.48 1.39 ;
 LAYER CO ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 6.19 2.17 6.32 2.3 ;
 RECT 5.41 1.915 5.54 2.045 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 3.51 0.94 3.64 1.07 ;
 RECT 3.81 0.285 3.94 0.415 ;
 RECT 5.88 0.625 6.01 0.755 ;
 RECT 0.845 2.125 0.975 2.255 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 6.855 0.645 6.985 0.775 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 7.365 1.555 7.495 1.685 ;
 RECT 4.11 0.625 4.24 0.755 ;
 RECT 6.29 0.64 6.42 0.77 ;
 RECT 7.365 0.675 7.495 0.805 ;
 RECT 2.31 0.625 2.44 0.755 ;
 RECT 5.055 1.125 5.185 1.255 ;
 RECT 1.715 0.625 1.845 0.755 ;
 RECT 4.765 2.01 4.895 2.14 ;
 RECT 0.655 0.605 0.785 0.735 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 3.2 2.05 3.33 2.18 ;
 RECT 2.185 2.42 2.315 2.55 ;
 RECT 6.185 0.295 6.315 0.425 ;
 RECT 5.41 0.625 5.54 0.755 ;
 RECT 6.895 1.855 7.025 1.985 ;
 RECT 6.29 1.555 6.42 1.685 ;
 RECT 2.095 1.415 2.225 1.545 ;
 RECT 2.91 1.65 3.04 1.78 ;
 RECT 1.715 2.07 1.845 2.2 ;
 RECT 7.04 1.225 7.17 1.355 ;
 RECT 1.13 0.605 1.26 0.735 ;
 RECT 7.365 2.425 7.495 2.555 ;
 RECT 7.365 2.13 7.495 2.26 ;
 RECT 6.895 2.385 7.025 2.515 ;
 RECT 6.895 2.12 7.025 2.25 ;
 RECT 7.87 2.38 8 2.51 ;
 RECT 7.87 2.115 8 2.245 ;
 RECT 7.865 0.645 7.995 0.775 ;
 RECT 7.87 1.855 8 1.985 ;
 RECT 3.2 0.625 3.33 0.755 ;
 RECT 4.115 2 4.245 2.13 ;
 RECT 7.365 1.815 7.495 1.945 ;
 RECT 4.915 0.625 5.045 0.755 ;
 RECT 0.655 1.525 0.785 1.655 ;
 RECT 1.13 1.59 1.26 1.72 ;
 RECT 4.3 1.215 4.43 1.345 ;
 RECT 5.88 2.025 6.01 2.155 ;
 LAYER M1 ;
 RECT 4.76 0.76 4.9 2.265 ;
 RECT 4.76 0.62 5.1 0.76 ;
 RECT 1.71 0.515 1.85 2.025 ;
 RECT 1.71 2.165 1.85 2.295 ;
 RECT 2.52 1.61 2.66 2.025 ;
 RECT 2.52 2.165 2.66 2.415 ;
 RECT 2.905 1.61 3.045 1.835 ;
 RECT 1.71 2.025 2.66 2.165 ;
 RECT 3.475 1.12 3.615 2.415 ;
 RECT 3.475 0.89 3.65 1.12 ;
 RECT 2.52 1.47 3.055 1.61 ;
 RECT 2.52 2.415 3.62 2.555 ;
 RECT 0.65 1.06 1.56 1.2 ;
 RECT 1.42 0.365 1.56 1.06 ;
 RECT 0.65 0.51 0.79 1.06 ;
 RECT 0.65 1.2 0.79 1.775 ;
 RECT 1.42 0.225 2.13 0.365 ;
 RECT 1.99 0.365 2.13 0.965 ;
 RECT 3.8 0.235 3.95 0.265 ;
 RECT 3.8 0.405 3.95 0.465 ;
 RECT 2.62 0.265 3.95 0.405 ;
 RECT 1.99 0.965 2.76 1.105 ;
 RECT 2.62 0.405 2.76 0.965 ;
 RECT 3.195 0.575 3.335 0.605 ;
 RECT 3.195 0.745 3.335 2.265 ;
 RECT 3.185 0.605 3.965 0.745 ;
 RECT 3.825 0.745 3.965 1.205 ;
 RECT 4.29 1.165 4.61 1.205 ;
 RECT 4.47 0.395 4.61 1.165 ;
 RECT 4.29 1.35 4.48 1.4 ;
 RECT 4.29 1.345 4.61 1.35 ;
 RECT 3.825 1.205 4.61 1.345 ;
 RECT 5.875 0.395 6.015 2.21 ;
 RECT 4.47 0.255 6.015 0.395 ;
 RECT 5.405 1.805 5.545 2.49 ;
 RECT 5.405 2.49 6.73 2.63 ;
 RECT 5.405 2.63 5.545 2.635 ;
 RECT 5.36 0.62 5.725 0.76 ;
 RECT 5.585 0.76 5.725 1.665 ;
 RECT 5.405 1.665 5.725 1.805 ;
 RECT 6.59 1.355 6.73 2.49 ;
 RECT 6.99 1.355 7.22 1.365 ;
 RECT 6.59 1.215 7.22 1.355 ;
 RECT 6.175 0.245 6.425 0.475 ;
 RECT 6.285 0.475 6.425 2.12 ;
 RECT 6.18 2.12 6.425 2.35 ;
 RECT 6.185 0.22 6.425 0.245 ;
 END
END XNOR3X2

MACRO XOR2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 4.8 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 4.8 2.96 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 4.375 1.515 4.515 2.8 ;
 RECT 1.115 1.825 1.255 2.8 ;
 RECT 2.92 2.12 3.06 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 4.8 0.08 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 4.375 0.08 4.515 0.785 ;
 RECT 1.115 0.08 1.255 0.82 ;
 RECT 2.94 0.08 3.08 0.82 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.195 1 4.44 1.365 ;
 END
 ANTENNAGATEAREA 0.134 ;
 END IN2

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.4 0.36 3.64 0.6 ;
 RECT 3.49 0.6 3.63 1.745 ;
 END
 ANTENNADIFFAREA 0.56 ;
 END Q

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.32 1.265 2.68 1.56 ;
 END
 ANTENNAGATEAREA 0.134 ;
 END IN1

 OBS
 LAYER PO ;
 RECT 3.21 0.38 3.31 1.175 ;
 RECT 3.21 1.39 3.31 2.77 ;
 RECT 3.085 1.175 3.315 1.39 ;
 RECT 2.32 0.425 2.42 0.975 ;
 RECT 2.2 0.21 2.43 0.425 ;
 RECT 1.815 1.665 1.915 2.53 ;
 RECT 1.7 1.45 1.93 1.665 ;
 RECT 1.41 0.395 1.51 2.425 ;
 RECT 1.37 2.425 1.58 2.655 ;
 RECT 2.32 1.56 2.42 2.53 ;
 RECT 1.81 0.195 1.91 1.165 ;
 RECT 0.9 0.195 1 2.255 ;
 RECT 2.31 1.265 2.52 1.56 ;
 RECT 1.81 1.165 2.42 1.265 ;
 RECT 0.9 0.095 1.91 0.195 ;
 RECT 2.705 0.2 2.805 2.545 ;
 RECT 4.155 0.2 4.255 1 ;
 RECT 4.155 1.23 4.255 1.945 ;
 RECT 4.155 1 4.43 1.23 ;
 RECT 2.705 0.1 4.255 0.2 ;
 LAYER CO ;
 RECT 3.135 1.215 3.265 1.345 ;
 RECT 4.26 1.05 4.39 1.18 ;
 RECT 2.35 1.38 2.48 1.51 ;
 RECT 1.41 2.475 1.54 2.605 ;
 RECT 2.25 0.25 2.38 0.38 ;
 RECT 1.75 1.49 1.88 1.62 ;
 RECT 3.495 0.625 3.625 0.755 ;
 RECT 3.495 1.56 3.625 1.69 ;
 RECT 2.945 0.625 3.075 0.755 ;
 RECT 2.925 2.17 3.055 2.3 ;
 RECT 2.035 2.115 2.165 2.245 ;
 RECT 2.035 1.81 2.165 1.94 ;
 RECT 2.035 0.625 2.165 0.755 ;
 RECT 1.12 0.625 1.25 0.755 ;
 RECT 1.12 1.875 1.25 2.005 ;
 RECT 0.65 1.81 0.78 1.94 ;
 RECT 0.65 0.625 0.78 0.755 ;
 RECT 4.38 0.605 4.51 0.735 ;
 RECT 3.905 0.605 4.035 0.735 ;
 RECT 4.38 1.59 4.51 1.72 ;
 RECT 3.905 1.525 4.035 1.655 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 0.205 2.065 0.335 2.195 ;
 LAYER M1 ;
 RECT 2.03 0.535 2.17 0.625 ;
 RECT 2.03 0.765 2.17 2.295 ;
 RECT 2.03 0.625 2.8 0.765 ;
 RECT 2.66 0.765 2.8 0.97 ;
 RECT 3.085 1.11 3.315 1.4 ;
 RECT 2.66 0.97 3.315 1.11 ;
 RECT 1.4 2.425 1.55 2.46 ;
 RECT 1.4 2.6 1.55 2.655 ;
 RECT 1.4 2.46 2.61 2.6 ;
 RECT 2.47 1.97 2.61 2.46 ;
 RECT 2.47 1.83 3.35 1.925 ;
 RECT 3.9 0.49 4.04 1.925 ;
 RECT 3.21 1.97 4.04 2.065 ;
 RECT 2.47 1.925 4.04 1.97 ;
 RECT 0.645 0.3 0.785 1.52 ;
 RECT 0.645 1.66 0.785 1.99 ;
 RECT 1.46 0.385 1.6 1.52 ;
 RECT 1.46 1.66 1.6 1.665 ;
 RECT 0.645 1.52 1.89 1.66 ;
 RECT 1.74 1.44 1.89 1.52 ;
 RECT 1.74 1.66 1.89 1.675 ;
 RECT 1.46 0.245 2.43 0.385 ;
 END
END XOR2X1

MACRO XOR2X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.49 1.4 3.63 1.745 ;
 RECT 3.49 1.16 3.8 1.4 ;
 RECT 3.49 0.515 3.63 1.16 ;
 END
 ANTENNADIFFAREA 0.7 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 1.115 1.825 1.255 2.8 ;
 RECT 2.92 2.12 3.06 2.8 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 4.005 2.27 4.145 2.8 ;
 RECT 4.895 1.515 5.035 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 4.895 0.08 5.035 0.785 ;
 RECT 1.115 0.08 1.255 0.82 ;
 RECT 2.94 0.08 3.08 0.82 ;
 RECT 4 0.08 4.14 0.82 ;
 END
 END VSS

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.325 1.32 2.68 1.56 ;
 RECT 2.325 1.56 2.495 1.65 ;
 RECT 2.325 1.16 2.495 1.32 ;
 END
 ANTENNAGATEAREA 0.134 ;
 END IN1

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.765 0.98 5.12 1.375 ;
 END
 ANTENNAGATEAREA 0.134 ;
 END IN2

 OBS
 LAYER PO ;
 RECT 2.32 0.425 2.42 0.975 ;
 RECT 2.2 0.21 2.43 0.425 ;
 RECT 2.32 1.42 2.42 2.53 ;
 RECT 0.9 0.215 1 2.255 ;
 RECT 1.81 0.215 1.91 1.165 ;
 RECT 1.81 1.19 2.525 1.265 ;
 RECT 2.315 1.265 2.525 1.42 ;
 RECT 1.81 1.165 2.42 1.19 ;
 RECT 0.9 0.115 1.91 0.215 ;
 RECT 1.815 1.665 1.915 2.53 ;
 RECT 1.7 1.45 1.93 1.665 ;
 RECT 3.77 1.225 3.87 2.77 ;
 RECT 3.21 0.375 3.31 1.125 ;
 RECT 3.21 1.125 3.87 1.175 ;
 RECT 3.77 0.375 3.87 1.125 ;
 RECT 3.085 1.175 3.87 1.225 ;
 RECT 3.085 1.225 3.315 1.39 ;
 RECT 3.21 1.39 3.31 2.77 ;
 RECT 1.41 0.395 1.51 2.425 ;
 RECT 1.37 2.425 1.58 2.655 ;
 RECT 2.705 0.195 2.805 2.545 ;
 RECT 4.675 0.195 4.775 1 ;
 RECT 4.675 1.23 4.775 1.945 ;
 RECT 4.675 1 4.95 1.23 ;
 RECT 2.705 0.095 4.775 0.195 ;
 LAYER CO ;
 RECT 1.12 1.875 1.25 2.005 ;
 RECT 2.035 1.81 2.165 1.94 ;
 RECT 2.945 0.625 3.075 0.755 ;
 RECT 4.9 0.605 5.03 0.735 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 4.005 0.625 4.135 0.755 ;
 RECT 4.01 2.375 4.14 2.505 ;
 RECT 2.355 1.24 2.485 1.37 ;
 RECT 4.78 1.05 4.91 1.18 ;
 RECT 1.75 1.49 1.88 1.62 ;
 RECT 2.25 0.25 2.38 0.38 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 2.925 2.17 3.055 2.3 ;
 RECT 3.495 0.625 3.625 0.755 ;
 RECT 1.12 0.625 1.25 0.755 ;
 RECT 4.9 1.59 5.03 1.72 ;
 RECT 0.65 0.625 0.78 0.755 ;
 RECT 3.135 1.215 3.265 1.345 ;
 RECT 2.035 0.625 2.165 0.755 ;
 RECT 4.425 1.525 4.555 1.655 ;
 RECT 4.425 0.605 4.555 0.735 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 3.495 1.56 3.625 1.69 ;
 RECT 0.65 1.81 0.78 1.94 ;
 RECT 1.41 2.475 1.54 2.605 ;
 RECT 2.035 2.115 2.165 2.245 ;
 RECT 0.205 1.545 0.335 1.675 ;
 LAYER M1 ;
 RECT 2.47 1.83 3.35 1.925 ;
 RECT 1.4 2.425 1.55 2.46 ;
 RECT 1.4 2.6 1.55 2.655 ;
 RECT 1.4 2.46 2.61 2.6 ;
 RECT 2.47 1.97 2.61 2.46 ;
 RECT 4.415 1.66 4.56 1.775 ;
 RECT 4.415 1.775 4.555 1.925 ;
 RECT 4.42 0.49 4.56 1.66 ;
 RECT 3.21 1.97 4.555 2.065 ;
 RECT 2.47 1.925 4.555 1.97 ;
 RECT 0.645 0.415 0.785 1.52 ;
 RECT 0.645 1.66 0.785 1.99 ;
 RECT 0.645 1.52 1.89 1.66 ;
 RECT 1.46 0.385 1.6 1.52 ;
 RECT 1.46 1.66 1.6 1.665 ;
 RECT 1.74 1.44 1.89 1.52 ;
 RECT 1.74 1.66 1.89 1.675 ;
 RECT 1.46 0.245 2.43 0.385 ;
 RECT 2.03 0.535 2.17 0.625 ;
 RECT 2.03 0.765 2.17 2.295 ;
 RECT 2.03 0.625 2.785 0.765 ;
 RECT 2.645 0.765 2.785 0.96 ;
 RECT 3.11 1.1 3.275 1.405 ;
 RECT 2.645 0.96 3.275 1.1 ;
 END
END XOR2X2

MACRO XOR3X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 7.68 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.345 1.11 7.595 1.4 ;
 RECT 7.36 1.4 7.5 2.62 ;
 RECT 7.36 0.49 7.5 1.11 ;
 END
 ANTENNADIFFAREA 0.468 ;
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 7.68 2.96 ;
 RECT 2.18 2.35 2.32 2.8 ;
 RECT 1.125 1.515 1.265 2.8 ;
 RECT 4.11 1.89 4.25 2.8 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 6.89 1.46 7.03 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 7.68 0.08 ;
 RECT 4.105 0.08 4.245 0.82 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 1.125 0.08 1.265 0.785 ;
 RECT 2.305 0.08 2.445 0.82 ;
 RECT 6.85 0.08 6.99 0.875 ;
 END
 END VSS

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.625 2.07 0.98 2.315 ;
 END
 ANTENNAGATEAREA 0.152 ;
 END IN2

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2 1.365 2.305 1.72 ;
 END
 ANTENNAGATEAREA 0.152 ;
 END IN1

 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.04 1.11 5.4 1.425 ;
 END
 ANTENNAGATEAREA 0.129 ;
 END IN3

 OBS
 LAYER PO ;
 RECT 7.145 0.24 7.245 1.115 ;
 RECT 7.145 1.325 7.245 2.76 ;
 RECT 6.945 1.115 7.245 1.325 ;
 RECT 0.905 0.355 1.005 2.075 ;
 RECT 0.905 2.305 1.005 2.68 ;
 RECT 2.575 0.395 2.675 2.68 ;
 RECT 0.805 2.075 1.015 2.305 ;
 RECT 0.905 2.68 2.675 2.78 ;
 RECT 2.98 1.83 3.08 2.78 ;
 RECT 2.87 1.6 3.08 1.83 ;
 RECT 4.365 0.385 4.465 1.175 ;
 RECT 4.365 1.39 4.465 2.39 ;
 RECT 4.25 1.175 4.48 1.39 ;
 RECT 3.77 0.39 3.99 0.465 ;
 RECT 3.89 0.465 3.99 2.78 ;
 RECT 3.77 0.235 3.98 0.39 ;
 RECT 3.485 0.21 3.585 0.89 ;
 RECT 3.47 0.89 3.68 1.12 ;
 RECT 5.19 0.21 5.29 0.935 ;
 RECT 5.19 0.205 6.355 0.21 ;
 RECT 5.19 0.11 6.35 0.205 ;
 RECT 6.145 0.21 6.355 0.475 ;
 RECT 5.045 1.235 6.64 1.31 ;
 RECT 5.505 1.31 6.64 1.315 ;
 RECT 5.14 1.215 6.64 1.235 ;
 RECT 5.14 1.21 5.76 1.215 ;
 RECT 6.54 0.385 6.64 1.215 ;
 RECT 6.54 1.315 6.64 2.1 ;
 RECT 5.66 0.39 5.76 1.21 ;
 RECT 5.14 1.465 5.24 2.43 ;
 RECT 5.045 1.31 5.26 1.465 ;
 RECT 5.66 2.31 6.36 2.32 ;
 RECT 5.66 1.495 5.76 2.31 ;
 RECT 5.66 2.41 5.76 2.415 ;
 RECT 5.66 2.32 6.285 2.41 ;
 RECT 6.15 2.09 6.36 2.31 ;
 RECT 3.535 1.4 3.635 2.78 ;
 RECT 2.975 0.945 3.08 0.985 ;
 RECT 2.975 0.985 3.075 1.3 ;
 RECT 2.98 0.2 3.08 0.945 ;
 RECT 1.965 0.2 2.065 1.365 ;
 RECT 1.965 1.365 2.18 1.595 ;
 RECT 1.965 1.595 2.065 2.5 ;
 RECT 2.975 1.3 3.635 1.4 ;
 RECT 1.965 0.1 3.08 0.2 ;
 LAYER CO ;
 RECT 5.88 2.025 6.01 2.155 ;
 RECT 5.41 0.625 5.54 0.755 ;
 RECT 5.41 1.915 5.54 2.045 ;
 RECT 2.91 1.65 3.04 1.78 ;
 RECT 3.81 0.285 3.94 0.415 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 2.185 2.42 2.315 2.55 ;
 RECT 2.31 0.625 2.44 0.755 ;
 RECT 1.715 0.625 1.845 0.755 ;
 RECT 3.2 2.05 3.33 2.18 ;
 RECT 0.655 0.605 0.785 0.735 ;
 RECT 4.915 0.625 5.045 0.755 ;
 RECT 4.11 0.625 4.24 0.755 ;
 RECT 4.3 1.215 4.43 1.345 ;
 RECT 1.13 0.605 1.26 0.735 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 3.2 0.625 3.33 0.755 ;
 RECT 0.655 1.525 0.785 1.655 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 4.765 2.035 4.895 2.165 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 0.845 2.125 0.975 2.255 ;
 RECT 1.715 2.07 1.845 2.2 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 4.115 2 4.245 2.13 ;
 RECT 1.13 1.59 1.26 1.72 ;
 RECT 5.88 1.76 6.01 1.89 ;
 RECT 6.895 1.55 7.025 1.68 ;
 RECT 6.895 2.15 7.025 2.28 ;
 RECT 7.365 2.165 7.495 2.295 ;
 RECT 3.51 0.94 3.64 1.07 ;
 RECT 5.09 1.285 5.22 1.415 ;
 RECT 6.19 2.14 6.32 2.27 ;
 RECT 2.01 1.415 2.14 1.545 ;
 RECT 6.185 0.295 6.315 0.425 ;
 RECT 6.995 1.155 7.125 1.285 ;
 RECT 7.365 1.88 7.495 2.01 ;
 RECT 7.365 0.6 7.495 0.73 ;
 RECT 7.365 1.525 7.495 1.655 ;
 RECT 6.855 0.645 6.985 0.775 ;
 RECT 6.895 1.825 7.025 1.955 ;
 RECT 6.29 0.64 6.42 0.77 ;
 RECT 6.29 1.525 6.42 1.655 ;
 RECT 5.88 0.625 6.01 0.755 ;
 LAYER M1 ;
 RECT 4.76 0.76 4.9 2.235 ;
 RECT 4.76 0.62 5.1 0.76 ;
 RECT 5.405 2.49 6.73 2.615 ;
 RECT 5.415 2.615 6.73 2.63 ;
 RECT 5.405 1.87 5.545 2.49 ;
 RECT 5.36 0.62 5.68 0.76 ;
 RECT 5.54 0.76 5.68 1.73 ;
 RECT 5.405 1.73 5.68 1.87 ;
 RECT 6.59 1.3 6.73 2.49 ;
 RECT 6.945 1.145 7.175 1.16 ;
 RECT 6.59 1.16 7.18 1.3 ;
 RECT 3.195 0.575 3.335 0.605 ;
 RECT 3.195 0.745 3.335 2.265 ;
 RECT 3.185 0.605 3.965 0.745 ;
 RECT 3.825 0.745 3.965 1.205 ;
 RECT 4.29 1.165 4.61 1.205 ;
 RECT 4.47 0.395 4.61 1.165 ;
 RECT 4.29 1.35 4.48 1.4 ;
 RECT 4.29 1.345 4.61 1.35 ;
 RECT 3.825 1.205 4.61 1.345 ;
 RECT 5.875 0.395 6.015 2.21 ;
 RECT 4.47 0.255 6.015 0.395 ;
 RECT 0.65 0.51 0.79 1.06 ;
 RECT 0.65 1.2 0.79 1.775 ;
 RECT 0.65 1.06 1.56 1.2 ;
 RECT 1.42 0.365 1.56 1.06 ;
 RECT 1.42 0.225 2.13 0.365 ;
 RECT 1.99 0.365 2.13 0.965 ;
 RECT 3.8 0.235 3.95 0.265 ;
 RECT 3.8 0.405 3.95 0.465 ;
 RECT 2.62 0.265 3.95 0.405 ;
 RECT 1.99 0.965 2.76 1.105 ;
 RECT 2.62 0.405 2.76 0.965 ;
 RECT 1.71 0.515 1.85 2.025 ;
 RECT 1.71 2.165 1.85 2.295 ;
 RECT 2.52 1.775 2.66 2.025 ;
 RECT 2.52 2.165 2.66 2.415 ;
 RECT 2.905 1.585 3.045 1.635 ;
 RECT 2.905 1.775 3.045 1.835 ;
 RECT 1.71 2.025 2.66 2.165 ;
 RECT 3.475 1.12 3.615 2.415 ;
 RECT 3.475 0.89 3.65 1.12 ;
 RECT 2.52 1.635 3.055 1.775 ;
 RECT 2.52 2.415 3.62 2.555 ;
 RECT 6.175 0.245 6.425 0.475 ;
 RECT 6.285 0.475 6.425 2.09 ;
 RECT 6.185 0.22 6.425 0.245 ;
 RECT 6.18 2.09 6.425 2.32 ;
 END
END XOR3X1

MACRO XOR3X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.32 BY 2.88 ;
 PIN IN3
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.04 1.16 5.4 1.425 ;
 END
 ANTENNAGATEAREA 0.128 ;
 END IN3

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.32 2.96 ;
 RECT 4.11 1.89 4.25 2.8 ;
 RECT 6.89 1.46 7.03 2.8 ;
 RECT 1.125 1.515 1.265 2.8 ;
 RECT 0.2 1.495 0.34 2.8 ;
 RECT 2.18 2.35 2.32 2.8 ;
 RECT 7.83 1.46 7.97 2.8 ;
 END
 END VDD

 PIN IN1
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.99 1.32 2.36 1.72 ;
 END
 ANTENNAGATEAREA 0.152 ;
 END IN1

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.36 1.4 7.5 2.62 ;
 RECT 7.36 1.16 7.64 1.4 ;
 RECT 7.36 0.49 7.5 1.16 ;
 END
 ANTENNADIFFAREA 0.6 ;
 END Q

 PIN IN2
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.68 2.075 0.98 2.36 ;
 END
 ANTENNAGATEAREA 0.152 ;
 END IN2

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.32 0.08 ;
 RECT 4.105 0.08 4.245 0.82 ;
 RECT 0.215 0.08 0.355 0.755 ;
 RECT 2.305 0.08 2.445 0.82 ;
 RECT 6.85 0.08 6.99 0.875 ;
 RECT 1.125 0.08 1.265 0.785 ;
 RECT 7.83 0.08 7.97 0.875 ;
 END
 END VSS

 OBS
 LAYER PO ;
 RECT 3.485 0.21 3.585 0.89 ;
 RECT 3.47 0.89 3.68 1.12 ;
 RECT 6.15 2.32 6.285 2.335 ;
 RECT 5.66 2.335 6.285 2.43 ;
 RECT 5.665 2.43 6.285 2.435 ;
 RECT 5.66 1.465 5.76 2.335 ;
 RECT 6.15 2.09 6.36 2.32 ;
 RECT 3.77 0.39 3.99 0.465 ;
 RECT 3.89 0.465 3.99 2.78 ;
 RECT 3.77 0.235 3.98 0.39 ;
 RECT 5.19 0.21 5.29 0.935 ;
 RECT 5.19 0.205 6.355 0.21 ;
 RECT 5.19 0.11 6.35 0.205 ;
 RECT 6.145 0.21 6.355 0.475 ;
 RECT 4.365 0.385 4.465 1.175 ;
 RECT 4.365 1.39 4.465 2.42 ;
 RECT 4.25 1.175 4.48 1.39 ;
 RECT 2.575 0.395 2.675 2.68 ;
 RECT 0.905 0.355 1.005 2.075 ;
 RECT 0.905 2.305 1.005 2.68 ;
 RECT 0.905 2.68 2.675 2.78 ;
 RECT 0.805 2.075 1.015 2.305 ;
 RECT 6.99 1.115 7.245 1.16 ;
 RECT 6.99 1.16 7.715 1.26 ;
 RECT 6.99 1.26 7.245 1.325 ;
 RECT 7.615 0.175 7.715 1.16 ;
 RECT 7.615 1.26 7.715 2.785 ;
 RECT 7.145 0.18 7.245 1.115 ;
 RECT 7.145 1.325 7.245 2.785 ;
 RECT 2.98 1.83 3.08 2.78 ;
 RECT 2.87 1.6 3.08 1.83 ;
 RECT 1.965 0.2 2.065 1.365 ;
 RECT 1.965 1.365 2.18 1.595 ;
 RECT 1.965 1.595 2.065 2.5 ;
 RECT 2.98 0.2 3.08 0.945 ;
 RECT 2.975 0.945 3.08 0.985 ;
 RECT 2.975 0.985 3.075 1.3 ;
 RECT 3.535 1.4 3.635 2.78 ;
 RECT 1.965 0.1 3.08 0.2 ;
 RECT 2.975 1.3 3.635 1.4 ;
 RECT 5.045 1.235 6.64 1.285 ;
 RECT 5.14 1.465 5.24 2.43 ;
 RECT 5.14 1.185 6.64 1.235 ;
 RECT 5.66 0.39 5.76 1.185 ;
 RECT 5.045 1.285 5.26 1.465 ;
 RECT 6.54 0.385 6.64 1.185 ;
 RECT 6.54 1.285 6.64 2.1 ;
 LAYER CO ;
 RECT 2.01 1.415 2.14 1.545 ;
 RECT 5.88 1.76 6.01 1.89 ;
 RECT 6.895 2.15 7.025 2.28 ;
 RECT 6.29 1.525 6.42 1.655 ;
 RECT 0.655 1.525 0.785 1.655 ;
 RECT 6.895 1.55 7.025 1.68 ;
 RECT 3.2 0.625 3.33 0.755 ;
 RECT 1.715 0.625 1.845 0.755 ;
 RECT 3.51 0.94 3.64 1.07 ;
 RECT 0.655 0.605 0.785 0.735 ;
 RECT 6.29 0.64 6.42 0.77 ;
 RECT 7.365 2.165 7.495 2.295 ;
 RECT 6.855 0.645 6.985 0.775 ;
 RECT 7.04 1.155 7.17 1.285 ;
 RECT 0.205 2.065 0.335 2.195 ;
 RECT 2.185 2.42 2.315 2.55 ;
 RECT 1.715 2.07 1.845 2.2 ;
 RECT 2.31 0.625 2.44 0.755 ;
 RECT 0.22 0.575 0.35 0.705 ;
 RECT 5.41 1.915 5.54 2.045 ;
 RECT 6.895 1.825 7.025 1.955 ;
 RECT 6.19 2.14 6.32 2.27 ;
 RECT 0.22 0.315 0.35 0.445 ;
 RECT 5.88 0.625 6.01 0.755 ;
 RECT 3.2 2.05 3.33 2.18 ;
 RECT 0.205 1.545 0.335 1.675 ;
 RECT 1.13 0.605 1.26 0.735 ;
 RECT 4.765 2.035 4.895 2.165 ;
 RECT 1.13 1.59 1.26 1.72 ;
 RECT 2.91 1.65 3.04 1.78 ;
 RECT 5.88 2.025 6.01 2.155 ;
 RECT 7.835 0.645 7.965 0.775 ;
 RECT 7.835 1.825 7.965 1.955 ;
 RECT 7.835 1.55 7.965 1.68 ;
 RECT 7.835 2.15 7.965 2.28 ;
 RECT 3.81 0.285 3.94 0.415 ;
 RECT 7.365 1.88 7.495 2.01 ;
 RECT 7.365 1.525 7.495 1.655 ;
 RECT 0.845 2.125 0.975 2.255 ;
 RECT 4.3 1.215 4.43 1.345 ;
 RECT 4.915 0.625 5.045 0.755 ;
 RECT 5.09 1.285 5.22 1.415 ;
 RECT 0.205 1.805 0.335 1.935 ;
 RECT 4.11 0.625 4.24 0.755 ;
 RECT 7.365 0.6 7.495 0.73 ;
 RECT 4.115 2 4.245 2.13 ;
 RECT 5.41 0.625 5.54 0.755 ;
 RECT 6.185 0.295 6.315 0.425 ;
 LAYER M1 ;
 RECT 4.76 0.76 4.9 2.235 ;
 RECT 4.76 0.62 5.1 0.76 ;
 RECT 3.195 0.575 3.335 0.605 ;
 RECT 3.195 0.745 3.335 2.265 ;
 RECT 3.185 0.605 3.965 0.745 ;
 RECT 3.825 0.745 3.965 1.205 ;
 RECT 4.29 1.165 4.61 1.205 ;
 RECT 4.47 0.395 4.61 1.165 ;
 RECT 4.29 1.35 4.48 1.4 ;
 RECT 4.29 1.345 4.61 1.35 ;
 RECT 3.825 1.205 4.61 1.345 ;
 RECT 5.875 0.395 6.015 2.21 ;
 RECT 4.47 0.255 6.015 0.395 ;
 RECT 1.71 0.515 1.85 2.025 ;
 RECT 1.71 2.165 1.85 2.295 ;
 RECT 2.52 1.775 2.66 2.025 ;
 RECT 2.52 2.165 2.66 2.415 ;
 RECT 2.905 1.585 3.045 1.635 ;
 RECT 2.905 1.775 3.045 1.835 ;
 RECT 1.71 2.025 2.66 2.165 ;
 RECT 3.475 1.12 3.615 2.415 ;
 RECT 3.475 0.89 3.65 1.12 ;
 RECT 2.52 1.635 3.055 1.775 ;
 RECT 2.52 2.415 3.62 2.555 ;
 RECT 5.405 2.49 6.73 2.615 ;
 RECT 5.415 2.615 6.73 2.63 ;
 RECT 5.405 1.87 5.545 2.49 ;
 RECT 5.36 0.62 5.68 0.76 ;
 RECT 5.54 0.76 5.68 1.73 ;
 RECT 5.405 1.73 5.68 1.87 ;
 RECT 6.59 1.3 6.73 2.49 ;
 RECT 6.59 1.16 7.22 1.295 ;
 RECT 6.99 1.145 7.22 1.16 ;
 RECT 6.59 1.295 7.18 1.3 ;
 RECT 6.175 0.245 6.425 0.475 ;
 RECT 6.285 0.475 6.425 2.09 ;
 RECT 6.18 2.09 6.425 2.32 ;
 RECT 6.185 0.22 6.425 0.245 ;
 RECT 0.65 0.51 0.79 1.06 ;
 RECT 0.65 1.2 0.79 1.775 ;
 RECT 0.65 1.06 1.56 1.2 ;
 RECT 1.42 0.365 1.56 1.06 ;
 RECT 1.42 0.225 2.13 0.365 ;
 RECT 1.99 0.365 2.13 0.965 ;
 RECT 3.8 0.235 3.95 0.265 ;
 RECT 3.8 0.405 3.95 0.465 ;
 RECT 2.62 0.265 3.95 0.405 ;
 RECT 1.99 0.965 2.76 1.105 ;
 RECT 2.62 0.405 2.76 0.965 ;
 END
END XOR3X2

MACRO ISOLANDAOX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.28 BY 2.88 ;
 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.315 0.91 2.71 1.24 ;
 END
 END ISO

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.8 1.185 5.22 1.565 ;
 END
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 5.36 1.16 6.71 1.3 ;
 RECT 6.57 1.44 6.71 1.565 ;
 RECT 6.265 1.3 6.71 1.44 ;
 RECT 6.57 0.885 6.71 1.075 ;
 RECT 6.265 1.075 6.71 1.16 ;
 RECT 4.275 0.365 4.415 0.825 ;
 RECT 4.275 0.825 5.5 0.965 ;
 RECT 5.36 0.965 5.5 1.16 ;
 END
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.28 2.96 ;
 RECT 4.345 2.27 4.575 2.8 ;
 RECT 4.98 2.57 5.12 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.28 0.08 ;
 RECT 2.44 0.305 2.705 0.445 ;
 RECT 4.96 0.08 5.45 0.42 ;
 RECT 3.805 0.08 3.945 0.57 ;
 RECT 2.505 0.445 2.645 0.48 ;
 RECT 2.505 0.08 2.645 0.305 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 1.445 1.99 7.745 2.13 ;
 RECT 2.44 1.395 2.72 1.535 ;
 RECT 7.56 0.935 7.79 1.425 ;
 RECT 1.365 1.1 1.595 1.59 ;
 RECT 7.1 0.43 7.24 1.99 ;
 RECT 2.505 1.535 2.645 1.99 ;
 RECT 7.605 1.425 7.745 1.99 ;
 RECT 1.45 1.59 1.59 1.99 ;
 END
 END VDDG

 OBS
 LAYER PO ;
 RECT 2.76 0.09 2.86 0.575 ;
 RECT 2.76 0.805 2.86 1.85 ;
 RECT 2.63 0.575 2.86 0.805 ;
 RECT 2.29 0.09 2.39 0.985 ;
 RECT 2.29 1.215 2.39 1.87 ;
 RECT 2.285 0.985 2.515 1.215 ;
 RECT 4.685 1.37 5.02 1.375 ;
 RECT 4.775 1.375 5.02 1.44 ;
 RECT 4.685 1.21 5.02 1.27 ;
 RECT 3.47 1.115 3.57 1.27 ;
 RECT 3.06 0.09 3.16 1.015 ;
 RECT 4.775 1.44 4.875 2.405 ;
 RECT 3.06 1.015 3.57 1.115 ;
 RECT 3.47 1.27 5.02 1.37 ;
 RECT 6.29 0.365 6.39 0.86 ;
 RECT 6.85 0.365 6.95 1.9 ;
 RECT 3.905 0.86 6.39 0.96 ;
 RECT 3.905 0.96 4.16 1.09 ;
 RECT 4.06 0.1 4.16 0.86 ;
 RECT 6.29 0.265 6.95 0.365 ;
 LAYER CO ;
 RECT 4.985 2.625 5.115 2.755 ;
 RECT 4.525 1.65 4.655 1.78 ;
 RECT 5.27 0.255 5.4 0.385 ;
 RECT 5.01 0.255 5.14 0.385 ;
 RECT 7.61 1.235 7.74 1.365 ;
 RECT 7.61 0.975 7.74 1.105 ;
 RECT 3.955 0.91 4.085 1.04 ;
 RECT 4.84 1.26 4.97 1.39 ;
 RECT 2.68 0.625 2.81 0.755 ;
 RECT 4.28 0.42 4.41 0.55 ;
 RECT 7.105 0.66 7.235 0.79 ;
 RECT 7.105 0.99 7.235 1.12 ;
 RECT 3.81 0.39 3.94 0.52 ;
 RECT 6.575 1.365 6.705 1.495 ;
 RECT 2.335 1.035 2.465 1.165 ;
 RECT 3.28 0.31 3.41 0.44 ;
 RECT 6.575 1.025 6.705 1.155 ;
 RECT 2.51 0.31 2.64 0.44 ;
 RECT 2.51 1.4 2.64 1.53 ;
 RECT 2.04 0.31 2.17 0.44 ;
 RECT 2.04 1.335 2.17 1.465 ;
 RECT 4.395 2.455 4.525 2.585 ;
 RECT 2.98 1.335 3.11 1.465 ;
 RECT 1.415 1.4 1.545 1.53 ;
 RECT 1.415 1.14 1.545 1.27 ;
 LAYER M1 ;
 RECT 2.035 0.24 2.175 0.62 ;
 RECT 2.035 0.76 2.175 1.725 ;
 RECT 2.035 0.62 2.88 0.76 ;
 RECT 3.275 0.89 3.415 1.185 ;
 RECT 2.975 1.115 3.115 1.185 ;
 RECT 2.975 1.325 3.115 1.535 ;
 RECT 3.275 0.24 3.415 0.75 ;
 RECT 3.885 0.89 4.135 1.185 ;
 RECT 3.885 1.325 4.135 1.33 ;
 RECT 3.275 0.75 4.135 0.89 ;
 RECT 4.52 1.325 4.66 1.85 ;
 RECT 2.975 1.185 4.66 1.325 ;
 END
END ISOLANDAOX1

MACRO ISOLANDAOX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.6 BY 2.88 ;
 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.315 0.915 2.71 1.24 ;
 END
 END ISO

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.8 1.185 5.22 1.565 ;
 END
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.57 0.31 7.71 0.45 ;
 RECT 5.36 1.16 6.71 1.3 ;
 RECT 6.265 1.075 6.71 1.16 ;
 RECT 7.57 0.45 7.71 1.565 ;
 RECT 6.57 0.45 6.71 1.075 ;
 RECT 4.275 0.365 4.415 0.825 ;
 RECT 6.57 1.44 6.71 1.565 ;
 RECT 6.265 1.3 6.71 1.44 ;
 RECT 4.275 0.825 5.5 0.965 ;
 RECT 5.36 0.965 5.5 1.16 ;
 END
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.6 2.96 ;
 RECT 4.345 2.27 4.575 2.8 ;
 RECT 4.98 2.57 5.12 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.6 0.08 ;
 RECT 2.44 0.305 2.705 0.445 ;
 RECT 5.15 0.08 5.64 0.42 ;
 RECT 3.805 0.08 3.945 0.57 ;
 RECT 4.75 0.08 4.89 0.57 ;
 RECT 2.505 0.445 2.645 0.48 ;
 RECT 2.505 0.08 2.645 0.305 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 2.44 1.395 2.72 1.535 ;
 RECT 8.065 0.925 8.295 1.415 ;
 RECT 1.365 1.1 1.595 1.59 ;
 RECT 7.1 0.59 7.24 1.99 ;
 RECT 1.45 1.99 8.25 2.13 ;
 RECT 2.505 1.535 2.645 1.99 ;
 RECT 8.11 1.415 8.25 1.99 ;
 RECT 1.45 1.59 1.59 1.99 ;
 END
 END VDDG

 OBS
 LAYER PO ;
 RECT 2.76 0.09 2.86 0.575 ;
 RECT 2.76 0.805 2.86 1.85 ;
 RECT 2.63 0.575 2.86 0.805 ;
 RECT 2.29 0.09 2.39 0.985 ;
 RECT 2.29 1.215 2.39 1.87 ;
 RECT 2.285 0.985 2.515 1.215 ;
 RECT 4.685 1.37 5.02 1.375 ;
 RECT 4.775 1.375 5.02 1.44 ;
 RECT 4.685 1.21 5.02 1.27 ;
 RECT 3.47 1.115 3.57 1.27 ;
 RECT 3.06 0.09 3.16 1.015 ;
 RECT 4.775 1.44 4.875 2.405 ;
 RECT 3.06 1.015 3.57 1.115 ;
 RECT 3.47 1.27 5.02 1.37 ;
 RECT 3.905 0.96 4.16 1.09 ;
 RECT 6.29 0.365 6.39 0.86 ;
 RECT 3.905 0.86 6.39 0.96 ;
 RECT 7.355 0.365 7.455 1.9 ;
 RECT 6.85 0.365 6.95 1.9 ;
 RECT 4.06 0.11 4.16 0.86 ;
 RECT 4.53 0.11 4.63 0.86 ;
 RECT 4.53 0.96 4.63 0.97 ;
 RECT 6.29 0.265 7.455 0.365 ;
 LAYER CO ;
 RECT 4.985 2.625 5.115 2.755 ;
 RECT 4.525 1.65 4.655 1.78 ;
 RECT 5.46 0.255 5.59 0.385 ;
 RECT 5.2 0.255 5.33 0.385 ;
 RECT 8.115 1.225 8.245 1.355 ;
 RECT 8.115 0.965 8.245 1.095 ;
 RECT 3.955 0.91 4.085 1.04 ;
 RECT 4.84 1.26 4.97 1.39 ;
 RECT 2.68 0.625 2.81 0.755 ;
 RECT 4.28 0.42 4.41 0.55 ;
 RECT 7.105 0.66 7.235 0.79 ;
 RECT 7.105 0.99 7.235 1.12 ;
 RECT 3.81 0.39 3.94 0.52 ;
 RECT 6.575 1.365 6.705 1.495 ;
 RECT 2.335 1.035 2.465 1.165 ;
 RECT 3.28 0.31 3.41 0.44 ;
 RECT 6.575 1.025 6.705 1.155 ;
 RECT 2.51 0.31 2.64 0.44 ;
 RECT 2.51 1.4 2.64 1.53 ;
 RECT 2.04 0.31 2.17 0.44 ;
 RECT 2.04 1.335 2.17 1.465 ;
 RECT 4.395 2.455 4.525 2.585 ;
 RECT 7.105 1.32 7.235 1.45 ;
 RECT 7.575 1.365 7.705 1.495 ;
 RECT 7.575 1.025 7.705 1.155 ;
 RECT 4.755 0.39 4.885 0.52 ;
 RECT 2.98 1.335 3.11 1.465 ;
 RECT 1.415 1.4 1.545 1.53 ;
 RECT 1.415 1.14 1.545 1.27 ;
 LAYER M1 ;
 RECT 2.035 0.24 2.175 0.62 ;
 RECT 2.035 0.76 2.175 1.535 ;
 RECT 2.035 0.62 2.88 0.76 ;
 RECT 2.975 1.325 3.115 1.605 ;
 RECT 3.275 0.24 3.415 0.75 ;
 RECT 3.885 0.89 4.135 1.185 ;
 RECT 3.885 1.325 4.135 1.33 ;
 RECT 3.275 0.75 4.135 0.89 ;
 RECT 4.52 1.325 4.66 1.85 ;
 RECT 2.975 1.185 4.66 1.325 ;
 END
END ISOLANDAOX2

MACRO ISOLANDAOX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.24 BY 2.88 ;
 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 2.44 1.465 2.72 1.605 ;
 RECT 2.505 1.45 2.645 1.465 ;
 RECT 1.45 1.99 9.025 2.13 ;
 RECT 1.365 1.1 1.595 1.59 ;
 RECT 8.78 0.935 9.01 1.425 ;
 RECT 2.505 1.605 2.645 1.99 ;
 RECT 6.9 0.59 7.04 1.99 ;
 RECT 7.84 0.595 7.98 1.99 ;
 RECT 1.45 1.59 1.59 1.99 ;
 RECT 8.825 1.425 8.965 1.99 ;
 END
 END VDDG

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.16 1.205 6.57 1.57 ;
 RECT 4.275 0.365 4.415 0.825 ;
 RECT 7.37 0.405 7.51 1.56 ;
 RECT 8.31 0.405 8.45 1.545 ;
 RECT 6.43 0.265 8.45 0.405 ;
 RECT 8.31 0.26 8.45 0.265 ;
 RECT 5.22 0.35 5.36 0.825 ;
 RECT 4.275 0.825 6.57 0.965 ;
 RECT 6.43 0.965 6.57 1.205 ;
 RECT 6.43 0.405 6.57 0.825 ;
 END
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.24 0.08 ;
 RECT 2.44 0.305 2.705 0.445 ;
 RECT 0.985 0.08 1.475 0.42 ;
 RECT 3.805 0.08 3.945 0.57 ;
 RECT 4.745 0.08 4.885 0.62 ;
 RECT 5.72 0.08 5.86 0.62 ;
 RECT 2.505 0.445 2.645 0.48 ;
 RECT 2.505 0.08 2.645 0.305 ;
 END
 END VSS

 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.315 1.025 2.71 1.285 ;
 END
 END ISO

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.24 2.96 ;
 RECT 4.345 2.27 4.575 2.8 ;
 RECT 4.98 2.57 5.12 2.8 ;
 END
 END VDD

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.8 1.185 5.22 1.565 ;
 END
 END D

 OBS
 LAYER PO ;
 RECT 2.76 0.09 2.86 0.645 ;
 RECT 2.76 0.875 2.86 1.85 ;
 RECT 2.63 0.645 2.86 0.875 ;
 RECT 2.29 0.09 2.39 1.03 ;
 RECT 2.29 1.26 2.39 1.87 ;
 RECT 2.285 1.03 2.515 1.26 ;
 RECT 4.685 1.37 5.02 1.375 ;
 RECT 4.775 1.375 5.02 1.44 ;
 RECT 4.775 1.44 4.875 2.405 ;
 RECT 4.685 1.21 5.02 1.27 ;
 RECT 3.47 1.115 3.57 1.27 ;
 RECT 3.06 0.09 3.16 1.015 ;
 RECT 3.06 1.015 3.57 1.115 ;
 RECT 3.47 1.27 5.02 1.37 ;
 RECT 5.975 0.365 6.075 0.87 ;
 RECT 8.095 0.365 8.195 1.9 ;
 RECT 7.625 0.365 7.725 1.9 ;
 RECT 7.155 0.365 7.255 1.9 ;
 RECT 6.685 0.365 6.785 1.9 ;
 RECT 3.905 0.86 4.16 0.87 ;
 RECT 3.905 0.87 6.075 0.97 ;
 RECT 3.905 0.97 4.16 1.09 ;
 RECT 5.505 0.1 5.605 0.87 ;
 RECT 5.005 0.1 5.105 0.87 ;
 RECT 4.53 0.1 4.63 0.87 ;
 RECT 4.06 0.1 4.16 0.86 ;
 RECT 5.975 0.265 8.2 0.365 ;
 LAYER CO ;
 RECT 6.435 1.025 6.565 1.155 ;
 RECT 1.415 1.14 1.545 1.27 ;
 RECT 1.415 1.4 1.545 1.53 ;
 RECT 8.315 0.66 8.445 0.79 ;
 RECT 8.315 0.99 8.445 1.12 ;
 RECT 7.845 0.66 7.975 0.79 ;
 RECT 7.845 0.99 7.975 1.12 ;
 RECT 7.375 0.66 7.505 0.79 ;
 RECT 7.375 0.99 7.505 1.12 ;
 RECT 5.725 0.42 5.855 0.55 ;
 RECT 5.225 0.42 5.355 0.55 ;
 RECT 4.75 0.42 4.88 0.55 ;
 RECT 8.83 0.975 8.96 1.105 ;
 RECT 6.905 0.66 7.035 0.79 ;
 RECT 6.905 0.99 7.035 1.12 ;
 RECT 2.335 1.08 2.465 1.21 ;
 RECT 3.81 0.39 3.94 0.52 ;
 RECT 4.84 1.26 4.97 1.39 ;
 RECT 3.955 0.91 4.085 1.04 ;
 RECT 2.98 1.405 3.11 1.535 ;
 RECT 8.83 1.235 8.96 1.365 ;
 RECT 4.28 0.42 4.41 0.55 ;
 RECT 2.51 0.31 2.64 0.44 ;
 RECT 3.28 0.31 3.41 0.44 ;
 RECT 4.395 2.455 4.525 2.585 ;
 RECT 2.68 0.695 2.81 0.825 ;
 RECT 6.435 1.365 6.565 1.495 ;
 RECT 2.04 1.405 2.17 1.535 ;
 RECT 1.035 0.255 1.165 0.385 ;
 RECT 1.295 0.255 1.425 0.385 ;
 RECT 2.04 0.31 2.17 0.44 ;
 RECT 4.525 1.65 4.655 1.78 ;
 RECT 2.51 1.47 2.64 1.6 ;
 RECT 4.985 2.625 5.115 2.755 ;
 LAYER M1 ;
 RECT 2.035 0.24 2.175 0.69 ;
 RECT 2.035 0.83 2.175 1.725 ;
 RECT 2.675 0.625 2.815 0.69 ;
 RECT 2.675 0.83 2.815 0.885 ;
 RECT 2.035 0.69 2.815 0.83 ;
 RECT 3.275 0.24 3.415 0.75 ;
 RECT 2.975 0.89 3.115 1.605 ;
 RECT 3.885 0.89 4.135 1.185 ;
 RECT 3.885 1.325 4.135 1.33 ;
 RECT 2.975 0.75 4.135 0.89 ;
 RECT 3.885 1.185 4.66 1.325 ;
 RECT 4.52 1.325 4.66 1.85 ;
 END
END ISOLANDAOX4

MACRO ISOLANDAOX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 15.36 BY 2.88 ;
 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.96 0.9 2.355 1.24 ;
 END
 END ISO

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.8 1.185 5.22 1.565 ;
 END
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 9.275 1.44 9.415 1.565 ;
 RECT 9.275 0.31 13.27 0.45 ;
 RECT 5.36 1.16 9.415 1.3 ;
 RECT 8.97 1.3 9.415 1.44 ;
 RECT 8.97 1.075 9.415 1.16 ;
 RECT 9.275 0.45 9.415 1.075 ;
 RECT 10.275 0.45 10.415 1.565 ;
 RECT 11.215 0.45 11.355 1.565 ;
 RECT 12.19 0.45 12.33 1.565 ;
 RECT 13.13 0.45 13.27 1.565 ;
 RECT 5.22 0.35 5.36 0.825 ;
 RECT 4.275 0.825 7.32 0.965 ;
 RECT 4.275 0.35 4.415 0.825 ;
 RECT 6.16 0.35 6.3 0.825 ;
 RECT 7.105 0.35 7.245 0.825 ;
 RECT 5.36 0.965 5.5 1.16 ;
 END
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 15.36 2.96 ;
 RECT 4.45 2.27 4.68 2.8 ;
 RECT 4.98 2.57 5.12 2.8 ;
 END
 END VDD

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 15.36 0.08 ;
 RECT 0.875 0.305 1.145 0.445 ;
 RECT 8.04 0.08 8.27 0.71 ;
 RECT 1.9 0.08 2.17 0.255 ;
 RECT 3.805 0.08 3.945 0.59 ;
 RECT 4.75 0.08 4.89 0.59 ;
 RECT 5.69 0.08 5.83 0.59 ;
 RECT 6.635 0.08 6.775 0.59 ;
 RECT 7.575 0.08 7.715 0.59 ;
 RECT 0.94 0.08 1.08 0.305 ;
 END
 END VSS

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 2.08 1.395 2.36 1.535 ;
 RECT 13.625 0.925 13.855 1.415 ;
 RECT 1.22 1.345 1.45 1.705 ;
 RECT 2.145 1.535 2.285 1.99 ;
 RECT 9.805 0.59 9.945 1.99 ;
 RECT 10.745 0.59 10.885 1.99 ;
 RECT 3.095 1.33 3.235 1.99 ;
 RECT 11.72 0.59 11.86 1.99 ;
 RECT 12.66 0.59 12.8 1.99 ;
 RECT 13.67 1.415 13.81 1.99 ;
 RECT 1.265 1.705 1.405 1.99 ;
 RECT 1.265 1.99 13.81 2.13 ;
 END
 END VDDG

 OBS
 LAYER PO ;
 RECT 0.725 0.09 0.825 1.015 ;
 RECT 1.93 0.985 2.16 1.015 ;
 RECT 1.93 1.115 2.16 1.215 ;
 RECT 0.725 1.015 2.16 1.115 ;
 RECT 1.93 1.215 2.03 1.87 ;
 RECT 8.995 0.365 9.095 0.86 ;
 RECT 8.995 0.265 13.015 0.365 ;
 RECT 12.915 0.365 13.015 1.9 ;
 RECT 11.975 0.365 12.075 1.9 ;
 RECT 11.47 0.365 11.57 1.9 ;
 RECT 12.445 0.365 12.545 1.9 ;
 RECT 11 0.365 11.1 1.9 ;
 RECT 10.53 0.365 10.63 1.9 ;
 RECT 10.06 0.365 10.16 1.9 ;
 RECT 9.555 0.365 9.655 1.9 ;
 RECT 3.905 0.86 9.105 0.96 ;
 RECT 3.905 0.96 4.16 1.09 ;
 RECT 7.36 0.11 7.46 0.86 ;
 RECT 7.36 0.96 7.46 0.97 ;
 RECT 6.415 0.11 6.515 0.86 ;
 RECT 6.415 0.96 6.515 0.97 ;
 RECT 6.89 0.11 6.99 0.86 ;
 RECT 6.89 0.96 6.99 0.97 ;
 RECT 5.945 0.11 6.045 0.86 ;
 RECT 5.945 0.96 6.045 0.975 ;
 RECT 5.475 0.11 5.575 0.86 ;
 RECT 5.475 0.96 5.575 0.97 ;
 RECT 5.005 0.11 5.105 0.86 ;
 RECT 5.005 0.96 5.105 0.97 ;
 RECT 4.53 0.11 4.63 0.86 ;
 RECT 4.53 0.96 4.63 0.97 ;
 RECT 4.06 0.11 4.16 0.86 ;
 RECT 4.775 1.375 5.02 1.44 ;
 RECT 4.775 1.44 4.875 2.405 ;
 RECT 3.47 0.925 3.57 1.27 ;
 RECT 3.17 0.09 3.27 0.825 ;
 RECT 2.69 0.09 2.79 0.825 ;
 RECT 4.685 1.21 5.02 1.27 ;
 RECT 4.685 1.37 5.02 1.375 ;
 RECT 5.28 1.37 5.38 2.405 ;
 RECT 2.69 0.825 3.57 0.925 ;
 RECT 3.47 1.27 5.385 1.37 ;
 RECT 2.4 0.76 2.5 1.75 ;
 RECT 2.88 1.105 2.98 1.75 ;
 RECT 2.22 0.09 2.32 0.66 ;
 RECT 1.75 0.09 1.85 0.66 ;
 RECT 1.005 0.575 1.235 0.66 ;
 RECT 1.005 0.76 1.235 0.805 ;
 RECT 1.005 0.66 2.5 0.76 ;
 RECT 2.4 1.75 2.98 1.85 ;
 LAYER CO ;
 RECT 4.28 0.42 4.41 0.55 ;
 RECT 9.81 0.66 9.94 0.79 ;
 RECT 9.81 0.99 9.94 1.12 ;
 RECT 3.81 0.39 3.94 0.52 ;
 RECT 9.28 1.365 9.41 1.495 ;
 RECT 1.98 1.035 2.11 1.165 ;
 RECT 2.92 0.505 3.05 0.635 ;
 RECT 9.28 1.025 9.41 1.155 ;
 RECT 0.945 0.31 1.075 0.44 ;
 RECT 2.15 1.4 2.28 1.53 ;
 RECT 0.475 0.31 0.605 0.44 ;
 RECT 1.68 1.335 1.81 1.465 ;
 RECT 7.11 0.42 7.24 0.55 ;
 RECT 6.64 0.39 6.77 0.52 ;
 RECT 6.165 0.42 6.295 0.55 ;
 RECT 12.665 1.32 12.795 1.45 ;
 RECT 11.725 1.32 11.855 1.45 ;
 RECT 12.665 0.66 12.795 0.79 ;
 RECT 12.195 1.365 12.325 1.495 ;
 RECT 12.665 0.99 12.795 1.12 ;
 RECT 13.135 1.365 13.265 1.495 ;
 RECT 12.195 1.025 12.325 1.155 ;
 RECT 13.135 1.025 13.265 1.155 ;
 RECT 11.725 0.66 11.855 0.79 ;
 RECT 11.725 0.99 11.855 1.12 ;
 RECT 5.5 1.65 5.63 1.78 ;
 RECT 1.495 0.31 1.625 0.44 ;
 RECT 4.5 2.455 4.63 2.585 ;
 RECT 3.39 0.31 3.52 0.44 ;
 RECT 2.44 0.31 2.57 0.44 ;
 RECT 1.97 0.11 2.1 0.24 ;
 RECT 3.1 1.4 3.23 1.53 ;
 RECT 11.22 1.365 11.35 1.495 ;
 RECT 11.22 1.025 11.35 1.155 ;
 RECT 10.75 1.32 10.88 1.45 ;
 RECT 10.75 0.66 10.88 0.79 ;
 RECT 10.75 0.99 10.88 1.12 ;
 RECT 5.695 0.39 5.825 0.52 ;
 RECT 5.225 0.42 5.355 0.55 ;
 RECT 9.81 1.32 9.94 1.45 ;
 RECT 10.28 1.365 10.41 1.495 ;
 RECT 10.28 1.025 10.41 1.155 ;
 RECT 4.755 0.39 4.885 0.52 ;
 RECT 2.62 1.335 2.75 1.465 ;
 RECT 1.27 1.515 1.4 1.645 ;
 RECT 7.58 0.39 7.71 0.52 ;
 RECT 4.985 2.625 5.115 2.755 ;
 RECT 4.525 1.65 4.655 1.78 ;
 RECT 8.09 0.53 8.22 0.66 ;
 RECT 8.09 0.27 8.22 0.4 ;
 RECT 13.675 1.225 13.805 1.355 ;
 RECT 13.675 0.965 13.805 1.095 ;
 RECT 3.955 0.91 4.085 1.04 ;
 RECT 4.84 1.26 4.97 1.39 ;
 RECT 1.055 0.625 1.185 0.755 ;
 LAYER M1 ;
 RECT 0.47 0.24 0.61 0.62 ;
 RECT 0.47 0.76 0.61 0.95 ;
 RECT 0.47 0.62 1.255 0.76 ;
 RECT 0.47 0.95 1.815 1.085 ;
 RECT 0.48 1.085 1.815 1.09 ;
 RECT 1.675 1.09 1.815 1.535 ;
 RECT 1.49 0.24 1.63 0.395 ;
 RECT 2.435 0.36 2.575 0.395 ;
 RECT 3.385 0.36 3.525 0.5 ;
 RECT 1.425 0.395 2.575 0.535 ;
 RECT 2.435 0.22 3.525 0.36 ;
 RECT 2.915 0.64 3.055 1.05 ;
 RECT 2.615 1.19 2.755 1.605 ;
 RECT 5.495 1.58 5.635 1.71 ;
 RECT 2.615 1.185 4.66 1.19 ;
 RECT 3.885 1.19 4.66 1.325 ;
 RECT 4.52 1.325 4.66 1.71 ;
 RECT 3.885 0.75 4.135 1.05 ;
 RECT 2.615 1.05 4.135 1.185 ;
 RECT 3.885 1.325 4.135 1.33 ;
 RECT 2.85 0.5 3.12 0.64 ;
 RECT 4.45 1.71 5.7 1.85 ;
 END
END ISOLANDAOX8

MACRO ISOLORAOX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.6 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.215 1.48 1.555 1.72 ;
 RECT 1.155 1.17 1.385 1.31 ;
 RECT 1.215 1.31 1.355 1.48 ;
 END
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.6 2.96 ;
 RECT 0.41 1.945 0.55 2.8 ;
 RECT 2.3 1.91 2.44 2.8 ;
 RECT 1.32 1.91 1.46 2.8 ;
 END
 END VDD

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 4.15 2.48 8.105 2.62 ;
 RECT 4.15 1.35 4.29 2.48 ;
 RECT 7.965 1.105 8.105 2.48 ;
 RECT 6.315 1.345 6.455 2.48 ;
 RECT 7.265 1.345 7.405 2.48 ;
 END
 END VDDG

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.56 0.79 6.935 1.07 ;
 RECT 6.795 1.07 6.935 1.845 ;
 RECT 6.795 0.22 6.935 0.79 ;
 END
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.6 0.08 ;
 RECT 5.1 0.08 5.24 0.545 ;
 RECT 3.6 0.34 3.875 0.48 ;
 RECT 1.32 0.08 1.46 0.715 ;
 RECT 0.41 0.08 0.55 0.765 ;
 RECT 6.31 0.08 6.45 0.535 ;
 RECT 7.28 0.08 7.42 0.535 ;
 RECT 3.67 0.08 3.81 0.34 ;
 RECT 2.3 0.08 2.44 0.73 ;
 END
 END VSS

 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.635 0.62 4 0.875 ;
 END
 END ISO

 OBS
 LAYER PO ;
 RECT 1.575 1.12 1.895 1.125 ;
 RECT 1.575 0.315 1.675 1.12 ;
 RECT 1.575 1.225 1.895 1.35 ;
 RECT 1.575 1.35 1.675 2.74 ;
 RECT 2.085 0.315 2.185 1.125 ;
 RECT 2.085 1.225 2.185 2.74 ;
 RECT 1.575 1.125 2.185 1.225 ;
 RECT 1.105 0.44 1.205 1.125 ;
 RECT 1.105 1.125 1.385 1.355 ;
 RECT 1.105 1.355 1.205 2.24 ;
 RECT 3.925 0.83 4.025 1.025 ;
 RECT 3.925 1.125 4.025 1.95 ;
 RECT 4.405 1.125 4.505 1.95 ;
 RECT 3.925 0.09 4.025 0.62 ;
 RECT 3.77 0.62 4.025 0.83 ;
 RECT 3.925 1.025 4.505 1.125 ;
 RECT 7.05 0.095 7.15 0.845 ;
 RECT 7.05 0.945 7.15 1.95 ;
 RECT 6.57 0.095 6.67 0.845 ;
 RECT 6.57 0.945 6.67 1.95 ;
 RECT 6.06 0.765 6.29 0.845 ;
 RECT 6.06 0.945 6.29 0.975 ;
 RECT 6.06 0.845 7.15 0.945 ;
 RECT 5.085 1.95 5.185 2.305 ;
 RECT 3.3 1.145 3.4 2.305 ;
 RECT 5.365 1.015 5.465 1.85 ;
 RECT 4.88 1.85 5.465 1.95 ;
 RECT 4.88 0.125 4.98 1.85 ;
 RECT 2.475 1.095 3.4 1.145 ;
 RECT 2.475 1.145 2.705 1.305 ;
 RECT 2.565 1.045 3.4 1.095 ;
 RECT 3.3 2.305 5.185 2.405 ;
 LAYER CO ;
 RECT 6.8 0.335 6.93 0.465 ;
 RECT 7.285 0.335 7.415 0.465 ;
 RECT 6.315 0.335 6.445 0.465 ;
 RECT 7.27 1.45 7.4 1.58 ;
 RECT 6.8 1.45 6.93 1.58 ;
 RECT 6.32 1.45 6.45 1.58 ;
 RECT 1.325 1.96 1.455 2.09 ;
 RECT 1.815 1.645 1.945 1.775 ;
 RECT 2.305 1.96 2.435 2.09 ;
 RECT 0.855 1.69 0.985 1.82 ;
 RECT 1.205 1.175 1.335 1.305 ;
 RECT 2.305 0.55 2.435 0.68 ;
 RECT 1.815 0.62 1.945 0.75 ;
 RECT 1.815 1.95 1.945 2.08 ;
 RECT 1.325 0.535 1.455 0.665 ;
 RECT 7.97 1.175 8.1 1.305 ;
 RECT 7.97 1.435 8.1 1.565 ;
 RECT 0.415 0.305 0.545 0.435 ;
 RECT 0.415 0.565 0.545 0.695 ;
 RECT 0.415 2.015 0.545 2.145 ;
 RECT 0.415 2.275 0.545 2.405 ;
 RECT 3.675 0.345 3.805 0.475 ;
 RECT 3.665 1.45 3.795 1.58 ;
 RECT 5.105 0.345 5.235 0.475 ;
 RECT 4.145 0.345 4.275 0.475 ;
 RECT 5.62 1.45 5.75 1.58 ;
 RECT 5.1 1.45 5.23 1.58 ;
 RECT 4.155 1.45 4.285 1.58 ;
 RECT 4.63 1.45 4.76 1.58 ;
 RECT 0.855 0.755 0.985 0.885 ;
 RECT 1.815 1.645 1.945 1.775 ;
 RECT 1.715 1.17 1.845 1.3 ;
 RECT 3.82 0.66 3.95 0.79 ;
 RECT 6.11 0.805 6.24 0.935 ;
 RECT 2.525 1.135 2.655 1.265 ;
 LAYER M1 ;
 RECT 0.85 0.995 0.99 1.87 ;
 RECT 0.85 0.7 0.99 0.855 ;
 RECT 1.71 1.26 1.85 1.35 ;
 RECT 1.53 1.12 1.85 1.26 ;
 RECT 0.85 0.855 1.67 0.995 ;
 RECT 1.53 0.995 1.67 1.12 ;
 RECT 3.66 1.155 3.8 1.7 ;
 RECT 5.615 1.155 5.755 1.71 ;
 RECT 4.625 1.155 4.765 1.675 ;
 RECT 3.66 1.015 5.755 1.155 ;
 RECT 4.14 0.265 4.28 0.735 ;
 RECT 5.095 1.35 5.235 1.945 ;
 RECT 6.035 0.975 6.175 1.945 ;
 RECT 4.14 0.765 6.29 0.875 ;
 RECT 4.14 0.735 6.175 0.765 ;
 RECT 6.035 0.875 6.29 0.975 ;
 RECT 5.095 1.945 6.175 2.085 ;
 RECT 1.81 1.685 1.95 2.36 ;
 RECT 1.81 0.57 1.95 0.835 ;
 RECT 2.02 0.975 2.16 1.13 ;
 RECT 2.02 1.27 2.16 1.545 ;
 RECT 1.81 0.835 2.16 0.975 ;
 RECT 1.81 1.545 2.16 1.685 ;
 RECT 2.475 1.095 2.705 1.13 ;
 RECT 2.475 1.27 2.705 1.305 ;
 RECT 1.99 1.13 2.705 1.27 ;
 END
END ISOLORAOX1

MACRO ISOLORAOX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 10.24 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 10.24 0.08 ;
 RECT 5.1 0.08 5.24 0.545 ;
 RECT 3.6 0.34 3.875 0.48 ;
 RECT 1.32 0.08 1.46 0.715 ;
 RECT 6.31 0.08 6.45 0.535 ;
 RECT 7.28 0.08 7.42 0.535 ;
 RECT 0.41 0.08 0.55 0.765 ;
 RECT 8.255 0.08 8.395 0.535 ;
 RECT 2.3 0.08 2.44 0.73 ;
 RECT 3.67 0.08 3.81 0.34 ;
 END
 END VSS

 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.635 0.62 4 0.875 ;
 END
 END ISO

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.795 1.07 6.935 1.845 ;
 RECT 6.795 0.22 6.935 0.79 ;
 RECT 6.56 0.87 7.91 1.01 ;
 RECT 6.56 1.01 6.935 1.07 ;
 RECT 6.56 0.79 6.935 0.87 ;
 RECT 7.77 1.01 7.91 1.845 ;
 RECT 7.77 0.22 7.91 0.87 ;
 END
 END Q

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 4.15 1.35 4.29 2.48 ;
 RECT 8.805 1.105 8.945 2.48 ;
 RECT 4.15 2.48 8.945 2.62 ;
 RECT 7.265 1.345 7.405 2.48 ;
 RECT 6.315 1.345 6.455 2.48 ;
 RECT 8.24 1.345 8.38 2.48 ;
 END
 END VDDG

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.215 1.48 1.555 1.72 ;
 RECT 1.155 1.17 1.385 1.31 ;
 RECT 1.215 1.31 1.355 1.48 ;
 END
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 10.24 2.96 ;
 RECT 0.41 1.945 0.55 2.8 ;
 RECT 2.3 1.91 2.44 2.8 ;
 RECT 1.32 1.91 1.46 2.8 ;
 END
 END VDD

 OBS
 LAYER PO ;
 RECT 1.105 0.44 1.205 1.125 ;
 RECT 1.105 1.125 1.385 1.355 ;
 RECT 1.105 1.355 1.205 2.24 ;
 RECT 1.575 1.12 1.895 1.125 ;
 RECT 1.575 0.315 1.675 1.12 ;
 RECT 1.575 1.225 1.895 1.35 ;
 RECT 1.575 1.35 1.675 2.74 ;
 RECT 2.085 0.315 2.185 1.125 ;
 RECT 2.085 1.225 2.185 2.74 ;
 RECT 1.575 1.125 2.185 1.225 ;
 RECT 5.085 1.95 5.185 2.305 ;
 RECT 3.3 1.145 3.4 2.305 ;
 RECT 5.365 1.015 5.465 1.85 ;
 RECT 4.88 1.85 5.465 1.95 ;
 RECT 4.88 0.125 4.98 1.85 ;
 RECT 2.475 1.095 3.4 1.145 ;
 RECT 2.475 1.145 2.705 1.305 ;
 RECT 2.565 1.045 3.4 1.095 ;
 RECT 3.3 2.305 5.185 2.405 ;
 RECT 3.925 0.83 4.025 1.025 ;
 RECT 3.925 1.125 4.025 1.95 ;
 RECT 4.405 1.125 4.505 1.95 ;
 RECT 3.925 0.09 4.025 0.62 ;
 RECT 3.77 0.62 4.025 0.83 ;
 RECT 3.925 1.025 4.505 1.125 ;
 RECT 8.025 0.095 8.125 0.845 ;
 RECT 8.025 0.945 8.125 1.95 ;
 RECT 6.06 0.845 8.125 0.945 ;
 RECT 7.05 0.095 7.15 0.845 ;
 RECT 7.05 0.945 7.15 1.95 ;
 RECT 6.57 0.095 6.67 0.845 ;
 RECT 6.57 0.945 6.67 1.95 ;
 RECT 7.545 0.095 7.645 0.845 ;
 RECT 7.545 0.945 7.645 1.95 ;
 RECT 6.06 0.765 6.29 0.845 ;
 RECT 6.06 0.945 6.29 0.975 ;
 LAYER CO ;
 RECT 1.325 1.96 1.455 2.09 ;
 RECT 2.305 1.96 2.435 2.09 ;
 RECT 7.27 1.45 7.4 1.58 ;
 RECT 6.8 0.335 6.93 0.465 ;
 RECT 6.32 1.45 6.45 1.58 ;
 RECT 0.415 2.015 0.545 2.145 ;
 RECT 3.665 1.45 3.795 1.58 ;
 RECT 0.415 0.305 0.545 0.435 ;
 RECT 1.815 1.645 1.945 1.775 ;
 RECT 4.145 0.345 4.275 0.475 ;
 RECT 5.105 0.345 5.235 0.475 ;
 RECT 0.415 0.565 0.545 0.695 ;
 RECT 8.81 1.435 8.94 1.565 ;
 RECT 6.8 1.45 6.93 1.58 ;
 RECT 0.855 1.69 0.985 1.82 ;
 RECT 6.315 0.335 6.445 0.465 ;
 RECT 0.415 2.275 0.545 2.405 ;
 RECT 1.815 1.645 1.945 1.775 ;
 RECT 4.155 1.45 4.285 1.58 ;
 RECT 8.81 1.175 8.94 1.305 ;
 RECT 1.325 0.535 1.455 0.665 ;
 RECT 1.715 1.17 1.845 1.3 ;
 RECT 1.205 1.175 1.335 1.305 ;
 RECT 2.305 0.55 2.435 0.68 ;
 RECT 3.675 0.345 3.805 0.475 ;
 RECT 1.815 1.95 1.945 2.08 ;
 RECT 1.815 0.62 1.945 0.75 ;
 RECT 5.1 1.45 5.23 1.58 ;
 RECT 4.63 1.45 4.76 1.58 ;
 RECT 5.62 1.45 5.75 1.58 ;
 RECT 0.855 0.755 0.985 0.885 ;
 RECT 8.26 0.335 8.39 0.465 ;
 RECT 7.775 1.45 7.905 1.58 ;
 RECT 8.245 1.45 8.375 1.58 ;
 RECT 7.775 0.335 7.905 0.465 ;
 RECT 7.285 0.335 7.415 0.465 ;
 RECT 2.525 1.135 2.655 1.265 ;
 RECT 3.82 0.66 3.95 0.79 ;
 RECT 6.11 0.805 6.24 0.935 ;
 LAYER M1 ;
 RECT 0.85 0.995 0.99 1.87 ;
 RECT 0.85 0.7 0.99 0.855 ;
 RECT 1.71 1.26 1.85 1.35 ;
 RECT 1.53 1.12 1.85 1.26 ;
 RECT 0.85 0.855 1.67 0.995 ;
 RECT 1.53 0.995 1.67 1.12 ;
 RECT 3.66 1.155 3.8 1.7 ;
 RECT 4.625 1.155 4.765 1.675 ;
 RECT 5.615 1.155 5.755 1.71 ;
 RECT 3.66 1.015 5.755 1.155 ;
 RECT 1.81 1.685 1.95 2.36 ;
 RECT 1.81 0.57 1.95 0.835 ;
 RECT 2.02 0.975 2.16 1.13 ;
 RECT 2.02 1.27 2.16 1.545 ;
 RECT 1.81 0.835 2.16 0.975 ;
 RECT 1.81 1.545 2.16 1.685 ;
 RECT 2.475 1.095 2.705 1.13 ;
 RECT 2.475 1.27 2.705 1.305 ;
 RECT 1.99 1.13 2.705 1.27 ;
 RECT 4.14 0.265 4.28 0.735 ;
 RECT 5.095 1.35 5.235 1.945 ;
 RECT 6.035 0.975 6.175 1.945 ;
 RECT 4.14 0.765 6.29 0.875 ;
 RECT 4.14 0.735 6.175 0.765 ;
 RECT 6.035 0.875 6.29 0.975 ;
 RECT 5.095 1.945 6.175 2.085 ;
 END
END ISOLORAOX2

MACRO ISOLORAOX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 12.16 BY 2.88 ;
 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.795 1.07 6.935 1.845 ;
 RECT 6.795 0.22 6.935 0.79 ;
 RECT 6.56 1.01 6.935 1.07 ;
 RECT 6.56 0.79 6.935 0.87 ;
 RECT 7.77 1.01 7.91 1.845 ;
 RECT 7.77 0.22 7.91 0.87 ;
 RECT 8.755 1.01 8.895 1.845 ;
 RECT 8.755 0.22 8.895 0.87 ;
 RECT 9.73 1.01 9.87 1.845 ;
 RECT 9.73 0.22 9.87 0.87 ;
 RECT 6.56 0.87 9.87 1.01 ;
 END
 END Q

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 12.16 2.96 ;
 RECT 0.41 1.945 0.55 2.8 ;
 RECT 1.32 1.91 1.46 2.8 ;
 RECT 2.3 1.91 2.44 2.8 ;
 END
 END VDD

 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 4.15 2.48 10.9 2.62 ;
 RECT 4.15 1.35 4.29 2.48 ;
 RECT 10.75 1.105 10.89 2.48 ;
 RECT 6.315 1.345 6.455 2.48 ;
 RECT 7.265 1.345 7.405 2.48 ;
 RECT 8.24 1.345 8.38 2.48 ;
 RECT 9.225 1.345 9.365 2.48 ;
 RECT 10.2 1.345 10.34 2.48 ;
 END
 END VDDG

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 12.16 0.08 ;
 RECT 5.1 0.08 5.24 0.545 ;
 RECT 3.6 0.34 3.875 0.48 ;
 RECT 1.32 0.08 1.46 0.715 ;
 RECT 8.255 0.08 8.395 0.535 ;
 RECT 7.28 0.08 7.42 0.535 ;
 RECT 6.31 0.08 6.45 0.535 ;
 RECT 0.41 0.08 0.55 0.765 ;
 RECT 9.24 0.08 9.38 0.535 ;
 RECT 10.215 0.08 10.355 0.535 ;
 RECT 2.3 0.08 2.44 0.73 ;
 RECT 3.67 0.08 3.81 0.34 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.215 1.48 1.555 1.72 ;
 RECT 1.155 1.17 1.385 1.31 ;
 RECT 1.215 1.31 1.355 1.48 ;
 END
 END D

 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.635 0.62 4 0.875 ;
 END
 END ISO

 OBS
 LAYER PO ;
 RECT 1.575 1.12 1.895 1.125 ;
 RECT 1.575 0.315 1.675 1.12 ;
 RECT 1.575 1.225 1.895 1.35 ;
 RECT 1.575 1.35 1.675 2.74 ;
 RECT 2.085 0.315 2.185 1.125 ;
 RECT 2.085 1.225 2.185 2.74 ;
 RECT 1.575 1.125 2.185 1.225 ;
 RECT 1.105 0.44 1.205 1.125 ;
 RECT 1.105 1.125 1.385 1.355 ;
 RECT 1.105 1.355 1.205 2.24 ;
 RECT 5.085 1.95 5.185 2.305 ;
 RECT 3.3 1.145 3.4 2.305 ;
 RECT 5.365 1.015 5.465 1.85 ;
 RECT 4.88 1.85 5.465 1.95 ;
 RECT 4.88 0.125 4.98 1.85 ;
 RECT 2.475 1.095 3.4 1.145 ;
 RECT 2.475 1.145 2.705 1.305 ;
 RECT 2.565 1.045 3.4 1.095 ;
 RECT 3.3 2.305 5.185 2.405 ;
 RECT 3.925 0.83 4.025 1.025 ;
 RECT 3.925 1.125 4.025 1.95 ;
 RECT 4.405 1.125 4.505 1.95 ;
 RECT 3.925 0.09 4.025 0.62 ;
 RECT 3.77 0.62 4.025 0.83 ;
 RECT 3.925 1.025 4.505 1.125 ;
 RECT 9.985 0.095 10.085 0.845 ;
 RECT 9.985 0.945 10.085 1.95 ;
 RECT 9.505 0.095 9.605 0.845 ;
 RECT 9.505 0.945 9.605 1.95 ;
 RECT 8.53 0.095 8.63 0.845 ;
 RECT 8.53 0.945 8.63 1.95 ;
 RECT 9.01 0.095 9.11 0.845 ;
 RECT 9.01 0.945 9.11 1.95 ;
 RECT 6.57 0.095 6.67 0.845 ;
 RECT 6.57 0.945 6.67 1.95 ;
 RECT 7.05 0.095 7.15 0.845 ;
 RECT 7.05 0.945 7.15 1.95 ;
 RECT 7.545 0.095 7.645 0.845 ;
 RECT 7.545 0.945 7.645 1.95 ;
 RECT 8.025 0.095 8.125 0.845 ;
 RECT 8.025 0.945 8.125 1.95 ;
 RECT 6.06 0.765 6.29 0.845 ;
 RECT 6.06 0.945 6.29 0.975 ;
 RECT 6.06 0.845 10.085 0.945 ;
 LAYER CO ;
 RECT 0.855 1.69 0.985 1.82 ;
 RECT 0.855 0.755 0.985 0.885 ;
 RECT 4.145 0.345 4.275 0.475 ;
 RECT 6.32 1.45 6.45 1.58 ;
 RECT 3.665 1.45 3.795 1.58 ;
 RECT 6.8 1.45 6.93 1.58 ;
 RECT 1.325 0.535 1.455 0.665 ;
 RECT 5.1 1.45 5.23 1.58 ;
 RECT 7.27 1.45 7.4 1.58 ;
 RECT 6.8 0.335 6.93 0.465 ;
 RECT 3.675 0.345 3.805 0.475 ;
 RECT 0.415 0.305 0.545 0.435 ;
 RECT 7.775 1.45 7.905 1.58 ;
 RECT 1.815 1.645 1.945 1.775 ;
 RECT 0.415 0.565 0.545 0.695 ;
 RECT 1.815 1.645 1.945 1.775 ;
 RECT 1.815 1.95 1.945 2.08 ;
 RECT 5.105 0.345 5.235 0.475 ;
 RECT 0.415 2.015 0.545 2.145 ;
 RECT 5.62 1.45 5.75 1.58 ;
 RECT 10.755 1.175 10.885 1.305 ;
 RECT 1.815 0.62 1.945 0.75 ;
 RECT 1.715 1.17 1.845 1.3 ;
 RECT 4.63 1.45 4.76 1.58 ;
 RECT 2.305 1.96 2.435 2.09 ;
 RECT 9.735 0.335 9.865 0.465 ;
 RECT 10.22 0.335 10.35 0.465 ;
 RECT 9.245 0.335 9.375 0.465 ;
 RECT 9.23 1.45 9.36 1.58 ;
 RECT 8.76 0.335 8.89 0.465 ;
 RECT 10.205 1.45 10.335 1.58 ;
 RECT 8.76 1.45 8.89 1.58 ;
 RECT 9.735 1.45 9.865 1.58 ;
 RECT 10.755 1.435 10.885 1.565 ;
 RECT 7.775 0.335 7.905 0.465 ;
 RECT 1.325 1.96 1.455 2.09 ;
 RECT 1.205 1.175 1.335 1.305 ;
 RECT 4.155 1.45 4.285 1.58 ;
 RECT 0.415 2.275 0.545 2.405 ;
 RECT 2.305 0.55 2.435 0.68 ;
 RECT 8.26 0.335 8.39 0.465 ;
 RECT 8.245 1.45 8.375 1.58 ;
 RECT 7.285 0.335 7.415 0.465 ;
 RECT 6.315 0.335 6.445 0.465 ;
 RECT 2.525 1.135 2.655 1.265 ;
 RECT 3.82 0.66 3.95 0.79 ;
 RECT 6.11 0.805 6.24 0.935 ;
 LAYER M1 ;
 RECT 3.66 1.155 3.8 1.7 ;
 RECT 5.615 1.155 5.755 1.71 ;
 RECT 4.625 1.155 4.765 1.675 ;
 RECT 3.66 1.015 5.755 1.155 ;
 RECT 0.85 0.7 0.99 0.855 ;
 RECT 0.85 0.995 0.99 1.87 ;
 RECT 1.53 1.12 1.85 1.26 ;
 RECT 1.71 1.26 1.85 1.35 ;
 RECT 1.53 0.995 1.67 1.12 ;
 RECT 0.85 0.855 1.67 0.995 ;
 RECT 1.81 1.685 1.95 2.36 ;
 RECT 1.81 0.57 1.95 0.835 ;
 RECT 2.02 0.975 2.16 1.13 ;
 RECT 2.02 1.27 2.16 1.545 ;
 RECT 1.81 0.835 2.16 0.975 ;
 RECT 1.81 1.545 2.16 1.685 ;
 RECT 2.475 1.095 2.705 1.13 ;
 RECT 2.475 1.27 2.705 1.305 ;
 RECT 1.99 1.13 2.705 1.27 ;
 RECT 4.14 0.265 4.28 0.735 ;
 RECT 5.095 1.35 5.235 1.945 ;
 RECT 6.035 0.975 6.175 1.945 ;
 RECT 4.14 0.765 6.29 0.875 ;
 RECT 4.14 0.735 6.175 0.765 ;
 RECT 6.035 0.875 6.29 0.975 ;
 RECT 5.095 1.945 6.175 2.085 ;
 END
END ISOLORAOX4

MACRO ISOLORAOX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 16.32 BY 2.88 ;
 PIN VDDG
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 4.15 1.35 4.29 2.48 ;
 RECT 14.7 1.105 14.84 2.48 ;
 RECT 4.15 2.48 14.84 2.62 ;
 RECT 6.315 1.345 6.455 2.48 ;
 RECT 9.225 1.345 9.365 2.48 ;
 RECT 7.265 1.345 7.405 2.48 ;
 RECT 8.24 1.345 8.38 2.48 ;
 RECT 10.2 1.345 10.34 2.48 ;
 RECT 12.165 1.345 12.305 2.48 ;
 RECT 14.125 1.345 14.265 2.48 ;
 RECT 13.15 1.345 13.29 2.48 ;
 RECT 11.19 1.345 11.33 2.48 ;
 END
 END VDDG

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 16.32 2.96 ;
 RECT 0.41 1.945 0.55 2.8 ;
 RECT 1.32 1.91 1.46 2.8 ;
 RECT 2.3 1.91 2.44 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 6.795 1.07 6.935 1.845 ;
 RECT 6.795 0.22 6.935 0.79 ;
 RECT 6.56 1.01 6.935 1.07 ;
 RECT 6.56 0.79 6.935 0.87 ;
 RECT 7.77 1.01 7.91 1.845 ;
 RECT 7.77 0.22 7.91 0.87 ;
 RECT 9.73 1.01 9.87 1.845 ;
 RECT 9.73 0.22 9.87 0.87 ;
 RECT 8.755 1.01 8.895 1.845 ;
 RECT 8.755 0.22 8.895 0.87 ;
 RECT 11.695 1.01 11.835 1.845 ;
 RECT 11.695 0.22 11.835 0.87 ;
 RECT 10.72 1.01 10.86 1.845 ;
 RECT 10.72 0.22 10.86 0.87 ;
 RECT 12.68 1.01 12.82 1.845 ;
 RECT 12.68 0.22 12.82 0.87 ;
 RECT 13.655 1.01 13.795 1.845 ;
 RECT 13.655 0.22 13.795 0.87 ;
 RECT 6.56 0.87 13.795 1.01 ;
 END
 END Q

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 16.32 0.08 ;
 RECT 5.1 0.08 5.24 0.545 ;
 RECT 3.6 0.34 3.875 0.48 ;
 RECT 1.32 0.08 1.46 0.715 ;
 RECT 6.31 0.08 6.45 0.535 ;
 RECT 8.255 0.08 8.395 0.535 ;
 RECT 10.215 0.08 10.355 0.535 ;
 RECT 7.28 0.08 7.42 0.535 ;
 RECT 0.41 0.08 0.55 0.765 ;
 RECT 9.24 0.08 9.38 0.535 ;
 RECT 11.205 0.08 11.345 0.535 ;
 RECT 12.18 0.08 12.32 0.535 ;
 RECT 14.14 0.08 14.28 0.535 ;
 RECT 13.165 0.08 13.305 0.535 ;
 RECT 3.67 0.08 3.81 0.34 ;
 RECT 2.3 0.08 2.44 0.73 ;
 END
 END VSS

 PIN ISO
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.635 0.62 4 0.875 ;
 END
 END ISO

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.215 1.48 1.555 1.72 ;
 RECT 1.155 1.17 1.385 1.31 ;
 RECT 1.215 1.31 1.355 1.48 ;
 END
 END D

 OBS
 LAYER PO ;
 RECT 1.575 1.12 1.895 1.125 ;
 RECT 1.575 0.315 1.675 1.12 ;
 RECT 1.575 1.225 1.895 1.35 ;
 RECT 1.575 1.35 1.675 2.74 ;
 RECT 2.085 0.315 2.185 1.125 ;
 RECT 2.085 1.225 2.185 2.74 ;
 RECT 1.575 1.125 2.185 1.225 ;
 RECT 1.105 0.44 1.205 1.125 ;
 RECT 1.105 1.125 1.385 1.355 ;
 RECT 1.105 1.355 1.205 2.24 ;
 RECT 11.95 0.095 12.05 0.845 ;
 RECT 11.95 0.945 12.05 1.95 ;
 RECT 10.975 0.095 11.075 0.845 ;
 RECT 10.975 0.945 11.075 1.95 ;
 RECT 12.935 0.095 13.035 0.845 ;
 RECT 12.935 0.945 13.035 1.95 ;
 RECT 10.495 0.095 10.595 0.845 ;
 RECT 10.495 0.945 10.595 1.95 ;
 RECT 13.91 0.095 14.01 0.845 ;
 RECT 13.91 0.945 14.01 1.95 ;
 RECT 6.06 0.845 14.01 0.945 ;
 RECT 11.47 0.095 11.57 0.845 ;
 RECT 11.47 0.945 11.57 1.95 ;
 RECT 13.43 0.095 13.53 0.845 ;
 RECT 13.43 0.945 13.53 1.95 ;
 RECT 12.455 0.095 12.555 0.845 ;
 RECT 12.455 0.945 12.555 1.95 ;
 RECT 7.545 0.095 7.645 0.845 ;
 RECT 7.545 0.945 7.645 1.95 ;
 RECT 6.57 0.095 6.67 0.845 ;
 RECT 6.57 0.945 6.67 1.95 ;
 RECT 7.05 0.095 7.15 0.845 ;
 RECT 7.05 0.945 7.15 1.95 ;
 RECT 9.985 0.095 10.085 0.845 ;
 RECT 9.985 0.945 10.085 1.95 ;
 RECT 9.505 0.095 9.605 0.845 ;
 RECT 9.505 0.945 9.605 1.95 ;
 RECT 9.01 0.095 9.11 0.845 ;
 RECT 9.01 0.945 9.11 1.95 ;
 RECT 8.025 0.095 8.125 0.845 ;
 RECT 8.025 0.945 8.125 1.95 ;
 RECT 8.53 0.095 8.63 0.845 ;
 RECT 8.53 0.945 8.63 1.95 ;
 RECT 6.06 0.765 6.29 0.845 ;
 RECT 6.06 0.945 6.29 0.975 ;
 RECT 5.085 1.95 5.185 2.305 ;
 RECT 3.3 1.145 3.4 2.305 ;
 RECT 5.365 1.015 5.465 1.85 ;
 RECT 4.88 1.85 5.465 1.95 ;
 RECT 4.88 0.125 4.98 1.85 ;
 RECT 2.475 1.095 3.4 1.145 ;
 RECT 2.475 1.145 2.705 1.305 ;
 RECT 2.565 1.045 3.4 1.095 ;
 RECT 3.3 2.305 5.185 2.405 ;
 RECT 3.925 0.83 4.025 1.025 ;
 RECT 3.925 1.125 4.025 1.95 ;
 RECT 4.405 1.125 4.505 1.95 ;
 RECT 3.925 0.09 4.025 0.62 ;
 RECT 3.77 0.62 4.025 0.83 ;
 RECT 3.925 1.025 4.505 1.125 ;
 LAYER CO ;
 RECT 2.305 1.96 2.435 2.09 ;
 RECT 4.63 1.45 4.76 1.58 ;
 RECT 0.415 2.275 0.545 2.405 ;
 RECT 4.155 1.45 4.285 1.58 ;
 RECT 2.305 0.55 2.435 0.68 ;
 RECT 9.735 1.45 9.865 1.58 ;
 RECT 5.62 1.45 5.75 1.58 ;
 RECT 14.705 1.175 14.835 1.305 ;
 RECT 11.7 1.45 11.83 1.58 ;
 RECT 11.195 1.45 11.325 1.58 ;
 RECT 14.13 1.45 14.26 1.58 ;
 RECT 13.66 0.335 13.79 0.465 ;
 RECT 11.21 0.335 11.34 0.465 ;
 RECT 14.145 0.335 14.275 0.465 ;
 RECT 13.155 1.45 13.285 1.58 ;
 RECT 13.17 0.335 13.3 0.465 ;
 RECT 12.685 0.335 12.815 0.465 ;
 RECT 10.725 0.335 10.855 0.465 ;
 RECT 12.17 1.45 12.3 1.58 ;
 RECT 12.185 0.335 12.315 0.465 ;
 RECT 11.7 0.335 11.83 0.465 ;
 RECT 10.725 1.45 10.855 1.58 ;
 RECT 12.685 1.45 12.815 1.58 ;
 RECT 13.66 1.45 13.79 1.58 ;
 RECT 6.315 0.335 6.445 0.465 ;
 RECT 3.675 0.345 3.805 0.475 ;
 RECT 0.415 0.305 0.545 0.435 ;
 RECT 1.815 0.62 1.945 0.75 ;
 RECT 7.775 1.45 7.905 1.58 ;
 RECT 4.145 0.345 4.275 0.475 ;
 RECT 0.415 0.565 0.545 0.695 ;
 RECT 5.105 0.345 5.235 0.475 ;
 RECT 7.285 0.335 7.415 0.465 ;
 RECT 3.665 1.45 3.795 1.58 ;
 RECT 7.27 1.45 7.4 1.58 ;
 RECT 1.815 1.645 1.945 1.775 ;
 RECT 6.8 0.335 6.93 0.465 ;
 RECT 1.325 0.535 1.455 0.665 ;
 RECT 6.11 0.805 6.24 0.935 ;
 RECT 2.525 1.135 2.655 1.265 ;
 RECT 3.82 0.66 3.95 0.79 ;
 RECT 0.415 2.015 0.545 2.145 ;
 RECT 0.855 1.69 0.985 1.82 ;
 RECT 0.855 0.755 0.985 0.885 ;
 RECT 6.32 1.45 6.45 1.58 ;
 RECT 1.815 1.95 1.945 2.08 ;
 RECT 8.245 1.45 8.375 1.58 ;
 RECT 10.205 1.45 10.335 1.58 ;
 RECT 10.22 0.335 10.35 0.465 ;
 RECT 8.76 0.335 8.89 0.465 ;
 RECT 9.23 1.45 9.36 1.58 ;
 RECT 7.775 0.335 7.905 0.465 ;
 RECT 6.8 1.45 6.93 1.58 ;
 RECT 1.815 1.645 1.945 1.775 ;
 RECT 9.245 0.335 9.375 0.465 ;
 RECT 14.705 1.435 14.835 1.565 ;
 RECT 9.735 0.335 9.865 0.465 ;
 RECT 5.1 1.45 5.23 1.58 ;
 RECT 1.325 1.96 1.455 2.09 ;
 RECT 8.76 1.45 8.89 1.58 ;
 RECT 1.205 1.175 1.335 1.305 ;
 RECT 8.26 0.335 8.39 0.465 ;
 RECT 1.715 1.17 1.845 1.3 ;
 LAYER M1 ;
 RECT 3.66 1.155 3.8 1.7 ;
 RECT 5.615 1.155 5.755 1.71 ;
 RECT 4.625 1.155 4.765 1.675 ;
 RECT 3.66 1.015 5.755 1.155 ;
 RECT 0.85 0.7 0.99 0.855 ;
 RECT 0.85 0.995 0.99 1.87 ;
 RECT 1.53 1.12 1.85 1.26 ;
 RECT 1.71 1.26 1.85 1.35 ;
 RECT 1.53 0.995 1.67 1.12 ;
 RECT 0.85 0.855 1.67 0.995 ;
 RECT 4.14 0.265 4.28 0.735 ;
 RECT 6.035 0.875 6.29 0.975 ;
 RECT 6.035 0.975 6.175 1.945 ;
 RECT 5.095 1.35 5.235 1.945 ;
 RECT 4.14 0.765 6.29 0.875 ;
 RECT 4.14 0.735 6.175 0.765 ;
 RECT 5.095 1.945 6.175 2.085 ;
 RECT 1.81 1.685 1.95 2.36 ;
 RECT 1.81 0.57 1.95 0.835 ;
 RECT 2.02 0.975 2.16 1.13 ;
 RECT 2.02 1.27 2.16 1.545 ;
 RECT 1.81 0.835 2.16 0.975 ;
 RECT 1.81 1.545 2.16 1.685 ;
 RECT 2.475 1.095 2.705 1.13 ;
 RECT 2.475 1.27 2.705 1.305 ;
 RECT 1.99 1.13 2.705 1.27 ;
 END
END ISOLORAOX8

MACRO LSDNENCLSSX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.985 0.825 1.255 1.095 ;
 END
 END D

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.265 0.655 2.535 0.925 ;
 END
 END ENB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 0.325 0.08 0.465 0.765 ;
 RECT 2.525 0.08 2.665 0.515 ;
 RECT 1.585 0.08 1.725 0.515 ;
 RECT 1.205 0.08 1.345 0.545 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 1.585 1.69 1.725 2.8 ;
 RECT 0.325 1.505 0.465 2.8 ;
 RECT 1.205 1.63 1.345 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.525 1.31 2.85 1.41 ;
 RECT 1.985 1.17 2.85 1.31 ;
 RECT 1.985 0.33 2.26 0.47 ;
 RECT 2.525 1.41 2.665 2.29 ;
 RECT 1.985 0.47 2.125 1.17 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 0.99 0.125 1.09 0.845 ;
 RECT 0.99 0.845 1.235 1.075 ;
 RECT 0.99 1.075 1.09 2.195 ;
 RECT 2.31 0.905 2.41 2.645 ;
 RECT 2.31 0.115 2.41 0.675 ;
 RECT 2.285 0.675 2.515 0.905 ;
 RECT 1.84 0.115 1.94 0.78 ;
 RECT 1.595 0.78 1.94 1.01 ;
 RECT 1.84 1.01 1.94 2.645 ;
 LAYER CO ;
 RECT 1.645 0.83 1.775 0.96 ;
 RECT 0.33 0.325 0.46 0.455 ;
 RECT 1.59 0.335 1.72 0.465 ;
 RECT 2.335 0.725 2.465 0.855 ;
 RECT 1.055 0.895 1.185 1.025 ;
 RECT 1.21 1.7 1.34 1.83 ;
 RECT 1.59 2.1 1.72 2.23 ;
 RECT 0.74 1.7 0.87 1.83 ;
 RECT 2.53 2.09 2.66 2.22 ;
 RECT 0.33 1.555 0.46 1.685 ;
 RECT 0.33 0.585 0.46 0.715 ;
 RECT 1.59 1.82 1.72 1.95 ;
 RECT 2.53 1.815 2.66 1.945 ;
 RECT 0.33 1.815 0.46 1.945 ;
 RECT 2.53 0.335 2.66 0.465 ;
 RECT 0.74 0.345 0.87 0.475 ;
 RECT 0.33 2.075 0.46 2.205 ;
 RECT 2.06 0.335 2.19 0.465 ;
 RECT 1.21 0.345 1.34 0.475 ;
 LAYER M1 ;
 RECT 0.735 0.275 0.875 0.47 ;
 RECT 0.695 0.47 0.875 0.61 ;
 RECT 0.695 0.61 0.835 1.235 ;
 RECT 0.695 1.235 0.875 1.375 ;
 RECT 0.735 1.375 0.875 2.005 ;
 RECT 1.64 0.755 1.78 1.37 ;
 RECT 0.735 1.235 1.785 1.375 ;
 END
END LSDNENCLSSX1

MACRO LSDNENCLSSX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 5.44 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 5.44 2.96 ;
 RECT 0.46 1.49 0.6 2.8 ;
 RECT 1.77 1.59 1.91 2.8 ;
 RECT 4.945 1.93 5.085 2.8 ;
 RECT 3.59 1.655 3.73 2.8 ;
 RECT 4.535 1.72 4.675 2.8 ;
 RECT 1.39 1.615 1.53 2.8 ;
 END
 END VDD

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.45 0.81 2.72 1.08 ;
 END
 END ENB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.305 0.825 1.575 1.095 ;
 END
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 5.44 0.08 ;
 RECT 1.77 0.08 1.91 0.5 ;
 RECT 2.71 0.08 2.85 0.5 ;
 RECT 0.415 0.08 0.555 0.75 ;
 RECT 4.945 0.08 5.085 0.76 ;
 RECT 3.595 0.08 3.735 0.525 ;
 RECT 4.54 0.08 4.68 0.585 ;
 RECT 1.39 0.08 1.53 0.53 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.94 1.7 4.26 2.075 ;
 RECT 4.065 0.5 4.205 1.7 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 1.175 0.845 1.555 1.075 ;
 RECT 1.175 0.11 1.275 0.845 ;
 RECT 1.175 1.075 1.275 2.34 ;
 RECT 3.66 1.27 3.95 1.4 ;
 RECT 3.66 1.17 4.42 1.27 ;
 RECT 4.32 0.095 4.42 1.17 ;
 RECT 4.32 1.27 4.42 2.78 ;
 RECT 3.85 0.095 3.95 1.17 ;
 RECT 3.85 1.4 3.95 2.78 ;
 RECT 2.495 0.1 2.595 0.83 ;
 RECT 2.495 1.06 2.595 2.63 ;
 RECT 2.47 0.83 2.7 1.06 ;
 RECT 2.025 0.98 2.125 2.63 ;
 RECT 2.025 0.1 2.125 0.75 ;
 RECT 1.835 0.75 2.125 0.98 ;
 RECT 3.22 2.265 3.475 2.42 ;
 RECT 3.22 2.42 3.47 2.495 ;
 RECT 3.375 0.095 3.475 2.265 ;
 LAYER CO ;
 RECT 1.775 1.9 1.905 2.03 ;
 RECT 1.775 1.64 1.905 1.77 ;
 RECT 2.715 2.075 2.845 2.205 ;
 RECT 1.775 0.32 1.905 0.45 ;
 RECT 0.925 1.685 1.055 1.815 ;
 RECT 0.465 1.8 0.595 1.93 ;
 RECT 2.52 0.88 2.65 1.01 ;
 RECT 1.395 1.685 1.525 1.815 ;
 RECT 2.715 1.8 2.845 1.93 ;
 RECT 1.775 2.16 1.905 2.29 ;
 RECT 0.42 0.57 0.55 0.7 ;
 RECT 3.6 0.325 3.73 0.455 ;
 RECT 4.54 2.305 4.67 2.435 ;
 RECT 4.54 1.79 4.67 1.92 ;
 RECT 2.245 0.32 2.375 0.45 ;
 RECT 0.465 2.06 0.595 2.19 ;
 RECT 1.395 0.33 1.525 0.46 ;
 RECT 1.375 0.895 1.505 1.025 ;
 RECT 0.465 1.54 0.595 1.67 ;
 RECT 2.715 0.32 2.845 0.45 ;
 RECT 0.42 0.31 0.55 0.44 ;
 RECT 0.925 0.33 1.055 0.46 ;
 RECT 1.89 0.81 2.02 0.94 ;
 RECT 3.27 2.31 3.4 2.44 ;
 RECT 3.12 1.81 3.25 1.94 ;
 RECT 4.07 0.565 4.2 0.695 ;
 RECT 4.95 0.3 5.08 0.43 ;
 RECT 4.545 0.385 4.675 0.515 ;
 RECT 3.595 2.305 3.725 2.435 ;
 RECT 3.125 0.325 3.255 0.455 ;
 RECT 4.07 1.61 4.2 1.74 ;
 RECT 4.07 1.91 4.2 2.04 ;
 RECT 3.12 1.54 3.25 1.67 ;
 RECT 4.95 2 5.08 2.13 ;
 RECT 4.95 2.26 5.08 2.39 ;
 RECT 3.71 1.225 3.84 1.355 ;
 RECT 3.595 1.73 3.725 1.86 ;
 RECT 4.95 0.56 5.08 0.69 ;
 LAYER M1 ;
 RECT 3.12 0.255 3.26 1.22 ;
 RECT 3.115 1.36 3.255 2.01 ;
 RECT 3.115 1.22 3.89 1.36 ;
 RECT 0.92 0.26 1.06 1.24 ;
 RECT 0.92 1.38 1.06 1.89 ;
 RECT 0.92 1.24 2.025 1.375 ;
 RECT 0.92 1.375 2.02 1.38 ;
 RECT 1.885 0.76 2.025 1.24 ;
 RECT 2.17 0.48 2.32 0.615 ;
 RECT 2.18 0.455 2.32 0.48 ;
 RECT 2.17 0.615 2.31 1.23 ;
 RECT 2.18 0.315 2.445 0.455 ;
 RECT 2.71 2.305 3.45 2.445 ;
 RECT 2.71 1.37 2.85 2.305 ;
 RECT 2.17 1.23 2.85 1.37 ;
 END
END LSDNENCLSSX2

MACRO LSDNENCLSSX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.72 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.72 0.08 ;
 RECT 1.41 0.08 1.55 0.535 ;
 RECT 6.195 0.08 6.335 0.89 ;
 RECT 0.92 0.08 1.06 0.685 ;
 RECT 3.635 0.08 3.775 0.785 ;
 RECT 2.35 0.08 2.49 0.535 ;
 RECT 2.745 0.08 2.885 0.525 ;
 RECT 4.63 0.08 4.77 0.785 ;
 RECT 5.645 0.08 5.785 0.785 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.72 2.96 ;
 RECT 1.41 1.42 1.55 2.8 ;
 RECT 0.92 1.64 1.06 2.8 ;
 RECT 6.195 1.935 6.335 2.8 ;
 RECT 3.635 1.735 3.775 2.8 ;
 RECT 2.745 1.565 2.885 2.8 ;
 RECT 4.635 1.735 4.775 2.8 ;
 RECT 5.65 1.735 5.79 2.8 ;
 END
 END VDD

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.175 0.745 2.495 1.105 ;
 END
 END ENB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.725 1.125 1.11 1.46 ;
 END
 END D

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.115 1.1 5.275 1.11 ;
 RECT 4.115 0.97 5.325 1.1 ;
 RECT 5.135 0.275 5.275 0.83 ;
 RECT 4.115 1.11 4.255 2.585 ;
 RECT 5.135 1.11 5.275 2.585 ;
 RECT 5.135 0.83 5.325 0.97 ;
 RECT 4.115 0.275 4.255 0.97 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 0.695 0.255 0.795 1.125 ;
 RECT 0.695 1.125 0.97 1.355 ;
 RECT 0.695 1.355 0.795 2.17 ;
 RECT 1.665 0.105 1.765 0.8 ;
 RECT 1.48 0.8 1.765 1.03 ;
 RECT 1.665 1.03 1.765 2.77 ;
 RECT 3 0.105 3.1 1.14 ;
 RECT 3 1.37 3.1 2.77 ;
 RECT 2.895 1.14 3.125 1.37 ;
 RECT 5.425 0.105 5.525 1.23 ;
 RECT 5.425 1.33 5.525 2.77 ;
 RECT 4.91 0.105 5.01 1.23 ;
 RECT 4.91 1.33 5.01 2.77 ;
 RECT 4.39 0.105 4.49 1.23 ;
 RECT 4.39 1.33 4.49 2.77 ;
 RECT 3.785 1.14 4.015 1.23 ;
 RECT 3.785 1.33 4.015 1.37 ;
 RECT 3.785 1.23 5.525 1.33 ;
 RECT 3.89 0.105 3.99 1.14 ;
 RECT 3.89 1.37 3.99 2.77 ;
 RECT 2.135 0.745 2.455 1.09 ;
 RECT 2.135 0.105 2.235 0.745 ;
 RECT 2.135 1.09 2.235 2.77 ;
 LAYER CO ;
 RECT 0.44 0.505 0.57 0.635 ;
 RECT 0.925 0.505 1.055 0.635 ;
 RECT 6.2 2.005 6.33 2.135 ;
 RECT 6.2 2.265 6.33 2.395 ;
 RECT 6.2 0.69 6.33 0.82 ;
 RECT 6.2 0.43 6.33 0.56 ;
 RECT 4.12 2.065 4.25 2.195 ;
 RECT 4.12 0.585 4.25 0.715 ;
 RECT 4.12 2.345 4.25 2.475 ;
 RECT 2.355 2.08 2.485 2.21 ;
 RECT 1.415 1.81 1.545 1.94 ;
 RECT 5.655 2.345 5.785 2.475 ;
 RECT 5.655 1.805 5.785 1.935 ;
 RECT 5.655 2.065 5.785 2.195 ;
 RECT 5.65 0.325 5.78 0.455 ;
 RECT 5.65 0.585 5.78 0.715 ;
 RECT 5.14 0.325 5.27 0.455 ;
 RECT 5.14 1.545 5.27 1.675 ;
 RECT 5.14 1.805 5.27 1.935 ;
 RECT 5.14 2.065 5.27 2.195 ;
 RECT 5.14 0.585 5.27 0.715 ;
 RECT 5.14 2.345 5.27 2.475 ;
 RECT 4.64 2.065 4.77 2.195 ;
 RECT 4.64 2.345 4.77 2.475 ;
 RECT 4.635 0.325 4.765 0.455 ;
 RECT 4.635 0.585 4.765 0.715 ;
 RECT 4.64 1.805 4.77 1.935 ;
 RECT 3.23 0.325 3.36 0.455 ;
 RECT 3.23 1.545 3.36 1.675 ;
 RECT 3.23 1.805 3.36 1.935 ;
 RECT 2.945 1.19 3.075 1.32 ;
 RECT 2.75 0.325 2.88 0.455 ;
 RECT 2.75 1.725 2.88 1.855 ;
 RECT 2.355 0.335 2.485 0.465 ;
 RECT 1.415 0.335 1.545 0.465 ;
 RECT 3.64 0.325 3.77 0.455 ;
 RECT 3.64 0.585 3.77 0.715 ;
 RECT 3.64 1.805 3.77 1.935 ;
 RECT 3.64 2.065 3.77 2.195 ;
 RECT 3.64 2.345 3.77 2.475 ;
 RECT 2.285 0.875 2.415 1.005 ;
 RECT 1.415 2.09 1.545 2.22 ;
 RECT 3.835 1.19 3.965 1.32 ;
 RECT 1.53 0.85 1.66 0.98 ;
 RECT 2.355 1.805 2.485 1.935 ;
 RECT 4.12 1.545 4.25 1.675 ;
 RECT 1.885 0.335 2.015 0.465 ;
 RECT 4.12 0.325 4.25 0.455 ;
 RECT 1.415 1.545 1.545 1.675 ;
 RECT 4.12 1.805 4.25 1.935 ;
 RECT 0.44 1.69 0.57 1.82 ;
 RECT 0.925 1.69 1.055 1.82 ;
 RECT 0.79 1.175 0.92 1.305 ;
 LAYER M1 ;
 RECT 0.435 0.435 0.575 0.845 ;
 RECT 0.435 0.985 0.575 1.87 ;
 RECT 0.435 0.845 1.73 0.985 ;
 RECT 3.225 0.275 3.365 1.26 ;
 RECT 3.225 1.4 3.365 2.095 ;
 RECT 3.225 1.26 3.975 1.4 ;
 RECT 3.82 1.14 3.975 1.26 ;
 RECT 2.35 1.4 2.49 2.28 ;
 RECT 1.88 0.265 2.02 1.26 ;
 RECT 1.88 1.26 3.085 1.37 ;
 RECT 2.93 1.14 3.085 1.26 ;
 RECT 1.88 1.37 3.075 1.4 ;
 END
END LSDNENCLSSX4

MACRO LSDNENCLSSX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 9.6 BY 2.88 ;
 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.985 0.825 1.255 1.095 ;
 END
 END D

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.335 0.825 2.605 1.095 ;
 END
 END ENB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 9.6 0.08 ;
 RECT 0.325 0.08 0.465 0.765 ;
 RECT 1.205 0.08 1.345 0.545 ;
 RECT 1.585 0.08 1.725 0.515 ;
 RECT 2.525 0.08 2.665 0.515 ;
 RECT 3.56 0.08 3.7 0.58 ;
 RECT 4.685 0.08 4.825 0.6 ;
 RECT 5.675 0.08 5.815 0.6 ;
 RECT 6.64 0.08 6.78 0.6 ;
 RECT 7.61 0.08 7.75 0.6 ;
 RECT 8.565 0.08 8.705 0.6 ;
 RECT 8.995 0.08 9.135 0.9 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 9.6 2.96 ;
 RECT 8.995 1.945 9.135 2.8 ;
 RECT 3.565 1.735 3.705 2.8 ;
 RECT 4.725 1.735 4.865 2.8 ;
 RECT 5.675 1.735 5.815 2.8 ;
 RECT 6.64 1.735 6.78 2.8 ;
 RECT 7.61 1.735 7.75 2.8 ;
 RECT 8.565 1.735 8.705 2.8 ;
 RECT 1.585 1.69 1.725 2.8 ;
 RECT 1.205 1.63 1.345 2.8 ;
 RECT 0.325 1.505 0.465 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 7.9 1.245 8.39 1.455 ;
 RECT 8.095 1.455 8.235 2.36 ;
 RECT 5.205 1.105 8.39 1.245 ;
 RECT 5.205 1.245 5.345 2.36 ;
 RECT 6.17 1.245 6.31 2.36 ;
 RECT 7.14 1.245 7.28 2.36 ;
 RECT 7.9 1.045 8.39 1.105 ;
 RECT 5.205 0.41 5.345 1.105 ;
 RECT 6.17 0.41 6.31 1.105 ;
 RECT 7.14 0.41 7.28 1.105 ;
 RECT 8.095 0.41 8.235 1.045 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 0.99 0.125 1.09 0.845 ;
 RECT 0.99 0.845 1.235 1.075 ;
 RECT 0.99 1.075 1.09 2.195 ;
 RECT 1.84 0.115 1.94 0.78 ;
 RECT 1.595 0.78 1.94 1.01 ;
 RECT 1.84 1.01 1.94 2.645 ;
 RECT 8.35 0.21 8.45 2.765 ;
 RECT 7.88 0.11 8.45 0.21 ;
 RECT 7.88 0.21 7.98 2.665 ;
 RECT 7.395 2.665 7.98 2.765 ;
 RECT 7.395 0.21 7.495 2.665 ;
 RECT 6.925 0.11 7.495 0.21 ;
 RECT 6.925 0.21 7.025 2.665 ;
 RECT 6.425 2.665 7.025 2.765 ;
 RECT 6.425 0.21 6.525 2.665 ;
 RECT 5.955 0.11 6.525 0.21 ;
 RECT 5.955 0.21 6.055 2.665 ;
 RECT 5.46 2.665 6.055 2.765 ;
 RECT 5.46 0.21 5.56 2.665 ;
 RECT 4.99 0.11 5.56 0.21 ;
 RECT 4.99 0.21 5.09 0.955 ;
 RECT 4.86 0.955 5.09 1.185 ;
 RECT 4.99 1.185 5.09 2.765 ;
 RECT 2.87 1.125 3.1 1.235 ;
 RECT 2.87 1.025 4.55 1.125 ;
 RECT 4.45 0.11 4.55 1.025 ;
 RECT 3.82 0.11 3.92 1.025 ;
 RECT 3.34 0.11 3.44 1.025 ;
 RECT 4.45 1.125 4.55 2.79 ;
 RECT 3.82 1.125 3.92 2.79 ;
 RECT 3.34 1.125 3.44 2.79 ;
 RECT 2.31 0.115 2.41 0.855 ;
 RECT 2.31 0.855 2.595 1.065 ;
 RECT 2.31 1.065 2.41 2.645 ;
 LAYER CO ;
 RECT 2.53 0.335 2.66 0.465 ;
 RECT 2.53 2.09 2.66 2.22 ;
 RECT 2.06 0.335 2.19 0.465 ;
 RECT 1.59 2.1 1.72 2.23 ;
 RECT 0.33 2.075 0.46 2.205 ;
 RECT 0.33 1.815 0.46 1.945 ;
 RECT 4.155 0.48 4.285 0.61 ;
 RECT 3.085 2.32 3.215 2.45 ;
 RECT 3.08 0.4 3.21 0.53 ;
 RECT 2.53 1.815 2.66 1.945 ;
 RECT 4.155 1.76 4.285 1.89 ;
 RECT 3.57 2.32 3.7 2.45 ;
 RECT 3.57 1.805 3.7 1.935 ;
 RECT 0.74 1.7 0.87 1.83 ;
 RECT 4.155 2.145 4.285 2.275 ;
 RECT 1.59 0.335 1.72 0.465 ;
 RECT 3.565 0.4 3.695 0.53 ;
 RECT 0.33 0.325 0.46 0.455 ;
 RECT 1.59 1.82 1.72 1.95 ;
 RECT 1.21 1.7 1.34 1.83 ;
 RECT 3.085 1.805 3.215 1.935 ;
 RECT 1.055 0.895 1.185 1.025 ;
 RECT 1.21 0.345 1.34 0.475 ;
 RECT 1.645 0.83 1.775 0.96 ;
 RECT 0.33 1.555 0.46 1.685 ;
 RECT 0.33 0.585 0.46 0.715 ;
 RECT 0.74 0.345 0.87 0.475 ;
 RECT 5.21 0.48 5.34 0.61 ;
 RECT 4.91 1.005 5.04 1.135 ;
 RECT 6.175 2.145 6.305 2.275 ;
 RECT 6.645 2.32 6.775 2.45 ;
 RECT 4.69 0.4 4.82 0.53 ;
 RECT 6.645 1.805 6.775 1.935 ;
 RECT 5.68 1.805 5.81 1.935 ;
 RECT 8.1 0.48 8.23 0.61 ;
 RECT 7.145 1.76 7.275 1.89 ;
 RECT 5.68 0.4 5.81 0.53 ;
 RECT 7.145 2.145 7.275 2.275 ;
 RECT 7.145 0.48 7.275 0.61 ;
 RECT 5.21 2.145 5.34 2.275 ;
 RECT 7.615 2.32 7.745 2.45 ;
 RECT 6.645 0.4 6.775 0.53 ;
 RECT 4.73 2.32 4.86 2.45 ;
 RECT 8.1 2.145 8.23 2.275 ;
 RECT 4.73 1.805 4.86 1.935 ;
 RECT 8.1 1.76 8.23 1.89 ;
 RECT 5.68 2.32 5.81 2.45 ;
 RECT 7.615 1.805 7.745 1.935 ;
 RECT 6.175 0.48 6.305 0.61 ;
 RECT 6.175 1.76 6.305 1.89 ;
 RECT 5.21 1.76 5.34 1.89 ;
 RECT 7.615 0.4 7.745 0.53 ;
 RECT 9 0.7 9.13 0.83 ;
 RECT 8.57 2.32 8.7 2.45 ;
 RECT 9 0.44 9.13 0.57 ;
 RECT 8.57 0.4 8.7 0.53 ;
 RECT 9 2.015 9.13 2.145 ;
 RECT 9 2.275 9.13 2.405 ;
 RECT 8.57 1.805 8.7 1.935 ;
 RECT 2.92 1.065 3.05 1.195 ;
 RECT 2.415 0.895 2.545 1.025 ;
 LAYER M1 ;
 RECT 0.735 0.275 0.875 0.47 ;
 RECT 0.695 0.47 0.875 0.61 ;
 RECT 0.695 0.61 0.835 1.235 ;
 RECT 0.735 1.375 0.875 2.005 ;
 RECT 1.64 0.755 1.78 1.235 ;
 RECT 0.695 1.235 1.785 1.375 ;
 RECT 4.15 0.41 4.29 1.335 ;
 RECT 4.435 1.15 4.575 1.335 ;
 RECT 4.15 1.475 4.29 2.36 ;
 RECT 3.245 1.335 4.575 1.475 ;
 RECT 3.075 0.33 3.215 0.72 ;
 RECT 3.075 0.72 3.385 0.86 ;
 RECT 3.245 0.86 3.385 1.335 ;
 RECT 3.245 1.475 3.385 1.545 ;
 RECT 3.08 1.545 3.385 1.69 ;
 RECT 3.08 1.69 3.22 2.52 ;
 RECT 4.905 0.935 5.045 1.01 ;
 RECT 4.905 1.15 5.045 1.205 ;
 RECT 4.435 1.01 5.045 1.15 ;
 RECT 2.055 0.265 2.195 1.245 ;
 RECT 2.87 1.235 3.03 1.245 ;
 RECT 2.525 1.385 2.665 2.29 ;
 RECT 2.055 1.245 3.03 1.385 ;
 RECT 2.87 1.025 3.1 1.235 ;
 END
END LSDNENCLSSX8

MACRO LSDNENSSX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.84 BY 2.88 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.475 0.755 1.835 1.14 ;
 END
 END ENB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.265 0.825 2.535 1.095 ;
 END
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.84 0.08 ;
 RECT 0.325 0.08 0.465 0.765 ;
 RECT 2.525 0.08 2.665 0.515 ;
 RECT 1.585 0.08 1.725 0.515 ;
 RECT 2.915 0.08 3.055 0.705 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.84 2.96 ;
 RECT 1.585 1.69 1.725 2.8 ;
 RECT 0.325 1.505 0.465 2.8 ;
 RECT 2.915 1.745 3.055 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 3.405 1.08 3.545 2.595 ;
 RECT 3.165 0.84 3.545 1.08 ;
 RECT 3.405 0.285 3.545 0.84 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 2.31 0.115 2.41 0.845 ;
 RECT 2.31 1.075 2.41 2.645 ;
 RECT 2.285 0.845 2.515 1.075 ;
 RECT 2.765 1.12 3.28 1.35 ;
 RECT 3.18 0.115 3.28 1.12 ;
 RECT 3.18 1.35 3.28 2.78 ;
 RECT 1.84 0.115 1.94 0.78 ;
 RECT 1.595 0.78 1.94 1.01 ;
 RECT 1.84 1.01 1.94 2.645 ;
 LAYER CO ;
 RECT 1.645 0.83 1.775 0.96 ;
 RECT 3.41 0.595 3.54 0.725 ;
 RECT 3.41 0.335 3.54 0.465 ;
 RECT 3.41 1.815 3.54 1.945 ;
 RECT 3.41 1.555 3.54 1.685 ;
 RECT 3.41 2.355 3.54 2.485 ;
 RECT 3.41 2.075 3.54 2.205 ;
 RECT 0.33 0.325 0.46 0.455 ;
 RECT 2.815 1.17 2.945 1.3 ;
 RECT 1.59 0.335 1.72 0.465 ;
 RECT 2.335 0.895 2.465 1.025 ;
 RECT 2.92 2.355 3.05 2.485 ;
 RECT 2.92 1.815 3.05 1.945 ;
 RECT 1.59 2.1 1.72 2.23 ;
 RECT 2.92 0.335 3.05 0.465 ;
 RECT 2.92 2.075 3.05 2.205 ;
 RECT 2.53 2.09 2.66 2.22 ;
 RECT 0.33 1.555 0.46 1.685 ;
 RECT 0.33 0.585 0.46 0.715 ;
 RECT 1.59 1.82 1.72 1.95 ;
 RECT 2.53 1.815 2.66 1.945 ;
 RECT 0.33 1.815 0.46 1.945 ;
 RECT 2.53 0.335 2.66 0.465 ;
 RECT 0.33 2.075 0.46 2.205 ;
 RECT 2.06 0.335 2.19 0.465 ;
 LAYER M1 ;
 RECT 1.985 0.33 2.26 0.47 ;
 RECT 1.985 0.47 2.125 0.63 ;
 RECT 1.985 0.495 2.125 1.245 ;
 RECT 2.525 1.305 2.85 1.385 ;
 RECT 1.985 1.245 2.66 1.385 ;
 RECT 2.525 1.245 2.665 2.29 ;
 RECT 2.71 1.165 3.015 1.245 ;
 RECT 2.525 1.245 3.015 1.305 ;
 END
END LSDNENSSX1

MACRO LSDNENSSX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 6.4 BY 2.88 ;
 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 6.4 2.96 ;
 RECT 0.46 1.49 0.6 2.8 ;
 RECT 1.77 1.59 1.91 2.8 ;
 RECT 5.785 1.93 5.925 2.8 ;
 RECT 4.43 1.655 4.57 2.8 ;
 RECT 5.375 1.72 5.515 2.8 ;
 RECT 3.1 1.73 3.24 2.8 ;
 END
 END VDD

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.45 0.81 2.72 1.08 ;
 END
 END D

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.76 0.75 2.03 1.02 ;
 END
 END ENB

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 6.4 0.08 ;
 RECT 1.77 0.08 1.91 0.5 ;
 RECT 2.71 0.08 2.85 0.5 ;
 RECT 0.415 0.08 0.555 0.75 ;
 RECT 5.785 0.08 5.925 0.76 ;
 RECT 4.435 0.08 4.575 0.525 ;
 RECT 5.38 0.08 5.52 0.585 ;
 RECT 3.1 0.08 3.24 0.775 ;
 END
 END VSS

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.78 1.7 5.1 2.075 ;
 RECT 4.905 0.5 5.045 1.7 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 4.5 1.27 4.79 1.4 ;
 RECT 4.5 1.17 5.26 1.27 ;
 RECT 5.16 0.095 5.26 1.17 ;
 RECT 5.16 1.27 5.26 2.78 ;
 RECT 4.69 0.095 4.79 1.17 ;
 RECT 4.69 1.4 4.79 2.78 ;
 RECT 2.495 0.1 2.595 0.83 ;
 RECT 2.495 1.06 2.595 2.63 ;
 RECT 2.47 0.83 2.7 1.06 ;
 RECT 2.025 0.98 2.125 2.63 ;
 RECT 2.025 0.1 2.125 0.75 ;
 RECT 1.835 0.75 2.125 0.98 ;
 RECT 4.06 2.265 4.315 2.42 ;
 RECT 4.06 2.42 4.31 2.495 ;
 RECT 4.215 0.095 4.315 2.265 ;
 RECT 3.185 1.105 3.465 1.335 ;
 RECT 3.365 0.1 3.465 1.105 ;
 RECT 3.365 1.335 3.465 2.765 ;
 LAYER CO ;
 RECT 3.235 1.155 3.365 1.285 ;
 RECT 0.465 1.8 0.595 1.93 ;
 RECT 2.52 0.88 2.65 1.01 ;
 RECT 2.715 1.8 2.845 1.93 ;
 RECT 1.775 2.16 1.905 2.29 ;
 RECT 3.105 2.34 3.235 2.47 ;
 RECT 0.42 0.57 0.55 0.7 ;
 RECT 4.44 0.325 4.57 0.455 ;
 RECT 5.38 2.305 5.51 2.435 ;
 RECT 5.38 1.79 5.51 1.92 ;
 RECT 3.105 2.06 3.235 2.19 ;
 RECT 2.245 0.32 2.375 0.45 ;
 RECT 0.465 2.06 0.595 2.19 ;
 RECT 3.595 1.54 3.725 1.67 ;
 RECT 3.105 1.8 3.235 1.93 ;
 RECT 3.595 1.8 3.725 1.93 ;
 RECT 0.465 1.54 0.595 1.67 ;
 RECT 2.715 0.32 2.845 0.45 ;
 RECT 0.42 0.31 0.55 0.44 ;
 RECT 3.595 0.58 3.725 0.71 ;
 RECT 3.595 2.34 3.725 2.47 ;
 RECT 1.89 0.81 2.02 0.94 ;
 RECT 4.11 2.31 4.24 2.44 ;
 RECT 3.96 1.81 4.09 1.94 ;
 RECT 4.91 0.565 5.04 0.695 ;
 RECT 5.79 0.3 5.92 0.43 ;
 RECT 5.385 0.385 5.515 0.515 ;
 RECT 4.435 2.305 4.565 2.435 ;
 RECT 3.965 0.325 4.095 0.455 ;
 RECT 4.91 1.61 5.04 1.74 ;
 RECT 4.91 1.91 5.04 2.04 ;
 RECT 3.96 1.54 4.09 1.67 ;
 RECT 5.79 2 5.92 2.13 ;
 RECT 5.79 2.26 5.92 2.39 ;
 RECT 4.55 1.225 4.68 1.355 ;
 RECT 4.435 1.73 4.565 1.86 ;
 RECT 5.79 0.56 5.92 0.69 ;
 RECT 3.105 0.58 3.235 0.71 ;
 RECT 1.775 1.9 1.905 2.03 ;
 RECT 3.595 2.06 3.725 2.19 ;
 RECT 1.775 1.64 1.905 1.77 ;
 RECT 3.595 0.32 3.725 0.45 ;
 RECT 2.715 2.075 2.845 2.205 ;
 RECT 3.105 0.32 3.235 0.45 ;
 RECT 1.775 0.32 1.905 0.45 ;
 LAYER M1 ;
 RECT 3.96 0.255 4.1 1.22 ;
 RECT 3.955 1.36 4.095 2.01 ;
 RECT 3.955 1.22 4.73 1.36 ;
 RECT 2.17 1.29 3.035 1.37 ;
 RECT 2.71 1.37 2.85 2.275 ;
 RECT 2.17 0.48 2.32 0.615 ;
 RECT 2.18 0.455 2.32 0.48 ;
 RECT 2.17 0.615 2.31 1.23 ;
 RECT 2.18 0.315 2.445 0.455 ;
 RECT 2.17 1.23 3.435 1.29 ;
 RECT 2.895 1.15 3.435 1.23 ;
 RECT 3.59 0.27 3.73 2.305 ;
 RECT 3.59 2.445 3.73 2.58 ;
 RECT 3.575 2.305 4.29 2.445 ;
 END
END LSDNENSSX2

MACRO LSDNENSSX4
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 3.2 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 3.2 0.08 ;
 RECT 0.45 0.08 0.59 0.535 ;
 RECT 2.68 0.08 2.82 0.89 ;
 RECT 1.785 0.08 1.925 0.785 ;
 RECT 1.39 0.08 1.53 0.535 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 3.2 2.96 ;
 RECT 0.45 1.42 0.59 2.8 ;
 RECT 2.68 1.935 2.82 2.8 ;
 RECT 1.785 1.735 1.925 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 2.265 0.83 2.455 1.1 ;
 RECT 2.265 1.1 2.405 2.585 ;
 RECT 2.265 0.275 2.405 0.83 ;
 END
 END Q

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.215 0.745 1.535 1.105 ;
 END
 END D

 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.385 0.73 0.77 1.065 ;
 END
 END ENB

 OBS
 LAYER PO ;
 RECT 1.175 0.745 1.495 1.09 ;
 RECT 1.175 0.105 1.275 0.745 ;
 RECT 1.175 1.09 1.275 2.77 ;
 RECT 0.705 0.105 0.805 0.8 ;
 RECT 0.52 0.8 0.805 1.03 ;
 RECT 0.705 1.03 0.805 2.77 ;
 RECT 2.04 0.105 2.14 1.14 ;
 RECT 2.04 1.37 2.14 2.77 ;
 RECT 1.935 1.14 2.165 1.37 ;
 LAYER CO ;
 RECT 1.325 0.875 1.455 1.005 ;
 RECT 0.455 2.09 0.585 2.22 ;
 RECT 1.985 1.19 2.115 1.32 ;
 RECT 0.57 0.85 0.7 0.98 ;
 RECT 1.395 1.805 1.525 1.935 ;
 RECT 2.27 1.545 2.4 1.675 ;
 RECT 0.925 0.335 1.055 0.465 ;
 RECT 2.27 0.325 2.4 0.455 ;
 RECT 0.455 1.545 0.585 1.675 ;
 RECT 2.27 1.805 2.4 1.935 ;
 RECT 2.685 2.005 2.815 2.135 ;
 RECT 2.685 2.265 2.815 2.395 ;
 RECT 2.685 0.69 2.815 0.82 ;
 RECT 2.685 0.43 2.815 0.56 ;
 RECT 2.27 2.065 2.4 2.195 ;
 RECT 2.27 0.585 2.4 0.715 ;
 RECT 2.27 2.345 2.4 2.475 ;
 RECT 1.395 2.08 1.525 2.21 ;
 RECT 0.455 1.81 0.585 1.94 ;
 RECT 1.395 0.335 1.525 0.465 ;
 RECT 0.455 0.335 0.585 0.465 ;
 RECT 1.79 0.325 1.92 0.455 ;
 RECT 1.79 0.585 1.92 0.715 ;
 RECT 1.79 1.805 1.92 1.935 ;
 RECT 1.79 2.065 1.92 2.195 ;
 RECT 1.79 2.345 1.92 2.475 ;
 LAYER M1 ;
 RECT 0.92 0.265 1.06 1.34 ;
 RECT 1.39 1.26 1.53 2.28 ;
 RECT 0.92 1.26 1.53 1.4 ;
 RECT 1.97 1.14 2.125 1.37 ;
 RECT 1.415 1.26 2.125 1.4 ;
 END
END LSDNENSSX4

MACRO LSDNENSSX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 8.96 BY 2.88 ;
 PIN ENB
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.3 0.735 0.57 1.005 ;
 END
 END ENB

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 1.305 0.825 1.575 1.095 ;
 END
 END D

 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 8.96 0.08 ;
 RECT 1.245 0.08 1.385 0.515 ;
 RECT 0.305 0.08 0.445 0.515 ;
 RECT 2.97 0.08 3.11 0.58 ;
 RECT 7.02 0.08 7.16 0.6 ;
 RECT 8.405 0.08 8.545 0.9 ;
 RECT 7.975 0.08 8.115 0.6 ;
 RECT 5.085 0.08 5.225 0.6 ;
 RECT 1.635 0.08 1.775 0.55 ;
 RECT 4.095 0.08 4.235 0.6 ;
 RECT 6.05 0.08 6.19 0.6 ;
 END
 END VSS

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 8.96 2.96 ;
 RECT 0.305 1.69 0.445 2.8 ;
 RECT 8.405 1.945 8.545 2.8 ;
 RECT 4.135 1.735 4.275 2.8 ;
 RECT 6.05 1.735 6.19 2.8 ;
 RECT 5.085 1.735 5.225 2.8 ;
 RECT 7.975 1.735 8.115 2.8 ;
 RECT 7.02 1.735 7.16 2.8 ;
 RECT 1.635 1.635 1.775 2.8 ;
 RECT 2.975 1.735 3.115 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 4.615 1.105 7.8 1.245 ;
 RECT 7.31 1.245 7.8 1.455 ;
 RECT 7.31 1.045 7.8 1.105 ;
 RECT 6.55 1.245 6.69 2.36 ;
 RECT 6.55 0.41 6.69 1.105 ;
 RECT 4.615 1.245 4.755 2.36 ;
 RECT 4.615 0.41 4.755 1.105 ;
 RECT 5.58 1.245 5.72 2.36 ;
 RECT 5.58 0.41 5.72 1.105 ;
 RECT 7.505 1.455 7.645 2.36 ;
 RECT 7.505 0.41 7.645 1.045 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 3.23 0.11 3.33 1.025 ;
 RECT 3.23 1.125 3.33 2.79 ;
 RECT 3.86 0.11 3.96 1.025 ;
 RECT 3.86 1.125 3.96 2.79 ;
 RECT 2.335 1.025 3.96 1.125 ;
 RECT 2.75 0.11 2.85 1.025 ;
 RECT 2.75 1.125 2.85 2.79 ;
 RECT 2.335 0.955 2.565 1.025 ;
 RECT 2.335 1.125 2.565 1.185 ;
 RECT 7.29 0.21 7.39 2.665 ;
 RECT 4.4 0.21 4.5 0.955 ;
 RECT 4.4 1.185 4.5 2.765 ;
 RECT 4.87 0.21 4.97 2.665 ;
 RECT 5.365 0.21 5.465 2.665 ;
 RECT 5.835 0.21 5.935 2.665 ;
 RECT 6.335 0.21 6.435 2.665 ;
 RECT 7.76 0.21 7.86 2.765 ;
 RECT 6.335 0.11 6.905 0.21 ;
 RECT 6.805 0.21 6.905 2.665 ;
 RECT 6.805 2.665 7.39 2.765 ;
 RECT 4.27 0.955 4.5 1.185 ;
 RECT 4.4 0.11 4.97 0.21 ;
 RECT 4.87 2.665 5.465 2.765 ;
 RECT 5.365 0.11 5.935 0.21 ;
 RECT 5.835 2.665 6.435 2.765 ;
 RECT 7.29 0.11 7.86 0.21 ;
 RECT 0.56 1.01 0.66 2.645 ;
 RECT 0.56 0.115 0.66 0.78 ;
 RECT 0.315 0.78 0.66 1.01 ;
 RECT 1.03 1.075 1.13 2.645 ;
 RECT 1.03 0.115 1.13 0.845 ;
 RECT 1.03 0.845 1.555 1.075 ;
 RECT 1.89 0.11 1.99 1.18 ;
 RECT 1.89 1.41 1.99 2.79 ;
 RECT 1.775 1.18 2.005 1.41 ;
 LAYER CO ;
 RECT 8.41 0.44 8.54 0.57 ;
 RECT 4.62 2.145 4.75 2.275 ;
 RECT 2.98 2.32 3.11 2.45 ;
 RECT 6.555 0.48 6.685 0.61 ;
 RECT 2.495 2.32 2.625 2.45 ;
 RECT 1.64 2.32 1.77 2.45 ;
 RECT 2.98 1.805 3.11 1.935 ;
 RECT 8.41 2.015 8.54 2.145 ;
 RECT 3.565 1.76 3.695 1.89 ;
 RECT 0.31 2.1 0.44 2.23 ;
 RECT 2.495 1.805 2.625 1.935 ;
 RECT 3.565 2.145 3.695 2.275 ;
 RECT 2.385 1.005 2.515 1.135 ;
 RECT 5.585 2.145 5.715 2.275 ;
 RECT 5.585 0.48 5.715 0.61 ;
 RECT 7.98 0.4 8.11 0.53 ;
 RECT 5.09 0.4 5.22 0.53 ;
 RECT 7.025 2.32 7.155 2.45 ;
 RECT 7.98 2.32 8.11 2.45 ;
 RECT 3.565 0.48 3.695 0.61 ;
 RECT 4.62 1.76 4.75 1.89 ;
 RECT 6.055 0.4 6.185 0.53 ;
 RECT 1.64 0.35 1.77 0.48 ;
 RECT 2.115 2.075 2.245 2.205 ;
 RECT 2.115 0.46 2.245 0.59 ;
 RECT 6.555 2.145 6.685 2.275 ;
 RECT 7.51 0.48 7.64 0.61 ;
 RECT 6.055 1.805 6.185 1.935 ;
 RECT 5.09 2.32 5.22 2.45 ;
 RECT 8.41 2.275 8.54 2.405 ;
 RECT 6.555 1.76 6.685 1.89 ;
 RECT 4.32 1.005 4.45 1.135 ;
 RECT 4.1 0.4 4.23 0.53 ;
 RECT 7.51 1.76 7.64 1.89 ;
 RECT 1.64 1.745 1.77 1.875 ;
 RECT 6.055 2.32 6.185 2.45 ;
 RECT 7.025 1.805 7.155 1.935 ;
 RECT 7.98 1.805 8.11 1.935 ;
 RECT 5.09 1.805 5.22 1.935 ;
 RECT 7.025 0.4 7.155 0.53 ;
 RECT 1.825 1.23 1.955 1.36 ;
 RECT 4.62 0.48 4.75 0.61 ;
 RECT 5.585 1.76 5.715 1.89 ;
 RECT 1.25 2.09 1.38 2.22 ;
 RECT 0.31 1.82 0.44 1.95 ;
 RECT 1.25 1.815 1.38 1.945 ;
 RECT 1.25 0.335 1.38 0.465 ;
 RECT 0.78 0.335 0.91 0.465 ;
 RECT 0.365 0.83 0.495 0.96 ;
 RECT 0.31 0.335 0.44 0.465 ;
 RECT 1.375 0.895 1.505 1.025 ;
 RECT 2.49 0.4 2.62 0.53 ;
 RECT 2.115 1.625 2.245 1.755 ;
 RECT 2.975 0.4 3.105 0.53 ;
 RECT 4.14 1.805 4.27 1.935 ;
 RECT 4.14 2.32 4.27 2.45 ;
 RECT 8.41 0.7 8.54 0.83 ;
 RECT 7.51 2.145 7.64 2.275 ;
 LAYER M1 ;
 RECT 2.11 0.355 2.25 1 ;
 RECT 2.11 1.14 2.25 2.3 ;
 RECT 2.11 1 2.58 1.14 ;
 RECT 2.49 1.335 3.985 1.475 ;
 RECT 3.56 0.41 3.7 1.335 ;
 RECT 3.56 1.475 3.7 2.36 ;
 RECT 3.845 1.15 3.985 1.335 ;
 RECT 2.72 0.86 2.86 1.335 ;
 RECT 2.49 1.475 2.63 2.52 ;
 RECT 2.485 0.33 2.625 0.72 ;
 RECT 2.485 0.72 2.86 0.86 ;
 RECT 4.315 0.935 4.455 1.01 ;
 RECT 4.315 1.15 4.455 1.205 ;
 RECT 3.845 1.01 4.455 1.15 ;
 RECT 1.245 1.385 1.385 2.29 ;
 RECT 0.775 0.265 0.915 1.245 ;
 RECT 1.82 1.16 1.96 1.245 ;
 RECT 0.775 1.245 1.96 1.385 ;
 RECT 1.82 1.385 1.96 1.435 ;
 END
END LSDNENSSX8

MACRO LSDNSSX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 SYMMETRY X Y ;
 SITE unit ;
 SIZE 1.92 BY 2.88 ;
 PIN VSS
 DIRECTION INOUT ;
 USE GROUND ;
 PORT
 LAYER M1 ;
 RECT 0 -0.08 1.92 0.08 ;
 RECT 1.54 0.08 1.68 0.765 ;
 RECT 0.615 0.08 0.755 0.575 ;
 END
 END VSS

 PIN D
 DIRECTION INPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.355 0.8 0.7 1.145 ;
 END
 END D

 PIN VDD
 DIRECTION INOUT ;
 USE POWER ;
 PORT
 LAYER M1 ;
 RECT 0 2.8 1.92 2.96 ;
 RECT 0.615 1.63 0.755 2.8 ;
 RECT 1.545 1.85 1.685 2.8 ;
 END
 END VDD

 PIN Q
 DIRECTION OUTPUT ;
 USE SIGNAL ;
 PORT
 LAYER M1 ;
 RECT 0.935 1.74 1.27 2.115 ;
 RECT 1.13 0.445 1.27 1.74 ;
 END
 END Q

 OBS
 LAYER PO ;
 RECT 0.915 0.095 1.015 1.14 ;
 RECT 0.915 1.37 1.015 2.79 ;
 RECT 0.805 1.14 1.035 1.37 ;
 RECT 0.395 0.1 0.495 0.865 ;
 RECT 0.395 1.095 0.495 2.185 ;
 RECT 0.395 0.865 0.625 1.095 ;
 LAYER CO ;
 RECT 1.55 2.18 1.68 2.31 ;
 RECT 1.55 1.92 1.68 2.05 ;
 RECT 0.855 1.19 0.985 1.32 ;
 RECT 1.135 0.515 1.265 0.645 ;
 RECT 0.62 0.375 0.75 0.505 ;
 RECT 0.62 2.26 0.75 2.39 ;
 RECT 1.135 1.92 1.265 2.05 ;
 RECT 1.135 1.62 1.265 1.75 ;
 RECT 0.62 1.7 0.75 1.83 ;
 RECT 0.445 0.915 0.575 1.045 ;
 RECT 0.145 1.525 0.275 1.655 ;
 RECT 0.145 0.33 0.275 0.46 ;
 RECT 1.545 0.305 1.675 0.435 ;
 RECT 1.545 0.565 1.675 0.695 ;
 LAYER M1 ;
 RECT 0.14 0.26 0.28 0.52 ;
 RECT 0.075 0.52 0.28 0.66 ;
 RECT 0.075 0.66 0.215 1.285 ;
 RECT 0.075 1.285 0.28 1.425 ;
 RECT 0.14 1.425 0.28 1.725 ;
 RECT 0.85 1.12 0.99 1.39 ;
 RECT 0.085 1.285 0.99 1.425 ;
 END
END LSDNSSX1

END LIBRARY
